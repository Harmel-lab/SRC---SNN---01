----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (    0,     0,     0,    -1,    -1,     1,     0,     0,     1,    -1,     0,     1,     0,    -2,    -2,     0,    -1,     1,     1,     0,    -1,    -1,    -1,     1,     1,     1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,     1,     2,     1,    -2,     1,     3,     1,     0,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     1,     3,     0,    -2,     0,    -2,    -5,    -1,    -1,     0,    -3,    -3,    -5,    -1,    -1,    -2,    -1,    -1,    -1,    -3,    -2,    -2,    -2,     0,    -1,     1,    -1,     0,     3,     0,     2,     1,    -4,    -3,    -2,    -3,    -3,    -5,    -3,    -5,    -5,    -1,     3,     0,    -4,    -3,    -2,    -3,    -2,     1,     1,    -1,     1,    -1,     1,     0,     0,    -2,    -4,     1,    -3,    -7,    -3,    -3,    -5,    -8,    -1,     0,    -2,    -1,    -4,    -3,    -3,     0,    -2,    -3,    -2,     1,    -1,    -2,     0,     0,     1,    -2,    -1,     0,    -2,    -1,     0,    -2,    -1,    -4,    -7,    -5,    -6,     1,     3,     0,    -3,     0,    -4,    -5,     0,    -1,    -1,    -1,    -6,    -2,    -1,    -1,     1,    -3,    -2,    -2,     0,    -1,    -1,    -3,    -3,    -2,    -8,    -6,    -2,    -1,    -3,     3,     2,     1,    -5,    -4,    -3,     1,    -5,    -2,    -5,    -1,     3,     0,    -2,    -2,    -2,     1,    -1,    -1,     1,    -2,    -2,    -5,    -8,    -8,    -3,     0,     0,     5,     3,    -5,     0,    -5,    -4,     2,    -3,    -5,    -2,    -5,     3,     4,    -6,     3,     2,    -1,    -1,    -1,     0,    -1,    -4,    -3,    -8,    -2,    -1,     2,    -3,     1,     6,    -2,     1,    -5,    -6,    -1,    -4,    -2,    -6,    -2,    -2,    -2,    -1,     6,    -1,    -1,    -1,    -4,    -1,    -3,    -7,    -3,    -1,    -2,     2,    -1,    -2,     4,     1,     0,    -4,    -9,    -1,    -1,    -2,    -3,    -5,     0,     1,    -1,    -1,     1,     2,    -2,    -3,    -1,     2,     0,    -1,    -3,    -2,    -1,     0,    -6,    -6,    -2,    -4,     1,    -4,    -4,    -2,    -4,    -5,    -2,    -2,    -4,     1,     1,     6,    -2,     1,    -3,     0,    -1,    -1,    -2,    -2,    -4,     0,     2,    -2,    -2,     1,    -3,     1,     7,    -5,    -4,     1,    -4,    -6,    -2,    -4,    -2,    -1,    -1,     2,     1,     0,     0,     1,     0,     0,    -6,     0,     1,    -1,     3,    -1,    -2,    -6,     1,     4,     6,    -1,     0,     4,     0,    -6,    -4,    -4,    -3,     1,     0,     3,     3,    -1,     0,     1,     3,    -4,    -3,     0,    -1,    -5,     2,    -4,   -11,    -9,    -1,     3,     6,     2,    -1,     4,    -2,    -4,    -3,    -2,    -5,     0,    -1,     0,     0,    -2,    -1,     2,    -3,    -4,    -3,    -1,     1,     2,     5,    -1,    -8,    -8,     0,     1,     3,     2,    -5,     0,     0,    -2,    -3,     1,    -4,     0,     0,    -1,    -2,    -2,     1,    -4,     0,    -6,    -3,    -5,    -1,     2,     7,     1,   -10,    -3,    -1,     1,    -1,    -2,    -5,     4,    -3,    -3,     0,    -3,    -3,     0,    -1,     0,    -1,    -3,     1,     0,    -7,    -2,    -5,    -5,    -3,     3,     3,    -3,   -13,     0,    -1,     8,    -2,    -1,    -4,    -3,     0,    -3,    -3,    -2,    -7,     3,     0,     0,    -4,    -2,    -6,    -2,    -4,    -3,    -4,   -10,     1,     1,     4,    -3,    -9,    -3,     0,     4,     1,     0,     2,    -3,    -1,     2,    -3,    -4,    -7,     2,     0,     1,    -2,     1,    -2,    -3,    -1,    -1,    -3,    -5,     4,     4,    -3,    -5,   -10,    -1,    -1,     1,    -1,     0,     0,    -1,     1,    -3,     0,    -1,    -3,    -2,     1,     2,     0,     2,     1,    -3,    -1,    -5,    -4,     1,     3,     3,     0,    -6,    -6,     4,     1,    -3,    -3,     0,    -5,    -2,    -2,    -2,     0,    -9,    -2,    -1,     0,     0,    -1,    -2,     1,    -1,    -3,    -6,    -5,     2,     1,    -3,    -4,    -1,    -1,     1,     1,    -3,     0,    -5,    -3,    -4,    -1,    -1,    -1,    -2,     1,     1,     0,    -1,    -3,    -3,    -1,    -2,     0,    -4,    -2,    -1,     1,    -1,     0,    -1,    -1,     2,    -1,    -1,    -3,    -5,    -5,    -3,     1,     0,    -5,     0,     2,     2,     0,     1,    -2,    -7,     1,     0,     1,     0,    -2,     2,     1,     3,    -1,    -5,     4,     3,     4,    -8,    -3,    -4,    -3,    -2,     1,    -1,     0,    -1,     2,     1,     0,     1,    -3,    -5,    -2,     1,    -2,    -1,    -2,    -5,     3,     2,     3,     3,    -4,    -3,    -4,    -9,     0,    -5,    -4,    -2,     3,     0,    -2,    -5,    -3,    -1,     1,    -1,    -1,     0,    -3,     3,     2,     1,    -5,    -6,    -4,    -4,     1,     6,     1,     1,    -6,    -2,    -1,    -4,    -4,     2,    -2,    -3,     0,    -1,    -1,     1,     0,     1,     0,    -1,    -9,    -4,    -3,    -3,    -1,    -3,    -5,    -6,    -9,    -9,   -11,    -4,    -3,    -3,    -3,    -2,    -5,    -2,    -3,    -2,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -4,    -6,     1,     0,    -4,    -2,    -1,    -3,    -3,    -3,    -3,    -2,    -5,    -7,    -3,    -5,    -3,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,    -1,    -1,     1,    -1,     1,    -3,     1,     0,    -2,     0,     1,     0,    -1,    -2,    -2,    -2,     0,     0,    -1,     1),
		     1 => (    0,    -1,     0,     1,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -1,     1,     1,     0,     0,    -1,     1,    -1,    -1,     1,    -1,     0,     0,    -1,     1,     1,     1,     1,     1,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,     4,     3,     0,    -2,    -1,     1,    -1,    -1,     0,    -1,    -1,     1,    -1,     1,     1,     0,     0,     1,     0,     0,     1,     1,    -4,    -3,     0,    -1,    -1,    -1,    -2,    -4,    -5,    -6,    -7,     1,     2,    -6,    -2,     0,    -1,    -2,     0,     1,     1,    -1,     8,     5,     0,     1,     1,     6,     5,     3,     3,     2,     1,    -9,   -10,   -10,    -8,    -2,    -3,    -1,     1,    -5,     2,     0,    -3,     0,     1,     1,     0,     0,     5,     4,     2,    -1,    -1,     0,     0,    -1,    -4,    -9,    -9,   -10,     1,     4,     0,     1,     2,     2,     1,     2,    -3,   -10,    -5,    -9,    -5,    -5,     0,    -1,     5,     7,     2,     1,    -2,    -2,   -12,    -5,    -4,    -8,   -10,    -6,    -1,     7,     0,    -1,     0,     3,     3,    -3,    -4,   -10,    -7,    -5,    -5,    -4,     0,    -1,     0,     3,     2,    -2,     0,     1,   -10,     1,     1,    -7,    -8,    -4,    -6,    -2,    -1,     2,     0,     3,    -3,    -3,    -2,   -10,    -7,    -3,     0,    -2,    -1,     0,    -2,     2,     1,     0,    -2,    -4,   -11,    -2,    -6,    -9,    -7,    -1,     4,     2,     2,    -1,     5,    -1,    -4,    -3,     0,    -7,    -7,    -3,    -3,    -2,     0,    -2,    -2,    -1,    -1,    -2,    -4,    -4,    -8,    -7,    -3,   -12,   -11,     0,     3,     2,     4,     3,     2,    -3,    -4,    -2,    -4,    -6,    -7,    -4,    -4,    -1,     1,     0,    -2,     2,    -1,     0,    -6,    -3,    -2,    -3,    -9,   -16,    -4,    -1,    -2,     0,     5,     1,    -5,    -3,    -7,    -3,    -2,    -4,    -7,    -3,     0,    -4,     0,     1,    -1,    -2,    -1,    -1,    -5,    -7,    -4,    -6,    -1,    -8,    -6,    -3,     1,     6,     5,    -1,    -5,    -5,    -7,    -3,    -2,    -3,    -7,    -8,     0,     8,     0,     0,     1,     2,     2,     1,    -3,    -4,    -6,   -10,    -5,    -9,    -2,    -4,     0,     7,     1,    -7,    -4,    -2,    -2,     1,    -2,    -4,    -8,    -7,     0,     7,     0,     0,    -2,     6,     1,    -1,    -2,    -2,   -10,    -9,    -5,    -5,     0,    -2,     5,    -1,     3,   -10,   -11,    -4,     5,     7,     7,     5,    -2,     0,    -1,     4,     0,    -1,     0,     2,     3,    -2,    -3,    -1,    -5,   -11,    -5,    -3,    -2,     1,     6,    -2,     2,    -9,   -11,     1,     4,     1,     0,    -8,    -5,     0,     2,     1,    -1,     1,     3,     3,     3,    -6,    -4,    -3,    -1,    -7,    -5,     2,    -1,    -4,     6,     0,    -4,    -9,    -1,     6,     6,     8,     5,    -2,    -4,     8,     7,     0,     1,     0,     3,     7,     3,    -1,    -2,    -1,     4,     0,    -2,     4,     0,    -2,    -2,    -6,    -5,    -7,    -3,    -6,    -1,     9,     4,    -4,   -10,     3,     2,    -1,     1,     1,     1,    -3,    -2,    -1,     2,     0,     4,     3,     2,     5,     2,     2,    -4,    -2,    -2,    -9,    -7,    -8,    -1,     6,     4,     8,    10,    -2,    -2,     0,     1,    -1,     1,    -4,     1,     1,     4,     1,     3,     1,     1,     2,    -1,     2,     2,    -2,    -4,    -3,     2,     4,     5,     8,     8,     9,     6,     0,    -2,    -3,    -3,    -1,     0,    -2,    -2,    -3,    -4,    -2,     1,    -4,     1,    -2,    -1,     3,    -4,   -10,    -7,     2,     5,     6,     3,     1,     1,     0,     3,     5,     1,     4,    -1,    -1,     4,     4,    -5,     4,     5,     1,     0,    -4,    -1,     2,     2,     3,    -6,    -7,   -11,    -2,     3,    -1,    -1,    -2,    -6,     1,     5,     7,     1,     3,     0,    -1,     4,     1,     0,     7,     3,    -4,     0,    -2,    -5,     2,     0,     3,    -3,    -8,    -9,    -2,    -2,    -1,     5,    -6,    -3,     0,     3,     2,     3,     0,     5,     3,    -2,     0,     0,    -6,    -9,    -3,     0,    -2,     0,    -2,     3,    -4,     0,    -2,    -8,    -8,    -7,    -2,     3,     2,     2,     2,     3,     3,     1,     1,     4,     4,     1,     0,     0,    -5,   -11,    -2,     0,    -3,     2,    -3,    -1,    -1,     3,    -4,    -3,    -7,     1,     5,     8,     3,     5,     4,     4,     7,    10,     1,    -1,    -1,    -1,     0,    -4,    -1,    -4,    -4,     4,    -3,    -1,     2,     0,     1,     2,    -1,     1,     1,     2,     6,     7,     1,    -1,    -2,     3,     5,    10,    -1,     0,     0,    -1,    -1,    -3,    -6,    -2,    -5,    -3,    -5,    -8,    -3,    -4,   -10,     4,     3,    -1,     1,     1,    12,     8,     1,    -1,     1,    -2,     2,     3,     0,     1,     1,     0,     0,     0,    -1,    -1,    -1,    -4,     3,    -8,    -4,    -7,    -6,    -6,    -9,    -4,    -5,    -4,    -4,    -5,    -4,    -3,    -2,    -2,     0,    -1,     1,    -1,    -1,    -1,    -1,    -2,    -4,    -5,    -3,    -3,    -4,     2,    -1,    -7,    -6,    -8,    -9,    -7,    -5,    -1,    -2,    -1,    -1,     0,     1,    -1,     1,    -1,     0,    -1,     0,    -1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -2,     1,     1,     2,     0,    -1,     0,    -1,    -1,     0,     1,    -1,     1,     1,     0,     1,     1),
		     2 => (    0,    -1,     1,    -1,    -1,     1,     1,     1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,     1,     1,    -1,     1,    -2,    -4,    -2,    -2,    -1,    -6,    -4,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -2,     0,     1,     1,     1,     0,    -1,     0,    -3,    -4,     0,     1,    -6,    -2,    -3,    -3,    -5,    -2,   -12,    -4,    -1,    -2,    -3,    -5,    -6,    -5,    -1,    -3,     1,     1,     3,     1,     1,     0,     1,    -2,    -5,    -5,     0,     6,    -2,    -1,     5,     5,     1,    -5,    -7,    -4,    -7,    -6,    -2,     3,    -2,    -7,    -4,    -1,    -3,    -4,     2,    -1,    -1,    -1,     1,     0,     3,    -2,    -3,    -1,     5,     1,    -1,    -5,    -4,    -3,    -8,    -8,    -5,     2,     2,     0,    -3,     3,     4,    -1,    -6,     1,     1,    -3,    -1,     0,     1,    -2,     1,     6,     1,     0,     0,    -1,    -2,    -6,    -8,    -9,    -9,    -7,    -3,    -1,     1,     4,     4,     3,     5,     1,    -5,    -4,     0,    -4,    -1,     1,     1,     2,     1,     1,    -1,    -2,     3,     2,    -2,    -2,    -3,    -1,    -9,    -7,    -6,    -3,     5,     2,     4,    -1,     2,     1,    -7,    -6,     6,    -4,    -1,     1,     1,     5,     0,     0,    -3,     0,     4,     0,     1,     0,     3,     2,     4,    -3,    -3,    -3,    -2,    -7,    -2,     2,     1,     1,   -12,    -1,     9,    -4,    -1,    -7,     6,     6,    -4,    -2,     2,     0,    -2,    -3,    -7,     1,     4,     0,     2,     3,    -8,   -10,    -4,    -4,     1,     3,    -1,    -1,     1,     1,     4,    -6,    -2,     0,    -3,     6,    -3,    -5,    -1,    -1,     0,    -4,    -3,     2,    -2,    -4,     0,     2,     1,    -3,    -3,    -1,     5,     2,     2,     2,    -1,    -1,    -6,     4,    -2,    -1,    -2,     5,    -7,    -4,     3,     3,     4,    -1,     0,     1,     0,     3,     6,    12,     4,    -4,    -2,     1,     6,     2,     3,     1,    -6,    -3,    -4,     3,    -3,     1,    -5,    -4,    -5,     3,     1,     3,     6,     6,     3,    -3,    -2,    -7,    -2,     0,     0,     0,    -6,     0,     3,     0,     2,     1,    -6,     0,    -2,     2,    -5,    -1,     0,   -10,    -3,     5,     4,     3,     3,     0,     2,     0,    -8,    -9,    -5,    -4,    -3,    -4,    -4,    -3,     1,     3,     0,    -1,    -9,    -2,     1,     7,     0,     0,     0,    -1,     4,    -1,    -5,    -6,    -7,   -12,    -4,    -3,     0,    -5,    -8,    -5,    -6,    -4,     0,    -1,    -1,    -2,    -5,    -2,    -2,     3,     4,    11,     2,    -1,     0,    -2,     0,    -6,    -9,    -3,    -4,    -7,    -9,    -7,     2,     3,    -6,    -8,    -3,     3,     2,    -2,    -3,    -8,    -5,     1,     2,     0,     4,     8,     3,     1,    -2,     1,     2,     2,    -2,    -5,   -10,    -5,    -6,     2,     1,     5,     2,     0,     2,    -2,     3,     3,     0,    -2,     0,     1,     2,     2,     2,     3,     5,    -1,     0,     1,     3,     5,     2,    -3,     1,    -2,    -1,     1,     2,     3,     0,     5,     6,     6,     9,     0,    -6,   -11,    -6,    -3,    -2,    -2,     2,     6,     5,     1,    -2,     3,     4,     0,     3,     0,    -4,     0,    -2,     3,    -2,     6,     0,     1,     0,     2,    -1,    -3,    -5,    -3,    -1,     1,    -1,     1,    -1,     5,     7,     1,     0,    -4,     8,     5,     8,     6,    -1,    -3,    -1,    -1,    -4,    -2,     3,     2,     5,     3,    -1,    -1,    -2,     0,    -2,     0,    -1,     7,     1,     7,    12,     1,    -1,    -1,     7,     9,     4,     4,     1,    -1,    -2,     6,     3,     3,    -1,    -1,     2,     3,     3,    -1,    -5,    -3,     0,     4,     2,     8,     5,     8,     9,    -1,     1,     2,     4,     5,     5,     6,     4,     1,     0,     0,     0,    -4,     0,     0,     5,     3,    -2,    -1,     0,    -3,     0,    -2,     4,     8,     2,     8,    -1,     0,     2,     1,    -1,     5,     7,    -1,    -2,    -2,    -2,    -2,    -4,    -4,    -9,    -5,     1,     1,     4,     8,     6,     3,    -6,     0,     5,     6,     5,     7,     0,     0,    -1,     4,     2,     6,     0,    -5,    -6,    -4,    -3,    -5,    -6,    -8,   -10,    -4,     1,    -1,     4,     3,     1,    -3,    -1,    -1,     1,     5,    -3,    -4,     0,    -1,     0,     2,     2,     3,     1,    -1,    -2,    -1,    -5,    -6,    -6,    -9,    -7,    -5,     1,    -8,   -15,    -5,     0,    -1,     1,    -4,    -4,    -1,     2,    -1,    -1,     1,     1,    -3,     2,    -4,    -5,    -1,    -3,    -1,    -9,   -10,    -9,    -9,   -10,    -5,    -4,   -11,   -17,    -9,     3,     1,     2,    -4,    -2,     3,     0,     0,    -1,     0,     0,    -1,    -3,    -5,    -7,    -7,    -6,    -7,    -8,    -8,    -5,    -3,    -8,     2,    -2,    -6,    -6,   -12,   -11,    -5,     1,    -4,    -5,    -2,     1,     1,     0,     0,    -1,     0,     1,    -4,    -4,    -4,    -5,    -3,   -10,    -5,    -2,    -3,    -4,    -2,    -6,    -6,    -7,   -10,   -10,    -7,    -7,    -6,     0,    -1,     1,     1,     0,     1,     1,     0,     1,     0,    -1,     0,     0,    -1,    -1,    -4,    -3,    -1,    -4,    -3,    -3,    -3,    -2,    -2,    -3,    -8,    -8,    -3,     0,     0,     0,     1,     0),
		     3 => (    0,    -1,     0,     1,     0,    -1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     1,     1,     0,     0,     0,     1,     1,     1,    -1,    -1,     1,     1,     1,     0,     1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -3,    -3,     1,     0,     1,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,     1,    -1,     1,    -2,    -1,    -1,    -5,    -5,    -2,    -4,    -5,    -3,    -4,    -7,    -8,    -7,    -4,   -11,    -9,   -10,    -3,    -1,     0,     0,     1,     1,    -1,     1,    -1,    -1,    -3,    -2,    -4,    -4,    -4,    -5,    -4,     0,    -1,    -5,    -5,     1,     6,     3,    -3,    -1,    -2,    -7,    -9,    -4,    -1,     0,    -1,     0,     1,    -1,     2,     6,     2,     0,     3,     4,     7,     6,    -1,     0,     3,     5,     1,    -4,    -1,     4,     0,    -1,    -8,    -4,   -16,   -10,    -1,    -3,     1,     1,     0,     1,    -2,     2,    -3,    -4,    -5,     1,    -4,     2,     2,     0,    -1,    -1,     0,     0,     2,     4,     2,     1,     4,     2,    -2,    -4,    -3,    -3,     0,     1,     1,     1,    -1,    -3,    -1,    -1,     0,     3,     0,     1,    -1,     2,     8,     3,     0,    -1,     0,     0,     5,    -5,    -3,     1,     0,     0,    -4,    -5,    -1,     1,     2,     0,    -5,    -2,     6,     0,    -1,     1,     0,     3,     5,     1,    -3,     1,     3,     5,     0,    -1,     0,     5,    -1,    -4,    -8,    -5,    -7,    -5,    -1,     1,    -1,     1,     7,     3,     2,    -4,     4,    -1,    -6,     4,     2,     5,     2,     0,    -2,    -1,     2,    -1,     1,     3,     3,    -1,   -13,   -14,    -4,    -6,    -1,    -1,    -3,     9,     8,     2,    -8,    -3,    -1,    -3,    -1,    -5,    -4,   -10,   -12,   -18,    -8,     2,     1,     2,     3,     3,     2,     1,    -9,   -18,    -8,    -8,     0,     0,    -2,    12,     5,    -5,    -9,   -10,   -15,   -12,   -13,   -12,   -22,   -18,   -16,    -7,    -2,     1,    -2,    -1,     1,     1,     4,     3,    -3,   -17,    -4,    -5,    -1,     0,    -2,    -2,    -3,    -7,    -9,   -14,   -10,   -15,   -20,   -14,   -12,    -6,     4,     7,     7,     1,     2,     0,     3,     8,     5,     4,    -9,    -8,    -7,    -3,     0,    -1,     0,    -5,    -7,     2,    -2,    -2,    -6,    -3,    -6,    -3,     1,     7,     6,     4,    -2,     1,    -2,     3,    -6,    -1,    -1,    -2,    -3,     0,    -1,    -2,    -1,     0,     0,    -6,     1,     8,     5,     0,    -3,     1,    -3,     2,     5,     3,     4,    -2,     0,     0,    -5,    -5,    -8,    -5,    -1,    -2,     0,    -5,    -5,    -2,    -1,    -2,     1,    -1,     0,     1,     7,    -3,    -5,     7,     2,    -1,     2,     2,     2,    -1,     1,     0,    -1,    -1,    -4,    -6,    -2,    -5,    -6,    -7,   -12,    -4,    -2,    -2,     4,     5,    -2,     4,    -1,    -9,   -11,    -7,    -4,     1,     2,     0,     5,     5,    -1,    -2,     1,    -1,     0,    -2,    -1,    -7,    -1,    -5,    -4,    10,     0,    -1,     1,     4,     5,     3,     0,   -14,   -10,   -15,    -8,    -5,     1,    -1,     3,    -2,    -3,     1,     0,     0,     3,     1,     3,    -5,    -3,    -8,    -4,     4,    -1,     0,     2,     6,    -1,    -6,    -2,    -9,    -3,   -10,   -19,   -23,   -10,   -10,   -10,    -6,    -4,     3,     2,     3,     0,    -2,     3,     1,    -4,    -8,    -8,    -3,    -1,    -2,     2,     8,     2,    -5,     4,     1,     6,    -1,    -3,    -8,    -6,   -12,   -11,    -5,     2,    -2,     0,    -2,     2,     4,     3,    -1,   -10,   -14,    -5,    -3,    -3,    -1,    -1,    -6,     9,     1,     2,     3,     1,     3,    -3,    -2,    -5,    -4,     3,     0,     0,    -1,    -2,     0,     0,    -1,    -3,    -5,    -6,   -11,    -4,    -4,    -2,    -1,     1,   -10,     7,     6,     0,     0,     0,     4,     1,     3,     2,     2,     2,    -2,    -4,     0,     0,    -2,    -2,     0,    -4,    -8,   -10,    -9,    -2,    -2,    -1,    -2,     1,    -1,     3,     8,     0,    -3,     2,     6,     0,     4,     2,     1,    -3,    -3,    -4,    -5,     2,    -1,    -6,    -3,    -3,    -5,   -10,    -8,    -3,     0,     1,    -1,    -2,    -1,     3,     2,     3,    -2,    -4,    -1,    -3,     0,    -1,    -4,    -3,    -4,    -2,    -1,     3,    -6,    -1,    -6,    -7,   -10,   -10,    -8,    -4,    -1,    -1,    -1,     1,     5,     5,     1,     7,    -4,     1,    -3,    -1,    -2,     1,    -1,     0,     2,     0,     7,     0,     0,     7,    -3,    -8,   -14,   -10,    -5,    -7,    -1,     0,     0,     0,    -1,     2,    -3,    -3,     1,    -2,    -3,     2,    -2,    -3,    -3,    -6,    -2,    -4,    -4,    -6,    -2,    -8,    -8,    -7,    -8,    -3,    -4,    -1,     0,     0,     0,     0,     0,    -5,    -2,    -1,    -4,    -6,    -4,    -1,     2,    -6,     0,    -1,    -3,    -9,    -9,    -8,    -3,    -2,     0,    -3,    -7,    -5,     0,    -2,     1,     0,    -1,    -1,     0,    -4,    -1,     1,    -3,    -6,    -9,   -10,    -4,    -6,     2,     6,     4,     1,    -4,    -5,    -3,    -4,    -7,    -4,    -5,    -1,     1,    -1,     1,    -1,     1,     1,     1,     0,     0,     0,    -1,     0,     0,    -3,     0,    -2,     0,    -2,    -4,     0,    -4,    -3,     0,    -1,    -3,    -1,    -1,    -1,     0,     1,    -1,     0),
		     4 => (    1,    -1,     0,     0,    -1,     1,     1,    -1,    -1,     0,    -1,     0,    -2,    -2,    -2,    -1,    -1,    -1,     0,     1,     0,     0,     1,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     0,     0,    -3,    -5,    -2,    -2,    -4,    -2,    -5,    -8,    -4,    -4,    -4,    -3,    -1,     1,    -3,    -2,    -3,    -3,     0,     0,     1,     0,     1,     0,    -1,     1,    -4,    -1,    -5,    -5,    -8,    -3,    -4,    -9,    -5,    -6,    -3,    -3,    -8,    -6,    -6,    -1,    -7,    -7,    -6,    -5,    -2,    -4,     1,    -1,    -1,     0,    -1,    -4,    -9,    -4,    -7,    -4,    -4,    -5,    -3,    -6,    -6,    -5,    -5,    -6,    -9,   -11,    -5,    -1,     1,    -1,    -2,    -2,    -5,    -3,    -1,    -1,    -1,    -1,    -2,    -8,    -1,     1,     6,     2,    -3,    -8,    -5,    -3,    -2,    -7,   -12,    -9,    -6,    -9,    -5,    10,     4,     1,     6,    -3,    -4,    -2,    -4,    -1,    -1,    -1,    -4,    -3,    -1,     1,     5,    -2,    -1,    -3,    -2,    -2,    -2,   -11,   -12,     1,    -5,     2,    -4,     1,     1,     1,     1,    -7,    -3,    -2,    -2,    -1,     1,     0,     0,    -1,    -3,    -3,     6,    -5,     2,     4,     1,    -4,    -8,   -17,   -16,    -9,    -2,     1,     6,     0,     0,     1,    -6,    -7,    -8,    -2,     0,    -3,     1,    -5,    -1,     1,    -1,    -2,     3,     0,     1,     1,     2,     2,    -8,   -14,   -19,    -8,    -3,     9,     6,     6,     2,    -1,    -5,    -7,    -7,     0,    -2,    -7,    -5,   -11,     1,    -1,     3,     2,     4,    -1,     2,     6,    -1,    -2,     1,   -15,   -13,    -6,     8,     6,     3,    -2,    -5,     3,    -1,    -3,    -4,     1,    -6,   -10,    -1,    -7,     1,     1,     7,     3,    -8,    -2,     5,     1,     3,     4,     5,    -7,   -11,    -1,    12,     2,     1,     0,    -6,    -2,    -3,     1,    -7,     1,    -6,    -5,     1,    -4,     0,     3,     2,    -1,   -14,    -4,     2,     5,    -1,     2,     5,    -8,    -9,     6,     6,     1,     4,     3,    -4,    -8,    -5,    -9,    -9,     2,     0,    -3,     0,    -5,     2,     1,     4,     1,    -5,    -1,     2,     1,     3,     3,     1,   -12,   -12,     1,     3,     0,     2,    -3,    -7,    -7,    -3,    -7,    -3,     2,    -2,    -7,     1,    -3,     3,     3,     4,     4,     1,     1,    -5,    -3,     3,     0,     1,    -3,    -8,     3,     0,     1,     0,     1,    -5,     0,     5,    11,    10,     9,    -8,    -6,     0,    -3,    -5,     0,     6,     2,    -2,     0,    -2,     3,     5,     0,    -1,    -1,    -3,    -3,     2,    -1,     3,     0,     1,     5,    10,     5,     1,    -1,    -8,     0,    -1,    -1,    -5,     0,     3,     8,     1,     5,     2,    -1,    -1,    -2,    -2,    -1,    -5,     0,    -2,     1,     2,     5,     1,     7,     6,    -1,     3,    -3,    -5,    -1,     1,     1,     1,    -1,     6,    -1,    -1,     5,     0,     1,     0,     2,     1,     4,     3,     5,     3,     2,     2,     5,     0,    -1,     2,    -4,    -6,    -6,     3,    -1,    -1,    -1,    -7,     4,     6,    -3,    -4,     6,     0,    -2,     1,     0,    -1,     2,     5,     4,     0,    -3,     3,     0,    -1,     2,    -5,    -6,    -1,    -2,    -3,     0,     0,    -1,     6,     5,    10,     0,    -6,     1,    -4,     1,    -6,    -4,    -2,    -3,     1,    -4,    -5,    -5,    -1,    -9,    -3,     2,    -3,    -4,     0,    -1,     1,     1,    -5,    -1,     5,     6,     7,    -5,    -6,    -6,    -3,    -1,    -4,    -5,    -3,    -2,    -3,    -9,    -7,    -3,    -6,    -6,    -2,     1,     1,    -2,    -2,    -3,     1,     0,     0,     0,    -2,     2,    -1,    -8,    -1,    -8,    -5,    -2,    -1,    -1,    -5,     0,     1,    -1,    -6,     2,    -5,    -1,    -2,     6,     2,     0,    -3,    -5,    -1,     0,     0,     0,    -1,    -5,   -12,    -8,    -7,    -2,    -5,    -7,    -4,     5,     2,    -1,     1,    -1,    -1,    -1,     4,     0,    -3,    -2,     0,    -1,    -1,   -10,    -1,    -1,    -3,    -3,    -2,    -7,    -4,    -7,    -5,    -5,    -2,    -6,    -2,     1,     1,    -2,     3,    -5,     1,    -4,    -2,    -4,    -5,    -8,    -2,     2,     1,    -9,    -5,    -1,    -1,    -3,    -1,    -3,    -1,     0,     0,    -6,     1,    -9,    -6,     0,     1,    -3,    -1,    -3,    -1,    -3,    -2,    -6,    -5,    -7,     1,     4,     0,     1,     2,    -1,    -1,    -1,    -2,    -3,     0,    -2,     4,     4,     1,   -11,    -1,    -3,    -4,    -3,    -2,    -4,     0,     0,     5,    -5,    -6,    -1,    -3,     2,    -3,     2,     1,    -1,    -1,     1,    -1,     1,    -9,    -2,    -4,    -2,    -1,    -2,    -5,    -2,    -4,    -3,     8,    -1,     5,     4,     6,    -6,    -1,     1,    -1,     0,    -7,     0,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -5,   -14,    -8,    -6,    -4,    -6,    -5,    -5,     1,     2,    -5,     0,     2,     0,    -3,    -1,     3,    -4,     2,    -3,    -1,    -2,     1,    -1,     0,     1,    -2,    -2,    -1,    -4,    -6,     1,    -1,    -8,   -13,   -11,    -8,    -4,    -6,   -11,    -3,    -7,    -9,   -11,   -11,    -9,    -2,    -3,     0,     1,    -1,     1,     0,     0,     0,    -1,     1,    -4,    -3,    -4,    -5,    -4,    -8,    -5,    -3,   -10,    -3,    -4,    -6,    -4,    -6,    -7,    -6,    -5,    -2,    -1,     0,     0,     1),
		     5 => (    1,     0,    -1,     1,     1,     0,     0,     1,    -1,     1,     1,     0,     0,     0,     0,     1,    -1,    -1,     1,     1,    -1,     0,     0,     0,     1,     1,     1,     1,     1,     1,     1,    -1,     1,    -1,     0,     0,     1,     1,     1,    -1,    -3,    -2,    -3,    -2,    -2,    -3,    -1,    -1,    -2,     0,     0,     0,    -1,     1,    -1,     1,     1,    -1,     0,    -1,    -1,    -1,     1,     1,    -1,     0,    -4,    -9,    -8,   -11,    -4,     4,     4,     5,     7,     6,     7,     5,     5,     6,    -3,    -1,     0,    -1,     1,     1,    -1,     2,     5,    -1,    -3,    -2,    -2,    -6,    -7,    -6,    -2,    -5,     4,    -2,    -8,    -6,    -1,    -2,     2,     4,    -2,    -1,     3,     3,     4,     1,     1,    -2,    -2,     1,    -6,    -6,    -8,    -9,   -13,    -4,   -10,    -7,    -7,     0,     7,     0,     2,     0,     0,    -1,     1,     4,     5,     5,     7,    13,     4,    -1,     0,    -1,    -1,    -1,    -6,    -6,   -11,   -11,   -14,    -7,    -1,    -1,     2,     0,     1,    -2,     2,     5,     3,     1,    10,     8,     4,     8,     9,    13,     6,    -2,     1,     0,     2,    -2,    -6,   -10,   -10,    -6,    -3,    -6,    -2,     1,     6,     0,     0,     1,     3,     5,    10,     1,     8,     0,     1,     8,     3,     6,     4,     1,     0,     1,    -1,    -3,    -5,    -7,    -3,    -1,    -2,     0,     0,     6,     4,     1,    -2,    -3,     1,     3,     4,     0,     4,     0,    -4,    -1,    -3,     3,     3,     2,    -1,    -1,    -4,    -3,    -4,    -3,    -6,    -3,    -5,    -7,     2,     7,     4,    -5,    -5,    -8,   -15,    -8,    -8,   -20,   -10,   -11,    -8,    -3,    -2,    -1,     2,     1,     0,    -2,    -8,    -9,    -8,    -1,    -7,    -8,    -7,    -4,    -4,    -2,    -3,    -4,    -8,   -19,   -24,   -27,   -30,   -29,   -20,   -15,   -14,    -8,    -5,    -4,     0,     1,     1,    -2,    -1,    -4,    -1,    -2,    -5,    -3,    -1,    -3,    -4,     1,    -4,     1,    -6,    -2,     0,    -6,   -17,   -18,   -17,   -14,   -14,    -9,    -5,     0,     1,     1,    -1,     0,    -1,    -3,    -1,    -3,    -5,    -5,    -4,    -5,    -4,    -2,    -2,     0,    -3,    -3,     2,     1,     2,    -3,    -9,   -14,   -10,    -5,    -6,    -1,     2,    -2,     1,    -1,     0,    -3,    -1,    -2,    -2,    -4,    -2,    -4,    -2,     2,     2,     2,     2,     1,     1,    -3,    -3,     0,    -3,    -5,    -8,    -5,    -2,    -2,     0,    -3,     0,     0,    -1,    -1,     0,     2,    -3,     1,    -5,     2,     4,     7,     3,    -1,     3,     1,    -1,    -1,    -4,     1,     1,     3,    -3,    -2,    -4,     0,    -1,    -2,     2,    -1,    -1,     1,     4,    -4,    -7,    -6,    -1,    -2,     4,     1,     0,    -3,     1,    -5,     4,     1,     1,    -4,     0,     1,     0,     0,    -2,    -1,    -2,    -2,     0,    -4,    -2,    -2,     4,    -4,    -7,    -5,    -6,    -3,    -3,    -2,     3,    -3,    -6,    -2,    -5,     3,    -2,    -1,    -3,     1,    -1,     1,     1,    -1,    -1,    -1,     0,     1,    -3,     1,     0,    -6,    -7,   -10,   -10,   -16,   -13,    -8,     1,     1,    -4,     2,     1,     8,    -2,     3,     2,     2,     3,    -4,    -5,    -3,    -3,    -4,    -1,    -2,    -7,     2,    -3,    -4,    -5,   -10,    -5,   -13,   -17,    -6,    -7,    -9,    -7,     2,    -2,    -3,     7,     4,     4,     3,    -2,    -3,    -8,    -4,    -1,    -2,     0,    -2,     0,     4,     0,    -3,    -5,    -1,     4,    -2,    -1,    -5,   -13,    -7,    -1,    -3,     2,     0,     5,    -2,    -1,     2,     0,    -3,    -7,     1,    -6,    -5,     0,     0,     5,     0,     1,    -4,    -1,    -2,     3,     4,     1,     4,     3,     2,     3,    -1,     2,    -1,     2,     2,     2,    -2,     0,    -4,    -7,     0,    -2,    -3,    -1,    -1,     3,     2,    12,    -1,     1,     0,     6,     5,     1,     2,    -5,     5,     5,     2,     1,     0,    -2,     4,     3,    -3,     4,    -7,    -5,    -3,    -1,     0,     1,    -2,    -3,    -2,     8,     6,     0,    -1,     1,     0,     2,     4,     2,     3,    -1,     2,     2,    -3,    -4,     3,     4,     5,     4,     1,    -3,    -4,     0,    -1,     1,     0,    -5,     1,    -4,    -2,    -4,    -2,    -3,    -2,     6,     1,     3,    -3,     0,    -3,     0,    -1,     2,     1,     6,    -2,    -2,    -3,    -4,    -4,     0,     0,     0,    -1,     2,     3,    -4,    -3,     1,     1,     7,     4,     1,    -6,    -2,    -2,     0,     7,    -1,    -7,    -6,    -5,    -6,    -5,     1,     2,   -10,   -10,     1,     0,    -1,     0,    -4,     0,     6,     5,    14,     7,    -1,     4,     8,     0,     2,     1,     5,    -4,    -7,    -3,    -5,    -6,    -1,     3,     4,    -1,     0,    -3,    -3,     1,    -1,     0,    -1,     5,    -3,    -1,     5,     7,     2,     5,     5,     4,     2,     1,    -3,    -2,    -3,    -7,     2,     3,     1,     2,     3,     1,    -1,     0,    -1,    -1,    -1,     1,     1,     0,    -3,    -3,    -2,    -1,     0,    -1,     3,     3,     2,    -2,    -3,    -1,    -1,    -1,    -2,    -1,     1,     1,     2,    -1,     1,     0,     1,     0,     0,     0,     1,    -1,     0,     0,    -1,     1,     0,    -1,     1,    -1,     0,     1,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -2,     1,     1,     0,     1,    -1),
		     6 => (   -1,     0,     1,     1,     1,    -1,    -1,    -1,     0,     1,     0,     1,     3,     2,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,    -1,     0,    -1,     1,     0,     1,     1,    -1,    -1,     1,     0,     2,     3,     5,     6,     5,     2,     6,     4,    -2,     0,     3,     5,     0,     4,     5,     4,     4,     5,     1,     1,    -1,     1,     1,     1,     2,     4,     5,     3,     4,     4,     1,    -1,    -3,     4,     7,     3,     3,     9,     5,     2,     3,    -1,    -2,     0,     1,     0,     2,     2,     0,    -1,     1,     0,     0,    11,     6,    -1,     5,     7,    -2,     1,    -3,     2,     2,     5,     2,    -2,    -2,     0,    -4,    -1,     4,     0,    -1,    -2,    -2,     0,     1,    -1,     0,     1,    -4,     5,     0,     3,     3,    -2,     1,     0,     2,     3,    -4,    -1,    -1,    -5,    -3,    -3,    -4,     7,     5,     3,    -3,    -6,    -3,    -4,    -1,     2,    -1,     1,     1,    -2,     0,    -7,    -6,    -2,    -4,     4,     0,    -3,     3,     4,    -2,    -3,    -6,     1,     2,     4,     2,     0,    -4,    -6,    -4,    -2,     1,     3,    -1,    -1,     1,    -5,    -5,   -10,    -8,    -1,    -4,     0,    -6,     4,     6,     1,    -1,    -2,    -2,    -5,     2,    -1,    -5,    -1,    -7,    -9,    -2,    -2,     4,    -1,     0,    -1,     0,    -5,    -5,   -12,    -8,    -4,    -2,    -2,     1,     7,     5,     0,     3,    -4,    -5,    -5,   -12,    -9,    -9,    -5,    -8,   -10,    -6,    -4,     2,    -6,     0,     0,     1,    -6,    -4,   -13,    -2,    -2,    -6,     3,     2,    -1,     5,     1,    -4,    -9,    -8,   -14,   -13,   -12,    -8,    -9,   -16,   -12,   -10,    -7,    -2,    -5,     1,    -1,    -2,    -3,    -3,   -14,    -1,     1,    -1,    -4,    -3,     1,    -3,    -6,    -5,   -11,   -10,   -14,   -14,   -12,    -8,   -14,   -13,    -9,    -2,    -3,    -3,    -2,    -1,     0,    -2,    -4,    -7,   -12,    -7,     1,     3,     0,    -4,     0,     3,    -4,   -12,   -12,    -3,     3,     0,    -6,    -4,    -3,    -6,    -2,    -2,     4,    -4,    -5,     1,     0,     1,    -7,    -5,    -2,    -5,     0,     4,    -3,    -1,     1,     3,   -10,    -9,    -2,     3,     4,     3,    -4,     0,    -8,    -4,    -6,    -6,    -1,    -7,    -4,     1,    -1,     1,    -4,    -5,    -6,    -3,     5,     3,    -1,    -4,     0,    -3,   -13,    -4,    -1,     5,     2,     0,     4,     4,    -1,    -3,    -4,     6,    -2,    -4,    -4,     0,     0,    -3,    -2,    -9,    -7,     0,     6,     3,    -8,    -6,     0,    -3,    -6,    -5,     1,    -1,    -1,    -1,     5,     8,     3,    -1,     2,     1,    -2,    -4,     3,     0,     0,    -1,    -6,   -10,    -4,     5,     3,     2,    -2,     2,     6,    -1,    -2,     3,    -1,     2,    -4,     4,     3,     2,     4,     5,     2,    -1,     1,    -3,    -1,     1,     0,    -1,    -5,    -8,     0,     8,     4,    -1,     0,    -1,     8,     1,    -4,     5,    -2,     0,    -2,     3,     1,     1,     3,     6,     3,     0,     2,    -6,    -8,    -1,    -1,    -1,    -4,    -3,     4,     9,    -1,    -2,    -7,     4,     7,    -1,    -4,     7,    -1,    -2,     0,    -1,    -1,     2,     6,     4,     1,     1,     0,    -8,    -7,     1,     0,     0,    -3,     0,    -3,     4,     2,    -4,    -4,     0,     3,     1,    -1,     1,    -1,    -2,    -4,     2,    -3,    -4,     5,     5,     1,     7,     6,    -3,    -6,     1,     0,     1,    -5,     0,    -2,     2,     4,     0,    -5,     1,    -1,     5,     2,     3,    -5,    -2,    -5,    -1,     2,    -2,     6,     2,     5,     4,     8,    -4,    -7,    -1,     0,    -1,    -5,     3,    -7,    -5,     2,    -1,    -3,    -4,     1,     4,     3,     5,     4,     1,     0,    -3,     2,    -4,    -2,    -5,     4,     2,     5,    -2,    -1,     1,    -2,     0,    -5,     2,    -3,    -5,     0,    -7,    -3,    -2,     0,    -3,     1,     7,     7,     2,     1,     5,    -1,    -2,    -2,     2,     4,     5,     7,     0,     1,    -1,     0,     0,     0,     0,    -2,     1,     0,    -6,    -7,    -1,    -5,    -8,    -6,     5,     5,    -2,     2,    -1,     1,     3,    -4,     4,     7,     3,     1,     2,     0,     1,     1,    -1,    -2,    -2,    -3,     3,    -8,   -15,   -15,    -1,    -4,    -4,    -4,    -5,    -3,    -8,    -5,     3,    -5,    -5,    -5,     2,    -2,   -12,    -8,     2,    -1,    -1,    -1,    -1,     0,    -4,     0,    -4,    -5,    -6,    -3,     7,     2,   -11,    -9,   -10,   -11,   -11,   -13,   -12,    -3,    -3,    -8,    -7,    -9,   -11,    -4,    -4,     0,     1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -4,     0,    -3,    -6,   -10,    -7,    -4,    -6,    -7,   -12,    -5,    -5,    -2,    -4,    -6,    -4,     0,     0,     0,     0,     1,    -1,     0,     1,    -1,    -2,     1,    -2,    -1,     2,     3,     1,     0,    -1,     0,    -2,     0,    -3,    -6,    -4,    -4,    -6,     0,    -1,     0,     0,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,     0,     1,     0,    -1,    -1,    -2,    -1,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,     1,     0,     0,    -1,     0,     1,     0,     1,     1,     0,     0,     1,    -1,     0,    -1,     1,     0,    -1,     1,     0),
		     7 => (    0,     0,    -1,     0,     1,    -1,    -1,     1,     0,     1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     1,     1,     0,    -1,     0,     1,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     1,    -2,    -3,    -1,    -3,    -3,    -3,    -5,    -6,    -3,    -1,    -1,     1,     2,    -1,     1,     0,    -1,     0,     0,    -1,     1,    -1,    -1,    -1,     0,    -2,    -3,    -1,    -6,   -10,    -5,    -3,    -2,    -2,    -3,    -1,     0,     0,    -2,    -1,    -1,     2,     1,    -1,     1,     0,     1,     0,     0,    -1,     0,    -4,    -6,    -5,    -6,    -1,    -1,    -4,    -7,    -9,    -5,    -4,    -4,    -2,     0,    -3,    -2,    -1,    -3,    -2,     0,     0,     1,    -1,     1,     0,    -1,     0,    -2,    -2,    -3,    -8,   -10,    -5,   -10,    -3,     1,    -1,    -5,    -8,    -9,   -10,    -7,    -5,    -4,    -3,    -7,    -9,    -7,    -6,    -4,     0,     0,    -1,     0,    -8,    -2,     5,     8,     5,     8,     2,    -4,     1,     1,     2,     4,     3,     1,    -1,    -6,    -8,   -12,    -8,    -7,   -11,   -17,   -12,    -3,     1,    -1,     1,    -2,    -5,    -1,     4,     4,     4,     2,     0,     4,     0,     6,     3,     3,    -3,    -5,    -3,    -6,     0,     0,    -2,    -7,    -6,   -13,    -7,    -7,    -2,    -1,     3,     0,     2,     2,     4,     2,     0,     0,    -4,     1,    -4,     3,    -2,    -4,    -7,    -3,    -4,    -6,    -6,    -1,    -5,     1,     2,    -2,    -7,    -8,    -3,    -4,     7,     4,     1,     6,     8,     0,     4,     1,     3,     1,    -5,    -3,    -2,    -3,     3,     2,     1,    -1,    -1,     0,     0,    -1,    -3,     0,   -11,   -10,    -4,     0,     5,     1,     4,     6,     8,     2,     2,     9,     3,    -4,    -5,    -4,     0,    -1,     2,    -3,     0,     3,    -1,     3,     3,     3,    -3,    -4,     0,     8,    10,     1,    -1,     1,    -2,     3,    -1,     4,     5,     5,     0,     0,     1,    -3,    -1,    -2,    -1,    -1,     3,     5,     2,     4,     3,     2,    -1,     0,     5,     3,     9,     0,    -3,     2,     5,    -1,    -2,     6,    10,     6,     5,     0,     0,     0,     1,     1,    -1,    -3,     6,    -3,     6,     3,    -2,    -4,    -5,    -2,    -7,    -2,     7,     0,     1,     1,    -3,    -6,   -10,     0,     0,     1,     0,    -4,    -3,    -3,    -7,    -4,    -1,    -3,    -5,     1,     0,     0,    -1,    -3,    -2,    -1,     1,     5,     8,    -1,     2,     5,    -6,    -7,    -8,    -3,    -3,    -6,    -7,    -8,    -8,   -12,   -13,    -2,    -1,     0,    -2,     5,     2,     3,    -2,     2,     7,     3,     3,    -6,    -5,    -2,    -2,    -2,    -6,    -5,    -8,    -6,    -8,   -13,   -11,    -9,    -9,   -11,    -6,     1,     1,     3,    -1,     3,     5,     6,    -3,     1,    -1,    -4,    -9,    -7,    -1,     0,     0,    -3,    -1,    -9,    -4,    -4,   -11,    -6,    -4,    -1,    -1,     2,     0,     4,     4,    -2,     2,     2,    -2,     7,     1,     4,    -2,    -2,   -11,    -5,    -2,    -1,    -2,    -2,    -2,    -6,    -5,    -6,    -8,     0,     5,     5,     4,     5,     3,     3,    -4,    -3,     0,    -1,     2,     0,     2,     3,    -4,   -13,   -12,    -5,    -3,    -1,    -1,     0,    -4,    -4,    -5,    -7,    -9,     0,     1,    -5,     0,     0,     2,     2,    -4,    -3,    -6,     2,     3,     1,    -2,     2,    -3,    -5,     1,    -1,    -2,     2,    -1,     6,    -3,    -6,   -10,   -11,    -7,    -4,   -11,    -8,    -1,     6,     6,    -6,    -6,    -5,    -2,    -1,    -5,    -4,    -6,    -3,    -5,    -5,    -3,     4,    -2,    -1,     2,     1,    -2,    -5,   -12,    -6,    -7,    -6,     2,    -4,    -3,     0,    -2,    -4,    -3,    -1,    -6,    -4,    -3,    -3,    -5,    -4,    -6,   -10,    -1,    -5,     0,     1,    -2,     0,    -2,    -7,    -1,     1,     3,    -3,    -1,    -1,    -1,     1,     2,    -6,    -7,    -5,    -9,    -8,    -6,    -2,     0,     2,     0,    -4,    -2,    -8,    -1,    -2,    -1,     0,    -7,    -5,     5,     6,    -3,     2,     0,    -2,    -4,    -2,     2,   -12,    -8,   -11,   -12,    -7,    -8,    -6,    -1,    -2,    -6,    -5,    -1,    -2,    -2,    -3,    -2,    -2,   -11,     4,     6,     5,     6,     8,     2,     2,     0,    -3,    -5,    -8,    -7,    -8,    -6,    -9,    -7,    -7,     1,     2,   -12,    -7,    -1,    -2,     0,     0,     1,    -3,   -12,     3,    -1,     4,    10,     1,     0,    -2,     3,    -4,    -3,    -8,    -3,    -9,   -14,   -11,   -10,   -10,    -1,     0,    -5,    -4,    -1,    -6,     0,    -1,     0,     3,    -1,     5,     8,     5,     2,     6,     1,    -2,     2,    -2,     3,    -5,    -4,   -12,   -13,   -10,    -6,    -9,     1,    -2,    -9,    -1,    -4,    -1,     1,    -1,     0,    -2,     5,    -5,     1,     0,     2,    -3,    -6,    -1,     3,    -1,    -7,    -9,    -7,    -8,    -5,    -3,    -4,   -11,    -1,    -2,    -7,     1,     0,    -1,    -1,     1,     1,    -1,    -6,    -7,    -7,    -2,     4,     6,     2,    -3,     0,     2,     4,    -4,    -2,     0,    -3,     1,     0,    -3,     3,     5,     2,    -2,     0,     1,    -1,     0,     0,     0,     1,     5,     5,    -1,    -1,    -1,     0,     3,     2,    -2,     7,     5,     0,     2,     1,     1,    -1,     1,     6,     4,     5,     0,     1,     0,     0),
		     8 => (   -1,     0,     0,     0,    -1,     1,    -1,     0,     1,    -1,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     1,    -1,    -1,     1,     0,     1,     1,    -1,     1,     1,     0,     0,     0,    -1,    -1,    -1,    -3,    -3,    -2,     1,    -1,     0,     1,     1,     0,     1,     1,    -1,     0,    -1,    -1,     1,    -1,     1,     0,     0,    -1,    -4,    -9,    -8,    -2,    -2,    -1,    -4,    -5,     4,     6,     2,    -4,    -4,    -4,    -4,    -1,    -2,     1,     0,     0,    -1,    -3,    -3,    -2,    -4,    -2,    -7,     5,     4,    -2,    -6,    -5,    -4,    -4,     1,     1,     1,     8,     4,     0,    -3,     5,     7,     0,    -2,    -3,     1,     0,    -1,    -3,    -4,    -7,    -9,     0,     4,    -1,    -5,    -5,     3,    -2,     0,     2,     2,     2,     1,    -1,     0,    -3,     0,     3,    -3,    -6,     4,     5,     0,    -1,    -1,    -2,    -4,    -4,    -7,     0,     0,    -7,    -4,    -2,     0,    -1,     3,    -1,     2,    -2,    -7,    -8,     5,    -1,     5,     0,    -2,    -2,    -1,    -2,    -2,     1,     0,    -4,    -7,    -5,     1,    -1,    -3,    -6,    -2,     1,    -3,    -2,    -2,    -6,     0,    -4,    -4,    -4,     2,     0,    -2,    -2,    -5,    -5,    -3,    -1,    -1,     1,    -5,    -2,    -3,    -1,    -1,    -3,    -3,    -1,    -1,    -4,    -1,    -3,    -7,    -4,     2,    -1,    -5,    -3,     1,     0,    -1,    -5,    -4,    -4,     0,     2,     4,    -2,    -4,    -1,    -1,    -3,     0,    -5,    -2,     1,     2,    -6,    -5,    -3,    -1,    -3,    -2,    -4,    -5,    -3,     1,     1,     2,    -7,    -8,    -2,     0,     8,     4,     0,    -2,    -4,     1,    -2,    -2,    -4,     2,     0,    -3,    -6,    -1,    -2,    -4,    -6,    -5,    -3,    -3,    -6,     3,     1,    -7,    -7,    -6,    -5,     0,     3,    -4,     1,    -2,    -3,     0,    -2,     1,    -3,    -3,    -1,     0,     3,     8,    -2,    -3,     2,     1,     1,     1,     2,     3,     0,    -2,    -5,    -8,    -3,    -4,     1,     2,     0,    -2,    -2,    -4,    -3,     3,     2,     0,     2,     5,     3,     1,    -3,    -5,    -2,    -1,     2,    -1,     0,    -5,    -5,     5,    -3,    -3,    -2,   -10,    -1,    -5,    -1,     0,    -4,     0,     4,     5,     3,    -1,     1,     4,     3,    -5,    -3,    -5,    -4,    -6,    -3,    -2,     0,    -5,    -1,     3,     3,     4,     1,    -9,    -9,    -7,     1,    -1,    -5,    -7,     1,     3,    -2,    -7,     3,    10,     4,     3,    -1,    -3,    -5,     0,     0,    -8,    -2,     0,     3,     6,     4,     4,    -1,    -8,   -12,     2,     0,     0,     0,    -9,    -4,    -1,    -3,    -7,     1,     1,    -1,     0,     1,     0,    -3,    -3,   -11,    -5,     3,     5,     5,     4,    -2,    -7,   -10,    -7,   -11,     0,    -1,     0,    -2,     2,     1,    -5,    -4,    -3,     0,    -1,     3,     4,     0,    -1,    -4,    -9,    -3,    -2,    -4,     1,    -2,    -6,    -7,    -4,    -3,     0,    -6,    -5,     0,    -1,    -1,     5,    -1,    -4,    -4,    -4,   -10,    -7,    -2,     3,     3,    -4,    -3,    -2,     0,    -1,    -1,    -4,    -1,     1,    -3,    -1,     1,    -1,    -6,    -3,     0,    -1,    -2,     3,    -3,    -4,    -6,    -3,    -9,   -16,    -6,     2,     5,    -1,    -1,     1,     1,    -3,    -6,    -6,     1,    -3,    -3,    -3,    -2,    -1,     1,    -2,    -1,     0,    -3,    -3,    -2,    -3,    -5,    -5,    -3,    -5,     0,     0,     3,     2,    -3,     3,     2,    -2,    -2,    -2,     0,    -4,    -2,    -4,    -2,    -1,    -1,    -3,     1,    -1,    -2,    -2,    -1,    -3,    -6,    -8,     2,     2,     0,    -2,     3,     2,    -1,     4,    -4,    -1,     0,     0,    -4,    -4,    -3,    -3,     0,     0,    -4,    -4,     1,    -1,    -2,     0,    -3,    -2,    -7,    -8,    -2,     2,    -2,    -2,    -1,     2,    -4,     1,    -6,    -6,    -2,     0,    -7,    -3,    -1,     0,     0,     0,    -3,     0,    -2,    -1,    -2,     0,    -3,    -4,    -6,    -1,    -5,    -4,    -2,     2,     7,     2,     2,     1,    -3,    -3,    -2,    -2,    -4,    -3,    -2,    -2,    -3,    -1,    -4,    -1,    -2,    -3,    -1,    -2,    -3,    -8,    -9,    -5,    -3,    -3,    -7,    -3,     4,     3,     3,    -5,    -1,     0,     0,     0,    -2,     0,     0,     0,    -2,    -1,    -3,     0,    -1,     0,    -3,    -1,    -1,    -4,    -8,   -10,    -3,    -1,    -4,     0,    -4,    -2,    -5,    -2,     1,    -4,    -3,     0,     2,     2,     1,    -1,     0,     0,    -4,     0,     1,    -1,    -1,    -1,    -2,    -3,    -3,    -5,    -4,    -3,    -9,    -3,    -4,    -4,    -2,     3,     3,    -3,     4,     2,     0,    -1,    -2,    -2,    -7,    -5,    -2,     1,     0,     1,    -2,    -1,    -2,    -4,    -3,    -2,    -3,    -3,    -5,    -6,    -1,     2,    -1,     3,    -1,    -1,     3,     2,     1,    -5,    -2,    -2,     0,    -2,    -1,     1,     0,    -1,    -1,    -2,    -1,    -3,    -5,    -2,    -1,    -2,    -4,    -8,    -9,    -7,    -8,   -11,     0,    -1,    -1,    -9,    -8,    -5,    -3,     1,    -1,    -1,     1,    -1,     0,    -1,    -1,     0,    -2,    -1,    -2,    -1,     0,    -2,    -1,    -3,     1,    -2,     0,     0,     0,     1,     0,     0,     0,     1,    -1,    -1,     1,     1,     0,     1),
		     9 => (    0,    -1,     1,    -1,    -1,    -1,    -1,     1,     1,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,    -1,     1,     0,    -1,     1,     1,     1,    -1,     0,     0,     1,    -1,     1,     1,    -1,     1,    -1,    -1,     1,     0,    -1,    -1,    -3,    -2,     0,     0,    -1,    -1,    -2,     1,     0,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     1,    -1,     1,     1,     0,     0,    -1,    -1,    -2,     0,     0,    -1,    -3,    -1,    -2,     0,    -1,     0,    -3,     1,    -1,    -2,    -1,     1,     0,    -1,     0,     0,     1,    -2,     0,    -2,    -1,     0,    -4,    -2,    -2,    -6,    -3,    -1,    -3,    -3,    -3,    -2,     3,    -2,    -3,    -4,    -3,     0,    -2,    -1,     0,    -1,     0,    -1,     0,    -2,    -2,     1,    -5,    -1,    -1,    -1,    -2,    -3,    -7,   -10,   -11,   -11,    -6,    -1,     4,    -5,    -8,    -6,    -4,    -4,    -3,    -7,    -5,     1,     0,     1,    -1,    -2,     0,    -1,    -2,    -3,    -7,    -4,    -6,    -2,    -2,     2,    -3,    -4,    -9,    -9,    -9,    -8,     1,    -4,    -5,    -6,    -4,    -3,    -8,     1,    -1,    -2,     0,    -2,     2,    -3,    -1,    -8,    -6,    -6,    -8,    -3,    -4,    -6,    -2,    -2,    -2,    -6,     0,    -4,     2,     4,     0,    -2,    -3,    -4,    -5,    -5,    -1,    -2,    -3,    -3,    -4,    -7,    -7,    -9,   -10,   -14,   -11,    -9,    -4,    -4,    -5,    -8,     3,     2,    -1,    -1,    10,     4,     4,     3,    -2,    -5,    -2,    -3,    -4,    -1,     1,     0,    -5,    -4,    -5,    -6,    -8,   -11,    -4,    -7,    -3,    -1,    -7,    -3,     1,     4,     4,     0,     1,    -1,     0,     4,     2,    -3,    -5,    -2,    -1,    -2,     6,    -1,    -3,    -4,    -3,    -1,    -8,    -2,    -2,    -3,    -3,    -7,     1,     5,     1,     0,    -1,     3,    -4,     1,     2,     0,     4,     3,   -10,    -5,     0,    -2,    -4,    -4,    -1,    -3,    -6,    -7,    -3,     0,    -1,     2,    -3,     2,    -1,    -5,    -5,    -4,    -9,    -8,    -4,    -2,    -3,    -1,     6,    12,    -4,    -7,     1,   -10,    -2,    -2,    -3,    -5,    -4,    -1,     6,     3,     4,    -1,     1,    -2,    -5,    -9,   -10,   -11,    -5,    -2,     3,    -1,     3,     1,     8,    11,    -1,    -6,     0,    -1,     1,    -6,     3,    -3,    -5,    -1,     3,     1,     5,    -2,    -7,    -5,    -8,    -6,    -3,    -9,     0,     0,     5,    -2,     4,     5,    -2,    -9,    -7,    -7,    -1,    -2,    -3,    -4,     3,    -4,     0,     2,     1,     3,     6,     1,     1,     1,    -4,     3,     6,     0,     0,     7,     2,     7,     1,    -3,    -6,    -4,    -4,     1,     0,    -2,     0,    -4,     3,    -4,     0,    -3,     6,     7,     6,     0,     3,     3,     3,     4,     1,     1,     0,     3,    -2,    -7,    -3,    -9,    -8,    -2,     1,     0,    -1,     1,    -7,    -5,     3,    -4,    -5,    -4,     1,    -3,     1,     3,     3,     7,     0,     2,    -1,     0,     4,     2,    -6,    -7,   -10,    -7,    -6,    -1,     6,    -1,    -1,    -2,    -5,    -4,     2,    -2,    -1,     0,    -3,    -2,     2,     2,    -2,     1,    -5,    -6,     0,     3,     1,    -1,    -8,    -3,    -3,    -9,    -4,     0,    -1,     0,     1,    -1,    -4,    -1,    -3,    -4,    -3,     4,    -4,    -6,    -4,    -3,    -2,    -1,    -3,    -1,     0,     4,     3,    -3,    -4,    -2,    -4,    -9,    -4,     5,    -1,    -2,     0,     1,    -4,    -2,    -8,    -6,     0,     3,    -4,    -7,    -1,     2,    -3,    -2,     3,    -3,    -1,    -2,     2,     0,    -4,    -3,    -1,    -3,    -2,     6,    -3,    -3,     0,    -1,    -5,    -3,    -9,    -7,    -3,    -3,    -5,    -8,    -5,    -7,    -1,    -4,    -1,    -4,    -5,    -3,    -1,     0,    -8,    -4,    -1,    -2,     2,     7,    -4,    -3,     1,     0,     3,    -2,    -6,    -4,   -11,    -9,     3,    -3,    -7,    -1,     4,     3,    -2,    -5,    -2,    -1,     0,    -2,    -5,    -4,    -3,    -1,     2,     6,    -1,    -1,     0,    -1,    -1,    -3,    -7,    -3,    -8,    -6,     2,     3,     0,    -3,    -1,    -4,    -3,    -9,     0,    -2,    -2,     2,    -4,    -3,    -5,    -2,     1,     5,    -5,     0,     1,     1,    -4,    -6,    -8,    -6,   -10,    -3,     2,     3,     4,     3,    -1,    -4,    -7,    -5,    -3,    -2,    -7,     0,     1,    -4,    -2,     0,     2,    -1,    -3,    -1,     0,     1,    -4,    -5,   -10,    -5,    -6,     1,     6,     4,     1,    -4,    -1,    -6,    -6,    -2,     0,    -1,    -1,    -1,     1,     0,     1,    -4,    -1,     2,    -3,     1,     1,     1,    -2,    -3,    -5,     0,     0,     3,     1,     4,     1,    -1,     0,    -6,     1,    -4,    -4,     0,    -3,     2,     1,     0,     2,     0,    -1,    -1,    -2,     0,    -1,     1,     4,    -2,     2,    -1,    -2,     0,     2,     1,     4,     0,     3,     0,    -4,    -4,     1,     5,     3,     1,    -2,    -2,    -3,     3,     1,    -1,    -1,     0,     1,     1,     0,     7,     3,    -1,     4,     3,    -3,     0,     2,     6,     1,     5,     4,     2,     7,     9,     5,     3,     7,     1,    -3,     2,    -1,     0,     0,    -1,    -1,     1,     1,    -1,    -2,    -1,     2,     7,     6,     4,     4,     8,     4,     4,     3,     3,     2,     3,     5,     6,    -2,    -3,    -2,    -2,     1,     0,    -1,     0),
		    10 => (    1,     1,     0,    -1,     0,     0,    -1,     0,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     1,    -1,     0,     0,     1,     0,    -1,    -1,    -1,     1,     1,    -1,     1,     1,    -1,    -1,     1,     3,     0,    -2,     4,     5,     6,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,     1,     1,     1,    -2,     5,     4,    -1,    -1,     1,    -2,    -2,    -4,     0,     0,    -3,    -1,    -6,    -1,    -7,    -6,    -6,    -5,    -2,    -6,    -4,    -3,    -1,    -1,     1,     1,     1,     1,     0,    -1,     0,    -2,     0,     2,    -4,   -10,    -6,     0,     1,    -1,    -5,    -4,    -8,    -1,     0,     1,    -5,    -5,    -3,    -1,     1,    -9,     0,     1,     1,    -1,    -2,     1,    -6,    -4,    -5,    -3,    -7,    -7,    -6,   -10,   -10,    -2,     2,    -5,     1,    -2,     0,    -1,     0,     2,     1,    -4,    -7,    -7,    -1,    -1,    -1,    -3,    -1,     1,    -7,    -4,    -7,    -2,     0,    -9,    -4,    -6,    -4,    -1,    -1,    -3,     0,    -3,    -1,    -9,    -4,     4,     0,    -7,    -5,    -6,    -4,     0,     1,    -5,    -1,    -1,    -1,    -3,    -3,     1,    -1,    -3,     0,    -3,     0,     0,    -3,    -2,     0,     1,     1,    -4,     3,     5,    -3,    -7,    -7,     0,    -1,     0,    -6,    -3,    -2,    -1,     1,    -1,    -5,    -1,    -2,    -1,     1,    -1,    -3,    -2,     1,    -3,     1,     3,     1,    -7,     0,    -2,    -3,   -10,    -7,    -5,     3,    11,    -8,     4,     2,    -1,    -2,    -2,    -6,    -3,    -3,     0,     0,     2,   -10,     2,     4,     0,     6,     4,    -5,    -7,    -2,    -3,    -3,   -10,    -4,    -8,    -1,     1,    -2,     6,    -1,    -1,     1,    -4,     1,     2,    -2,     1,    -1,     0,     0,    -3,    -3,     4,     2,     4,    -2,     4,    -2,    -4,    -4,    -4,    -9,    -8,     0,     0,     1,     4,     2,    -1,    -1,    -1,    -2,    -2,    -1,     1,    -1,     0,    -2,     1,    -8,    -3,     3,     0,     0,    -2,    -4,     1,    -1,    -6,    -6,    -7,    -1,    -1,    13,    -4,    -4,    -5,     1,     2,    -4,    -8,    -7,    -1,     1,    -2,     2,    -5,    -9,    -7,    -1,     2,     3,     0,    -7,    -8,    -6,    -8,    -7,    -4,     1,     0,     2,    -2,    -5,     5,     5,     1,    -3,   -11,    -1,     2,     1,     4,    -1,    -7,   -10,    -4,     1,     4,     6,     2,    -6,    -7,    -3,    -6,    -8,    -3,    -1,    -1,     3,     3,    -5,     9,     4,     3,     1,    -4,     4,     2,    -1,     1,    -5,   -12,   -16,    -6,     0,     1,     6,     8,    -5,    -3,     3,     1,    -1,    -5,    -2,     1,     1,    -1,    -6,     0,     5,    -4,     1,     3,     3,     1,     7,     5,    -1,    -9,    -7,    -5,    -4,     3,     8,     7,    -5,     0,     5,     0,    -3,    -3,    -2,     1,    -1,    -4,    -8,    -5,    -3,    -3,    -1,     2,     1,     3,     6,    12,    -5,   -12,    -6,    -2,     0,     7,    -2,     3,    -7,    -1,     3,    -2,    -2,   -10,    -2,     1,     1,    -4,    -4,    -3,    -1,    -5,    -5,     4,    -1,    -2,     3,     4,    -9,   -13,    -1,     2,     2,     3,     2,    -5,    -9,    -6,    -2,    -4,    -6,    -8,     8,     1,    -2,    -4,    -5,    -1,    -4,    -7,    -2,     1,    -2,     0,     0,     2,    -7,    -7,    -1,     2,     2,    -2,     2,    -1,    -8,    -3,    -4,    -4,    -5,    -5,    13,     0,    -2,    -5,    -5,    -4,    -9,    -5,    -3,     0,    -2,     2,     1,    -5,    -6,    -4,     0,     6,     2,     1,    -3,    -4,    -5,     0,    -4,    -2,    -4,    -6,    -3,     0,     4,     0,    -3,    -5,    -5,    -8,    -3,     5,     1,     0,     1,    -1,     1,    -3,    -2,    -6,    -3,     4,    -2,    -2,     0,    -4,    -4,    -1,    -7,    -4,    -1,    -1,     4,    -2,    -4,    -1,    -5,    -9,    -4,     2,     1,     3,     4,     4,     3,    -1,    -8,    -6,    -1,    -4,     0,    -2,     2,    -4,    -1,    -5,     1,     3,     1,     1,     0,    -2,    -5,    -6,    -3,    -5,    -4,     0,     1,     7,     1,     6,     3,    -4,    -4,    -3,    -3,     1,     3,     0,    -3,    -5,    -1,     0,     1,    16,     4,     1,    -1,    -5,    -8,    -7,    -4,    -6,    -5,    -3,     4,     0,     0,     0,    -7,     1,     3,     3,    -4,    -7,    -1,    -6,    -5,    -4,    -2,    -1,     2,     9,     3,    -1,     1,    -1,    -5,    -6,   -10,    -4,    -3,    -4,     5,     9,     3,     2,    -2,    -1,    -4,     1,    -3,     0,    -1,    -6,    -5,    -1,    -2,     0,     0,    -7,     0,    -1,     0,    -2,     0,     3,     2,    -7,    -9,    -9,    -7,    -6,    -4,    -1,    -5,    -6,    -4,    -4,    -2,     3,    -8,    -5,    -4,    -3,    -1,     1,     1,     1,     1,     1,     0,    -2,     0,    -5,    -4,    -5,    -7,    -2,    -4,    -9,   -11,   -18,   -17,   -18,   -14,    -8,    -7,    -7,    -6,    -8,    -6,    -3,    -3,     0,     0,     0,     0,     1,    -1,     1,     1,    -3,    -5,   -11,    -3,    -4,    -9,    -6,    -6,    -4,    -5,    -2,    -6,    -6,    -6,    -8,    -7,    -6,    -5,    -3,    -3,     0,     1,     1,     0,     0,    -1,    -1,     1,     0,     1,    -1,    -2,    -3,     0,    -1,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,     1,    -1,     0,    -1,     1,    -1,    -1,     0),
		    11 => (    0,     0,    -1,    -1,     1,    -1,     1,     1,     0,     1,     1,    -1,    -1,    -1,     1,    -1,     0,     1,    -1,     0,     0,    -1,     0,    -1,     1,     0,     1,    -1,     0,     0,    -1,     1,     0,    -1,     0,     1,     1,     0,     0,    -1,    -1,    -2,     0,    -2,    -2,    -2,     0,    -1,     0,    -1,    -1,     1,    -1,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,    -2,    -1,     2,     1,     0,    -1,    -1,    -4,    -9,   -11,    -9,     2,     3,    -4,    -2,    -3,    -1,    -1,     0,     0,     1,    -1,     3,     1,    -1,    -1,    -1,     4,     4,     5,     4,     1,     1,     0,     1,    -6,    -9,    -7,    -1,    -3,    -3,    -5,     1,     4,    -4,     0,     0,     1,    -1,     1,     3,     3,     1,     3,     4,     3,    -1,     0,    -3,    -3,    -3,    -3,    -4,    -7,    -6,    -3,     1,     2,     5,     0,     0,    -2,    -6,    -4,    -6,    -5,     0,    -1,     0,     5,     4,     4,    -1,     0,    -6,    -4,    -5,    -6,    -3,    -2,   -11,   -12,    -8,     1,     2,     1,     0,     5,     4,     2,     1,    -4,    -5,     0,     0,     0,    -1,     5,     9,    -1,    -3,    -1,    -7,     5,     4,     0,   -11,   -13,   -16,   -13,    -6,    -4,     0,    -1,    -2,     1,     0,     1,    -3,    -5,    -4,    -2,     1,    -2,    -3,     0,    -4,    -4,    -3,    -4,    -8,     0,     5,     0,    -7,   -10,   -11,    -9,    -3,    -2,     3,     0,     1,    -1,    -1,     1,    -7,   -10,    -6,    -2,     0,    -4,    -3,    -1,    -2,    -2,    -3,    -5,    -5,    -2,     1,    -7,    -5,    -6,   -11,    -5,     0,     2,     1,     0,     2,    -2,     0,    -1,    -7,    -8,    -6,    -2,    -1,     0,    -3,    -1,    -2,    -3,    -2,    -2,    -2,     0,    -9,   -10,   -11,   -18,   -15,     0,     4,     1,     2,    -1,    -1,    -2,     0,     0,    -2,    -5,    -2,    -4,    -1,     0,    -2,    -1,     0,     0,    -6,    -6,    -8,    -5,    -9,    -9,   -12,   -15,    -7,    -1,     7,     1,    -2,    -1,     0,     2,     2,    -1,     1,    -2,    -3,    -2,    -1,     0,     1,     1,    -2,     1,    -3,    -7,    -7,    -6,    -8,    -5,    -7,    -5,    -4,     8,     3,     3,     8,    -2,     0,     1,    -5,    -7,    -4,     1,    -4,     1,    -1,     0,    -4,     2,     0,     2,     1,    -5,     1,    -9,    -6,    -6,    -2,    -4,     2,     6,     0,     3,     1,     2,    -6,     0,    -5,    -1,    -3,     0,    -2,     0,    -1,     0,    -3,     0,     0,    -3,    -1,    -3,    -2,    -5,    -2,    -1,    -4,     1,     6,     4,     1,     4,     3,    -3,   -14,    -6,    -6,    -2,    -3,    -1,     0,     0,    -1,     0,     0,     0,     2,    -2,    -2,     0,    -1,     4,     4,    -2,     0,     4,     2,     2,     3,    -5,    -7,   -16,   -17,    -2,     2,     0,    -1,    -3,    -2,    -1,     0,    -1,     3,     6,     0,    -7,     0,     1,     9,     3,     3,     1,    -1,     1,     1,     3,     1,    -5,   -14,   -18,   -10,    -2,     2,     0,   -11,    -8,    -5,     0,     1,     0,     1,    -2,     2,    -2,    -4,     0,     3,     3,    -5,     0,    -2,     0,    -4,     3,     3,    -1,   -10,   -10,    -1,     3,     3,     7,     9,    -4,    -6,    -2,     0,     0,     0,    -3,     0,    -7,    -3,     2,     0,     0,    -1,     4,     3,     0,     1,    -5,     1,    -1,     2,     4,     5,     8,    11,    10,     7,    -1,   -11,    -4,     0,     0,    -1,     0,    -5,   -12,    -7,     1,     1,    -1,    -2,     3,    -2,    -1,     0,    -1,    -4,     0,     2,     3,     3,    -1,     6,     5,     0,     2,    -1,     3,     0,     1,     1,    -4,    -7,    -2,     1,     2,     1,    -1,    -2,    -1,    -1,    -5,   -10,    -7,    -5,    -7,    -6,    -3,    -3,    -2,     4,     5,     5,     5,     0,     2,    -1,     0,     0,    -3,     2,     4,     3,     1,     2,     0,    -3,     3,    -3,    -7,    -7,    -5,     2,    -3,    -7,    -5,    -5,    -2,     4,     4,     7,     0,     1,     2,     3,     3,     0,     0,    -1,     0,    -1,     1,     1,    -2,    -2,    -1,    -3,    -1,    -2,     1,     4,     3,    -4,    -3,    -5,    -2,     1,     7,     6,     3,     1,     1,     4,     3,     0,     0,     1,     7,     2,     0,     2,     4,    -2,    -3,    -5,     0,    -5,     4,     5,     0,    -4,    -5,    -5,    -5,     1,     1,     1,     0,     1,     0,     0,     0,    -2,     3,     1,     0,     0,     0,     5,     3,    -2,    -5,     1,     2,     3,     4,     2,    -3,    -3,    -4,    -2,     0,    -1,    -1,     3,     6,     8,     1,     0,     0,     1,     2,    -6,    -4,    -6,    -8,    -1,     5,    -1,    -3,     4,     7,     1,     1,     0,     0,     0,    -2,     0,     1,     1,     1,    -4,     1,     0,     1,     0,     0,     1,    -3,    -5,    -5,    -2,   -10,    -3,     2,    -2,     2,     5,     2,    -8,    -5,    -4,    -7,    -4,    -2,    -1,    -4,    -3,    -2,    -3,    -1,     0,    -1,     0,    -1,     0,    -1,    -5,    -4,    -4,    -5,    -7,    -6,    -4,    -2,    -4,    -4,    -3,    -3,    -5,    -5,    -2,     0,    -1,    -1,     0,    -1,     1,     0,    -1,    -1,     1,     0,    -1,     1,     0,    -1,     0,     0,     1,    -1,    -4,    -2,    -1,    -1,    -2,    -1,     1,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,    -1,     1),
		    12 => (    1,    -1,     1,    -1,     0,     0,     0,     1,     0,     1,    -1,     1,     1,    -1,     2,     1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,    -4,    -2,    -2,    -2,    -2,    -3,    -1,     1,     1,     0,    -1,    -4,    -3,    -2,     0,     1,     0,     1,    -1,     0,     1,     0,    -2,    -4,    -3,     1,     0,    -1,     0,     1,     1,     4,     1,    -2,    -2,    -4,    -4,    -3,     1,     1,     1,     1,    -3,    -1,    -2,     1,     1,     1,     0,     1,    -1,    -7,     0,    -4,    -2,    -3,     0,     4,     7,     5,     4,     1,     0,     1,     0,     0,    -2,     0,     1,     1,    -4,    -6,    -3,    -3,    -1,     1,     0,     0,     0,    -3,     1,     2,     5,     6,     1,     0,     2,     6,     5,     6,     0,    -1,     0,    -3,    -1,    -4,    -2,    -3,    -4,    -4,    -7,    -6,    -5,    -1,     1,     1,    -4,    -1,     0,     2,     5,     8,     4,     2,     2,     1,     1,     1,    -3,    -2,    -3,    -2,    -3,    -1,     0,     1,    -2,    -3,    -6,    -3,    -3,    -1,    -1,    -1,     0,     0,    -1,     0,     6,     5,     3,     3,     1,     0,    -2,     0,    -2,    -3,    -2,    -2,    -1,    -4,    -1,     2,     1,    -4,     0,     5,    -3,     0,     1,    -1,    -1,    -1,    -1,     1,     0,     2,     0,    -3,    -2,     0,    -2,    -3,    -1,     1,     1,    -4,    -4,    -4,     1,     3,    -1,    -4,     2,     7,    -9,    -4,    -4,     2,    -2,     0,    -1,     0,    -1,     1,    -4,    -5,    -3,    -3,    -1,     1,     0,     1,     1,    -1,    -3,    -1,    -1,     0,    -1,     2,     1,    -1,    -8,    -4,     1,    -3,     4,     0,    -2,    -1,    -3,    -2,    -4,    -5,    -2,    -3,     0,    -1,     4,     1,    -3,    -1,    -2,    -2,    -1,     2,     1,     0,    -2,    -4,     0,    -3,     1,    -1,     1,    -1,    -4,    -2,    -3,    -5,    -8,    -7,    -7,    -3,    -1,    -2,    -2,     0,    -4,    -1,    -5,    -1,    -4,     2,     3,    -2,    -5,    -2,     2,    -4,     0,    -3,    -1,    -4,    -3,    -2,     0,    -7,    -7,    -7,    -7,    -2,    -1,     1,     2,    -2,    -5,    -3,     1,    -1,    -2,    -2,    -1,    -2,    -3,    -2,     0,    -2,    -1,    -2,    -4,    -5,    -2,    -1,    -3,    -4,    -2,    -2,    -2,     1,     3,     0,    -1,    -1,    -3,    -2,    -3,     0,    -5,    -5,    -2,    -4,    -5,     0,     2,     1,     1,    -2,    -3,    -3,    -3,    -5,    -2,    -5,    -3,    -1,     0,    -1,     0,    -1,    -1,    -1,    -3,    -3,     1,     0,    -2,    -2,    -4,    -4,    -1,     2,     4,     0,     0,    -3,    -2,    -1,    -4,    -6,    -1,    -4,    -3,    -3,    -3,    -4,    -4,    -3,    -2,    -3,    -4,    -5,     0,    -1,    -1,    -5,    -4,    -4,    -1,     3,     5,     3,     0,    -4,    -2,     0,    -3,     1,    -3,    -2,     0,    -3,    -2,    -2,    -4,     0,    -1,    -4,    -7,    -5,     0,     0,     0,    -2,    -4,    -5,     2,     5,     7,     5,     0,    -2,    -1,     4,     3,     0,    -2,    -2,    -1,    -1,     1,     0,     1,     1,     1,    -3,    -4,    -4,    -4,    -3,    -2,    -1,    -3,    -4,     1,     4,     8,     5,    -1,    -1,     1,     4,     3,    -1,     0,    -4,    -2,    -1,    -2,    -2,     3,     1,    -2,    -2,    -5,    -5,    -3,    -4,    -5,    -3,    -3,    -6,     0,     6,     5,     6,     1,     0,    -1,     1,     4,     0,    -4,    -2,     0,     1,    -1,    -3,     0,    -1,     0,    -1,    -5,    -2,    -4,    -4,    -2,    -2,     1,     0,     4,     4,     4,     5,     0,     0,     0,     2,     1,    -2,    -1,    -2,    -1,    -2,     1,     1,     0,     0,    -3,    -2,     0,    -1,     3,    -6,    -2,     2,     3,     5,     5,     5,     9,     9,     0,    -2,     1,    -1,     2,     2,    -1,    -1,    -2,     0,     0,     3,     0,    -2,    -3,    -3,    -2,    -2,     2,    -4,    -1,     2,     4,     5,     6,     3,     3,    -1,     1,     0,     2,     3,    -2,     1,     0,    -3,    -4,    -3,    -3,    -1,    -3,    -2,    -3,    -2,    -1,     1,    -1,    -2,     1,     3,     6,     5,     3,    -1,     1,    -2,     0,     1,     1,     2,     3,    -2,    -1,    -2,    -1,    -2,    -4,    -2,    -1,    -1,     2,    -2,     2,    -2,    -3,     0,     1,     2,     5,     5,     1,     4,    -4,    -2,     0,     0,     1,     1,     1,     0,    -1,     0,     2,    -2,    -1,     2,     0,     1,     2,     1,     0,    -4,    -5,    -3,     1,     2,     5,     6,     0,     3,    -2,     1,     0,     1,    -3,    -1,    -3,    -3,    -3,     0,    -1,    -1,    -3,     0,     3,     0,     3,     0,    -4,    -2,    -3,     0,    -3,    -1,    -3,     2,     2,     1,     0,     0,    -1,     0,    -5,    -1,    -1,    -1,     0,    -1,    -3,    -4,    -4,    -1,    -4,    -7,    -3,    -3,    -5,    -1,    -3,     0,    -3,    -3,    -4,    -2,    -2,    -1,     0,     1,     0,     1,     0,     1,    -2,    -4,    -3,    -3,    -4,    -6,    -5,    -2,    -2,    -3,    -6,    -5,   -10,   -11,    -9,    -7,    -4,    -3,    -5,    -3,     0,     0,     1,    -1,     1,     0,     1,     0,     0,     1,    -1,    -2,    -3,    -1,    -3,    -3,    -2,    -6,    -3,    -3,    -4,    -3,    -4,    -2,    -3,    -2,    -3,     1,     0,     0,    -1,     1),
		    13 => (   -1,    -1,     1,    -1,    -1,     0,    -1,    -1,     1,     0,     1,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,     1,     1,    -1,    -1,     1,     0,     0,     0,     1,     0,    -1,     1,     0,    -1,    -1,     0,     1,     0,    -1,     1,     0,    -1,    -2,    -1,    -2,    -1,     1,     0,    -1,     0,    -1,     1,    -1,    -1,     1,     0,     0,     1,     0,     0,     1,    -1,     1,     0,    -3,    -5,     4,     3,     5,    -2,    -2,    -3,    -1,     0,    -1,     0,    -3,    -2,    -4,    -2,     0,     0,     0,     1,     0,     1,    -1,     0,     0,    -2,     1,    -2,    -3,    -5,    -6,    -4,    -5,   -12,   -18,   -14,   -11,    -1,     2,     0,    -5,    -4,    -3,    -6,    -1,    -1,     0,    -1,     1,     3,     0,     2,    -4,    -6,    -3,    -3,     5,    -3,     3,     6,    -5,    -3,     0,    -2,    -5,     4,     1,    -5,    -2,     3,    -2,    -2,    -5,    -2,    -2,     0,     1,     0,     5,     0,     6,     8,     4,     3,    -3,    -5,     0,     0,    -1,    -2,     1,     0,    -3,    -2,    -1,    -1,    -7,    -6,    -3,    -6,    -2,    -5,    -3,    -1,     0,     0,     1,     2,     5,     6,     2,     0,    -2,     0,     0,     4,     0,     4,     2,     1,     0,     3,     0,   -12,    -1,    -4,    -8,    -4,    -2,    -2,     0,    -1,    -1,     1,     2,    -3,     7,    -3,     7,     2,     1,     4,     1,     2,     1,     2,     2,    -6,    -3,     0,     1,    -3,    -2,     0,    -8,    -5,    -3,    -3,    -4,    -1,     0,    -1,     2,    -3,     7,     1,     1,     2,     0,     8,     4,     2,    -2,    -1,    -3,     0,     0,     2,     3,    -2,    -5,     0,    -4,   -12,    -7,    -2,    -5,     1,     1,    -3,     4,     2,     5,     1,     8,     9,     4,     4,     0,    -7,    -5,    -1,     1,     3,     0,     1,     1,     3,     1,    -2,    -9,    -9,   -10,    -4,    -3,     0,     1,    -4,     5,     8,     6,     4,     4,     2,    -8,   -11,   -15,    -8,    -6,     2,     2,     5,    -1,     7,    -1,     1,     1,    -3,    -7,     0,    -5,    -4,    -3,     0,     1,    -3,     0,     7,     3,    -4,    -7,   -12,   -19,   -10,    -2,    -3,     3,     7,     1,    -1,    -4,    -3,     1,    -1,     2,     0,    -9,    -6,    -4,    -3,    -1,     0,    -1,    -1,     6,     7,    -4,   -10,   -16,   -10,   -10,     1,     6,     4,     5,     4,     1,    -3,    -6,    -5,    -5,   -10,    -6,   -13,    -6,   -10,    -4,     0,     0,    -2,    -1,     1,    -2,    -2,    -1,    -6,   -10,    -8,    -4,     0,     5,     2,     3,     2,     1,    -5,    -2,    -3,    -5,    -5,    -7,    -8,    -3,    -2,    -2,    -4,    -3,    -2,    -1,     2,     0,     3,     0,    -5,    -6,    -3,     6,     0,     2,    -1,     1,     0,     4,    -2,    -2,    -3,    -7,     2,    -5,    -4,    -5,     2,    -1,    -9,    -5,    -2,    -2,     2,     2,     5,    -3,    -4,    -2,    -1,    -1,     3,     5,     9,     0,     1,     1,     3,     0,    -5,    -6,     0,     0,     4,    -5,     6,    -1,    -5,    -2,    -3,     1,     1,     2,     5,    -6,    -7,    -4,    -3,     2,     6,     0,     0,     5,     4,     4,    -1,     0,    -1,     0,    -3,     1,     7,     3,     4,    -1,    -7,    -7,    -3,     1,     1,     2,     5,    -6,   -11,   -11,    -9,    -4,    -2,    -7,    -1,     1,     3,     0,     1,     3,     1,    -1,     1,    -2,     6,     6,     1,    -3,   -11,    -5,    -2,    -2,     0,     4,     9,    -2,    -6,    -9,   -11,   -18,   -24,   -20,   -21,   -20,   -15,   -10,   -13,    -3,     8,     1,     2,     3,     2,     9,     5,    -4,    -9,    -4,    -4,     0,    -1,    -7,     5,     4,     5,    -4,    -4,    -8,   -11,   -16,   -18,   -16,   -14,   -11,   -12,    -7,    -3,     1,     6,     5,     4,     6,     7,    -1,    -6,    -7,    -4,     1,     1,    -5,    -3,    -1,     5,     2,    -1,    -1,    -6,    -6,    -5,    -4,    -1,    -2,    -7,    -8,    -1,     0,     4,     3,    -1,     1,    13,    -1,    -6,     0,     0,    -1,     1,     3,     4,     3,     0,     4,     2,    -1,    -2,     1,     0,     2,     3,    -2,    -1,    -3,     0,     2,     1,     6,    -3,    -3,    -1,    -4,    -5,    -1,     1,     1,    -1,     5,     5,     7,     4,     2,     3,     6,     2,    -1,    -3,     0,     3,    -4,     0,    -1,    -4,     1,     1,     3,     2,     0,     2,    -8,    -6,     0,    -1,     0,     0,     5,     7,     6,    -1,     0,     3,     2,     1,    -1,     3,    -2,     2,    -2,    -2,    -3,    -3,    -6,     0,    -5,    -2,    -5,     0,    -6,    -1,     1,     1,     1,     1,     2,    -1,     8,     5,     2,     7,     5,     0,     5,     4,     2,    -1,     1,    -2,    -3,     1,    -1,    -5,    -8,     0,     3,     1,    -5,     0,     0,     0,     1,     0,    -1,    -4,     2,     6,     1,     3,     5,     3,    -1,    -3,    -4,    -5,    -7,    -4,    -1,    -8,    -8,    -8,    -6,    -5,    -3,   -14,    -6,    -1,    -1,     0,     1,     0,     1,    -3,     0,     0,    -4,    -2,    -6,    -7,    -7,    -8,    -7,     2,    -2,    -5,     5,     0,     1,    -1,    -1,     0,    -4,    -1,     0,    -1,     1,     0,     1,    -1,     0,    -1,    -1,     1,    -1,     1,     0,    -6,    -5,    -3,     0,    -4,    -3,    -3,    -2,     0,    -2,    -5,    -5,    -1,    -2,    -1,     0,    -1,    -1,     0),
		    14 => (    0,    -1,     1,    -1,     1,     1,     1,    -1,     0,    -1,     0,     0,    -3,    -2,     0,     0,     0,    -1,     0,    -1,     1,     0,    -1,     1,     1,     1,     1,     1,     0,     0,     1,     1,     0,     0,     0,    -2,    -1,    -2,    -4,    -3,    -5,    -3,    -1,   -10,    -9,    -7,    -2,    -1,    -4,    -2,    -1,    -1,    -1,     0,     0,     1,     1,    -1,     0,    -4,   -11,     0,    -1,    -3,    -6,    -4,    -9,    -8,    -9,     0,     2,     2,    -8,    -5,    -3,    -3,    -8,    -4,     1,    -1,    -1,    -5,     0,    -1,     0,     0,     0,    -4,   -10,    -8,    -4,    -2,    -2,    -3,    -8,    -8,    -6,     0,     3,     0,    -6,    -8,     0,     4,     5,     4,    -2,    -5,    -8,    -4,     0,     0,     1,     0,    -2,    -7,    -3,    -4,    -2,     2,     3,     5,     0,    -8,    -8,     1,     1,    -1,    -2,    -2,     3,    -1,     4,     1,    -1,    -4,    -8,    -5,    -6,    -1,     0,     1,    -3,    -1,    -3,     0,     3,     2,     5,     3,    -1,    -7,    -7,    -5,     0,    -3,    -5,     1,     1,     4,     0,    -1,     0,     0,    -2,     3,    -7,    -2,    -1,     0,    -5,    -2,     3,     4,     1,     1,     0,    -3,     1,    -3,     3,     2,     6,    12,    12,     9,     6,     5,     1,     6,    -3,    -1,    -2,    -4,     0,    -3,     0,    -9,    -2,     1,     2,     2,     6,     5,     0,     2,     2,    -1,     3,     3,     3,     8,     9,     7,     1,    -1,     0,     0,     1,     1,    -2,     1,    -1,    -9,    -4,   -11,    -1,     1,     0,     1,     6,     4,     5,    -1,    -5,    -1,    -3,     0,    -2,     1,     0,    -2,     0,     0,    -1,     1,    -1,     0,     2,     3,    -1,    -8,     0,    -5,    -6,     0,     0,     1,     0,    -1,    -1,    -8,    -8,    -1,    -4,    -7,    -8,    -4,    -3,    -3,     0,    -3,     0,     3,     1,     1,    -3,    -1,    -3,    -6,     0,    -4,     1,     0,    -3,    -2,    -4,    -3,    -4,    -5,    -3,    -3,    -4,   -10,   -11,    -7,    -6,    -4,     1,    -2,    -4,     4,    -2,    -8,   -10,    -6,    -3,    -2,     0,    -4,    -3,     0,    -4,     0,    -4,    -2,    -5,    -5,    -4,    -5,     0,    -4,    -9,    -1,    -3,     2,     1,     2,    -2,     2,    -4,   -12,   -11,    -7,    -5,    -8,    -1,     1,     1,     2,    -2,     2,     3,    -1,     3,     3,     3,     1,     4,     3,    -5,     3,     2,     0,     0,     2,     3,     9,     2,    -2,    -7,    -4,    -9,    -9,    -1,    -2,    -4,     0,     5,    -1,     0,    -1,     3,     2,     0,     4,     2,    -1,     2,     7,     3,     4,     4,     5,     3,     2,    -2,    -2,    -7,    -3,    -7,     0,    -1,    -2,   -10,    -2,     5,    -2,    -1,    -1,    -1,     0,    -4,    -1,    -5,    -2,     1,     7,     2,     5,     7,     5,     5,     1,     0,    -3,     1,    -4,     6,     1,     1,     0,     5,     1,     4,    -6,    -3,     0,    -2,    -4,   -10,    -6,    -3,     3,     5,     9,     9,     7,     7,    -1,     0,     2,     2,    -2,    -5,    -6,     6,    -5,     0,     0,     1,     3,     4,    -5,    -5,    -3,    -3,    -6,    -8,    -1,     2,     7,    11,     9,    10,     2,     7,    -2,     0,    -1,    -2,    -3,    -3,     1,     1,    -2,     1,     0,     3,    -2,     8,    -6,    -3,    -3,    -1,    -6,    -1,     3,     7,     7,     6,     7,    10,     3,     5,    -4,    -2,    -1,     1,     0,    -4,     1,     4,    -5,    -7,    -1,     0,    -1,     6,    -4,    -3,    -3,   -11,    -3,     2,     3,     6,     1,     6,     6,     7,     2,    -1,    -5,     1,     1,    -1,     7,    -6,    -7,    -2,    -1,     0,    -2,    -4,     5,     0,    -1,     0,     0,    -1,     2,     3,     8,     0,    -4,     4,     4,    -1,    -3,     4,     1,    -2,     1,    -1,    -1,    -5,    -4,    -2,    -1,     1,     1,    -2,    -4,    -7,    -6,    -4,     1,     5,     4,     5,     5,     4,     4,    -1,     2,     7,     1,     5,     3,     4,     2,     1,     0,    -6,    -9,    -5,     0,    -1,    -2,    -7,    -3,    -8,    -1,    -9,     0,     2,     2,     0,    -3,    -6,    -6,     6,     5,     3,     2,    -1,     3,     2,    -2,     3,     1,    -2,   -13,    -8,     0,    -1,    -2,    -1,    -6,   -17,    -8,    -2,    -1,     1,    -8,     1,    -3,    -4,    -2,    -1,     3,     0,    -5,    -2,     2,    -1,     3,     0,     3,    -4,    -7,    -3,    -2,     0,     0,     0,    -9,   -14,   -12,     4,     0,    -5,    -6,    -3,    -4,    -4,    -2,     2,    -2,    -2,    -2,     1,     5,     1,    -2,    -5,    -1,    -3,    -1,    -2,    -1,     1,     0,    -2,    -2,   -10,     2,     0,    -4,    -7,    -5,    -6,    -3,    -3,     1,    -1,    -3,     0,    -3,     0,     7,    -4,    -6,    -2,     2,    -6,     3,    -5,     1,     0,     1,     0,     0,     6,     5,    -6,    -7,    -6,     0,    -6,     2,    -1,     4,     2,     2,    -1,    -5,    -3,    -2,    -6,    -8,    -3,     3,    -2,    -5,    -5,    -1,    -1,     1,     1,    -5,     7,     1,    -4,    -9,    -6,    -5,    -6,    -4,   -11,    -9,   -10,   -10,    -7,   -10,    -8,    -4,   -11,   -16,   -17,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     0,    -1,    -2,    -2,    -4,    -5,    -5,    -9,    -7,    -5,    -6,   -10,    -1,    -5,    -7,    -4,    -6,    -7,    -6,    -7,     0,    -1,     0,     0,     1),
		    15 => (    0,    -1,     0,     1,    -1,     0,     0,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     0,    -1,     0,     1,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     1,     1,    -1,     1,     1,     0,    -1,    -1,    -3,    -3,    -3,    -2,    -3,    -5,    -3,    -2,    -2,    -1,     1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,     1,    -2,    -4,    -3,    -7,    -3,    -1,    -3,    -5,    -6,    -9,    -4,    -2,     1,     0,    -2,    -4,    -1,     1,    -2,    -1,    -1,    -1,     0,     0,    -2,     2,     1,    -3,     0,    -5,    -5,    -5,    -5,    -3,    -2,    -6,    -6,    -9,   -10,    -6,    -2,    -1,    -1,     2,     2,    -1,    -3,    -3,     1,    -1,    -1,     0,    -1,     2,    -1,    -1,    -1,     2,    -2,     1,    -5,    -4,    -7,    -7,    -1,     2,    -5,    -2,    -3,    -2,    -5,    -1,    -3,     2,     3,    -3,    -5,    -6,     0,    -1,    -2,     0,    -1,     1,     3,     3,    -5,    -5,     1,    -1,    -4,    -6,     1,     2,    -2,    -4,    -4,    -3,     1,    -1,    -6,    -8,    -6,    -1,    -3,    -4,     1,    -1,    -1,    -3,    -2,     3,     2,    -1,    -4,    -4,    -3,     1,    -2,    -1,     4,    -3,    -5,    -7,    -6,    -1,    -1,    -3,    -1,    -1,    -3,     0,     0,     4,     1,    -2,    -1,    -5,    -1,     1,     1,    -3,    -4,    -7,     1,     1,    -2,    -4,     2,    -4,    -6,    -6,   -12,   -12,   -10,    -4,    -1,    -2,     2,     2,     2,     3,     0,    -6,    -5,    -6,    -4,     5,     0,    -2,    -8,    -2,     3,    -4,    -1,     0,    -5,   -10,    -5,    -4,   -10,    -9,    -5,    -4,    -4,    -1,     1,    -4,    -9,     0,     0,    -1,    -2,    -5,    -3,     4,    -4,    -7,    -3,    -1,     2,     0,     0,    -8,    -2,    -7,     2,     2,     3,    -3,    -4,     0,    -2,     1,     6,     2,    -2,    -2,    -1,    -2,     0,    -1,    -4,    -2,     0,    -6,    -1,    -1,     3,     0,    -2,     4,    -1,     2,     6,     6,     6,     7,     5,     3,     4,    11,     7,     9,     2,    -2,     1,    -1,    -1,    -2,    -2,    -3,     3,    -3,     0,     1,     2,     5,     1,    -2,    -2,    -1,     5,     0,     4,     4,     8,     9,    10,    11,     3,     5,     0,     0,    -1,     0,    -1,    -4,    -7,    -2,    -1,    -2,    -1,     5,     5,     1,     2,     0,     3,     0,    -2,    -1,     0,     2,     9,     5,     8,     5,     1,     5,    10,    -1,    -1,    -1,    -1,    -2,    -8,    -2,    -4,    -4,     2,     1,     4,     1,     1,    -1,    -3,    -9,    -2,    -1,   -12,    -8,    -5,    -7,    -1,    -2,    -1,     0,     9,    -3,     0,    -1,    -3,    -6,     4,     3,    -1,    -1,     5,     2,     3,     6,     3,     3,    -8,    -9,    -7,    -6,    -4,    -9,    -3,    -5,    -2,    -4,    -5,    -6,    -3,     0,     1,     1,    -2,    -3,     9,    -1,     2,    -1,    -2,     4,    -1,     1,     6,     0,    -6,    -5,    -8,    -8,    -2,    -6,    -4,    -3,    -3,    -6,    -1,    -9,    -2,    -3,    -2,    -2,    -2,     0,    -7,    -5,    -8,    -3,    -6,    -4,    -2,    -2,     0,     0,    -2,    -1,    -1,     0,    -1,    -5,    -6,    -2,    -6,    -2,    -3,    -8,    -4,    -3,    -1,    -1,    -2,    -3,    -4,    -6,    -7,   -11,    -9,    -2,    -8,     0,    -2,    -6,     1,     0,    -3,    -1,     0,    -2,     0,    -2,    -8,     4,    -5,    -9,    -5,    -8,    -1,     0,    -2,     1,     0,    -1,     0,    -2,    -6,    -3,    -3,     2,     2,    -4,    -6,    -7,     4,     2,     1,    -4,    -1,    -4,    -4,     2,    -3,    -2,    -5,    -4,     0,    -1,     3,    -5,    -1,    -5,     4,     3,    -4,    -2,    -1,     1,    -2,     0,     2,     1,     5,     1,     3,     0,    -2,    -5,     2,     5,    -2,    -6,    -6,    -5,    -1,    -3,     2,    -5,    -4,    -3,     3,     5,    -1,     2,     4,    -3,    -1,     1,    -4,     0,     4,     3,    -2,    -1,    -4,     2,     4,     1,    -2,     0,    -7,     1,     0,    -1,    -1,     0,    -4,     2,     5,     6,     1,     0,     1,    -3,    -5,     2,    -4,     2,     2,    -1,     4,     1,     3,     3,     0,     0,    -6,    -1,    -6,    -1,     0,     1,    -1,     3,    -1,    -2,     2,    -2,     3,     0,     3,     2,     6,     2,     3,     3,     0,     2,     0,     2,     3,     1,    -2,    -1,    -5,     0,    -2,    -1,     0,     1,     3,    -2,    -4,    -6,    -2,    -1,     4,     2,     2,     1,     3,     7,     4,    -2,    -1,     1,    -4,     2,     3,    -2,    -4,     1,     0,     0,    -1,     0,    -1,    -1,    -3,    -1,    -1,    -6,    -5,    -5,     4,     5,     3,     2,     1,    -2,     4,     1,     1,     4,    -2,     2,     1,    -6,    -3,     1,    -1,    -6,    -2,     1,     0,    -1,    -1,     1,    -3,    -8,    -4,    -9,    -6,    -8,    -6,    -4,    -5,    -7,    -5,    -3,    -6,    -8,    -5,    -4,    -2,    -2,    -2,    -1,     0,    -1,     1,    -1,     0,     1,    -1,    -1,    -1,    -5,    -7,    -6,     0,    -3,     2,    -2,    -5,    -9,    -8,    -9,    -7,    -4,    -6,    -1,    -2,     1,     0,    -3,     0,     1,     1,    -1,     1,    -1,    -1,    -1,    -2,     0,    -1,    -2,     0,     0,     0,    -1,    -1,    -2,    -7,    -3,    -3,    -1,    -1,    -3,    -4,    -5,    -5,    -1,    -1,    -1,     0,    -1),
		    16 => (    1,    -1,     1,     0,     1,    -1,    -1,     0,     1,     0,     0,    -1,     2,     0,    -1,     0,     0,    -1,     1,     1,     0,     0,     0,    -1,     0,     0,     1,    -1,     0,     0,     0,    -1,     1,    -1,     0,     4,     1,     1,     1,     1,     4,     2,    -3,     0,     2,     2,     1,     0,     6,     1,     2,     1,     1,     0,     0,     1,     0,     0,     2,     0,     1,     1,     2,     3,     3,    -2,    -2,     0,    -4,    -3,     2,     2,     7,     9,     1,    -4,    -6,     3,     5,     4,     2,    -2,     0,     0,    -1,     0,    -1,     0,     2,     4,    -1,    -1,     0,    -2,    -2,    -1,    -5,    -2,     4,     4,     8,     3,    -1,     2,     7,     3,    -3,    -1,     0,     0,     0,    -1,     1,     0,    -4,    -3,     6,     6,    -1,    -1,    -3,    -2,    -2,    -5,    -6,    -2,    -5,     0,    -1,     0,    -3,    -2,     0,    -5,     1,    -4,    -4,    -2,     3,     3,     1,     0,    -2,     0,     7,     6,     1,    -1,    -1,    -1,    -6,   -10,    -3,    -6,    -2,    -2,     3,     3,    -2,    -1,    -8,    -7,    -1,    -5,    -1,     0,     3,     1,     1,     0,     1,    -3,     4,     4,    -1,     0,    -2,    -3,    -9,   -10,    -6,    -1,     1,     5,     0,    -6,     3,     3,    -1,    -8,    -1,    -2,     0,    -1,    -1,     1,     1,    -1,     0,    -6,     3,     4,     0,    -3,    -3,    -4,    -7,   -10,    -5,     0,     1,    -7,    -4,    -8,    -4,     1,     1,     3,     3,     0,    -1,     2,     1,    -2,     0,     0,    -1,    -6,     3,     4,     1,     0,    -4,    -5,    -7,   -10,    -2,     1,     1,    -5,    -3,    -5,    -7,    -5,    -2,     5,     2,    -2,    -1,    -1,    -4,    -6,     1,     0,     0,    -3,     6,     5,     1,     2,    -2,    -5,    -5,    -1,     2,     3,    -1,     1,    -5,    -3,    -6,    -5,    -5,    -5,    -4,     0,    -1,     0,     0,    -2,     1,    -1,    -2,    -4,     6,     6,    -1,    -2,    -3,    -2,    -1,    -4,     3,     0,     0,    -8,    -5,    -6,   -10,    -7,    -6,    -7,    -4,     1,     1,     0,    -2,    -1,    -1,     1,     0,    -4,     7,     7,    -1,    -2,    -3,    -6,    -4,     1,     0,    -3,    -4,    -6,    -4,    -7,    -9,    -8,    -5,    -8,    -6,     1,     2,     1,    -1,    -3,     0,     0,    -1,    -3,     4,     6,    -2,    -4,    -4,    -2,    -1,     5,     2,    -3,    -2,     0,    -6,    -9,    -6,    -3,    -3,    -7,    -6,     4,     3,     0,    -4,    -3,     1,     0,     1,    -3,     4,     4,     0,    -3,    -2,    -3,     0,     3,    -1,    -1,     1,     2,     5,     2,    -3,    -3,    -2,    -5,    -5,     2,    -4,    -5,    -4,     0,     1,     1,    -1,    -1,     0,     3,     2,     1,    -1,    -7,     0,     0,     0,    -2,    -4,    -1,     4,    -3,    -6,     0,     3,    -4,    -4,    -1,    -2,    -2,    -2,    -1,     1,     0,    -1,    -4,    -1,     1,     1,     0,    -3,    -5,     0,     0,     0,    -9,    -1,    -1,     2,     6,     0,     6,     5,    -3,    -1,    -2,    -3,    -3,    -2,    -5,    -1,     1,    -1,    -4,    -2,     2,     0,     3,     2,    -5,    -1,     6,     5,    -5,    -1,    -6,    -1,     2,    -3,     3,     0,    -5,    -2,    -4,    -2,    -1,    -2,    -2,     0,     1,     1,    -4,    -3,    -1,     1,     2,     2,    -5,     3,     8,     2,    -9,    -8,    -3,     1,    -4,    -1,     2,     0,    -4,    -4,    -2,    -3,    -6,    -1,    -4,     1,     0,     0,     1,    -3,     0,     0,     0,    -6,    -4,     0,     1,     3,     0,    -7,    -5,     0,     2,     2,     2,    -7,    -4,    -6,    -5,    -6,    -7,    -1,    -3,     0,    -1,     0,     0,    -2,    -3,    -4,    -4,    -4,    -6,    -1,     7,     4,     4,     0,    -2,    -4,     3,     1,     1,    -4,    -3,    -5,    -4,    -5,    -3,    -4,    -1,     1,    -1,    -1,    -1,     0,    -2,    -3,    -5,    -5,    -8,    -7,    -1,     2,     4,    -1,     0,    -1,     5,    -1,     3,     2,    -3,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,     1,     0,     1,    -1,    -2,    -3,    -5,    -7,    -7,    -7,     0,     3,     0,    -1,    -3,    -1,     0,    -1,    -6,    -3,    -2,    -1,    -3,    -3,     0,     1,     1,     0,     0,    -2,     0,    -1,     1,     0,    -4,    -8,     1,    -3,     0,     1,     4,     4,    -3,    -6,    -6,     2,    -1,    -2,     1,    -2,    -5,    -1,     1,     1,     1,    -1,    -1,    -2,     1,    -1,     0,    -1,    -1,    -5,    -6,    -4,     1,    -2,     1,    -2,    -2,    -3,    -1,     1,    -2,    -2,     1,    -1,     0,    -1,     1,     0,     1,     1,     0,    -1,    -2,    -2,    -1,     0,    -3,    -2,    -3,     1,     2,     2,     0,     5,    10,     4,    -6,    -9,    -3,     0,     0,    -1,    -1,    -2,     0,     0,     0,    -1,     0,    -1,     1,    -1,    -1,    -1,     0,    -2,    -1,     0,     3,     2,    -1,    -1,    -2,    -1,    -1,    -2,    -3,     0,    -1,    -2,     0,     1,     1,     0,     0,     1,     1,     0,    -1,     0,     1,     0,     1,     0,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     0,    -1,     0,    -2,     0,     0,     1,     1,    -1,     1,    -1,    -1,     1,     1,     0,     0,    -1,    -1,     1,    -1,     0,     1,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,    -1,     1,     0,     0,     0),
		    17 => (    0,     0,    -1,     1,     0,    -1,    -1,    -1,     1,     1,    -1,     1,     0,     1,     1,    -1,     0,    -1,     1,    -1,    -1,     1,    -1,     1,     0,     0,     0,     1,    -1,     0,     1,     0,     1,     1,     0,     0,    -1,     0,    -1,    -5,    -4,    -3,    -1,    -4,    -4,    -3,     0,     1,     1,     1,     0,    -1,     1,     0,     0,     0,     0,     1,     0,    -3,    -2,     0,    -1,     0,    -2,    -1,    -1,    -4,    -2,    -2,     0,    -3,    -3,     0,     0,     1,    -1,     0,    -1,     0,     1,     0,     1,     0,     1,     0,     1,    -4,    -1,    -2,    -2,    -3,    -5,    -3,    -3,    -2,    -2,    -3,    -2,    -3,    -1,    -1,    -2,    -1,    -1,    -2,    -6,    -2,     0,    -2,     1,    -1,     0,     0,    -1,     0,    -6,    -3,    -1,    -8,    -8,    -4,    -8,   -13,   -11,   -10,    -8,    -4,    -2,     0,     0,    -1,    -5,    -6,    -3,    -6,    -2,    -3,    -1,     0,     1,     1,     0,    -1,    -6,    -3,    -2,     2,     2,    -1,    -5,    -3,     1,     0,    -7,    -8,    -9,   -17,   -19,   -18,   -17,   -10,    -1,    -6,    -4,    -3,    -1,    -1,    -1,     1,     6,     6,    -1,    -1,     0,    -3,    -3,    -6,    -8,     3,     5,     2,    -3,   -10,    -8,     0,    -1,    -1,    -2,     6,     4,     1,    -4,    -5,    -8,    -2,    -1,    12,    11,     7,     1,    -1,     0,     5,    -1,     0,     1,    -3,     3,    -1,    -4,    -5,    -5,    -2,    -1,    -2,    -4,     1,    -1,     3,     3,    -1,    -6,    -3,    -7,    12,     4,     1,    -3,    -4,    -3,    -1,    -5,    -1,     5,     0,     2,    -4,    -4,    -2,    -4,     2,     3,     0,    -2,    -4,    -2,     5,     8,     2,    -5,    -4,     1,     7,    -5,    -1,     2,     0,     3,    -1,    -3,     1,     1,     2,     1,     0,     6,     0,    -4,     2,     4,     3,     1,     1,     1,     3,     9,    -1,    -8,     0,     1,     5,     4,     1,     2,     1,     5,     2,     2,     0,     0,     5,     5,     6,     0,    -5,    -4,     2,     0,     3,     5,     4,    -3,    -2,    -4,    -3,    -7,     2,     0,     1,     5,     6,     2,     7,     1,    -3,    -5,     5,     2,     9,    10,     0,    -8,    -5,    -3,    -1,     7,     4,     5,    -2,    -4,     0,    -2,    -6,    -3,     1,     1,     2,     3,     4,     1,     4,     1,     5,     3,     3,     5,     3,     6,   -15,   -17,    -3,     2,     2,     4,     0,     2,    -2,    -5,    -5,    -3,    -4,    -1,     3,     0,     2,     6,    -1,    -1,     6,     4,     5,     4,    -1,     1,     0,    -3,   -21,   -14,    -7,     3,     0,     4,    -3,     0,     2,    -4,    -8,     0,    -7,    -2,    -1,    -1,     4,    11,     4,    -3,     7,     2,    -2,    -1,     4,     6,     1,   -10,   -28,   -13,    -5,     3,    -1,     5,     3,    -1,    -1,    -1,    -1,     0,    -4,    -3,    -1,    -1,     0,     3,     4,   -10,     3,     4,     3,    -4,    -3,     7,    -4,   -24,   -17,    -9,    -4,     3,     3,     2,     5,     0,    -2,     1,    -4,    -6,    -5,    -1,    -2,    -2,    -2,     2,     2,    -5,    -4,     1,     7,    -1,    -1,     8,   -10,   -23,    -3,     0,    -1,    -2,     1,     4,     4,    -5,     0,     3,    -3,    -3,    -5,     0,    -5,    -1,     1,     3,    -2,     1,    -3,     1,    -1,    -4,    -8,   -12,   -16,   -13,    -1,     2,    -1,    -2,    -3,     4,    -3,     1,    -1,     4,   -12,   -15,    -3,     0,    -6,     3,    -1,     7,   -10,    -4,    -1,     2,     1,    -6,   -12,   -20,    -5,    -2,     3,     6,    -1,     2,     3,     3,    -3,     4,    -3,    -4,   -15,   -14,     2,     0,    -2,    -1,     4,     2,    -8,    -1,     2,     2,   -13,   -13,   -15,   -16,    -5,    -1,     0,     1,     0,    -2,    -3,     2,     0,    -2,    -6,    -9,   -11,    -7,     5,     0,    -1,     0,     4,     0,    -5,    -3,    -3,    -5,   -12,   -12,   -16,    -3,     6,     4,    -3,     0,    -4,    -3,     1,    -3,    -1,    -4,    -9,    -8,   -12,    -4,     0,     0,     0,    -1,     0,    -2,    -6,   -11,    -3,   -11,   -10,    -9,    -3,     8,     3,    -3,    -4,    -3,    -7,    -4,    -1,     3,     1,    -1,    -2,     0,    -2,    16,     1,    -1,     1,     0,     1,    -1,    -3,    -7,     1,     1,     0,     1,     3,     1,     2,    -3,     0,     1,     0,    -1,     1,     2,     3,     1,    -3,     0,    -2,    -1,     0,    -3,     0,     1,     1,    -1,    -7,    -4,     4,     6,     3,     4,     0,     2,    -8,     0,     3,     0,     0,    -3,    -2,     3,    -5,    -2,    -1,   -11,    -7,    -1,    -2,    -1,    -1,    -1,     0,     2,     2,     0,     5,    -2,    -6,     4,    -1,     1,     2,     1,     0,     3,    -2,    -3,    -3,    -8,    -5,    -2,     2,    -9,    -9,    -2,    -7,     1,     0,     1,     0,    -1,     0,    -9,   -11,    -4,    -3,     0,    -1,     2,     2,     2,     0,     4,     0,     2,     3,    -5,    -2,    -2,     2,     0,    -6,     2,    -1,    -1,     1,     0,     0,     1,    -1,   -10,    -9,    -7,    -8,    -3,    -5,    -5,    -6,     1,     5,     5,     1,     3,    -1,     0,     2,    -2,    -2,    -1,     0,    -2,     1,     0,     0,     1,     1,     1,    -1,     3,     3,     1,     3,     5,     2,     3,     1,    -2,    -1,     1,    -3,    -3,     6,     5,    -5,     3,     9,     2,     5,    -1,     1,     0,     0),
		    18 => (    1,    -1,     0,     0,     1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     1,    -1,    -1,     0,     0,    -1,     1,     1,    -1,     0,     0,    -1,     1,    -1,    -1,     1,    -1,     0,     0,    -1,    -2,    -3,    -5,    -9,    -4,    -2,    -2,    -2,    -3,    -2,     0,     1,     1,    -1,     0,     1,     0,    -2,     0,     0,    -1,    -3,    -2,    -3,    -7,    -9,    -5,    -1,     0,    -2,    -6,    -4,    -1,     2,    -3,   -10,    -8,    -9,    -3,    -2,    -2,     1,     1,    -1,     0,    -4,    -4,     0,    -3,    -4,   -10,     2,     1,    -1,    -4,    -5,    -7,   -11,     0,     2,     1,     4,     2,     9,     8,     3,     3,    -3,    -1,    -3,     0,     0,     1,     0,    -6,    -6,    -9,     0,     0,    -4,    -6,     1,    -3,    -8,    -7,     3,     0,     1,    -1,    -1,     3,     7,     7,     4,     3,     0,     9,     4,    -1,    -1,     0,    -5,    -6,   -10,    -3,    -1,     1,     3,    -1,     0,     0,    -3,    -3,    -3,     1,     0,    -4,    -5,    -2,     6,     3,     2,     8,     8,     4,    -3,     0,     0,     0,    -4,    -6,    -2,    -5,     1,     2,     3,    -1,    -2,    -3,     2,     0,     1,     0,    -6,    -6,    -2,     3,     0,    -3,    -6,     2,    -1,    10,     1,    -5,    -1,    -7,    -4,    -1,     0,    -6,     2,     7,     0,    -3,    -2,    -1,     1,     0,     1,     2,    -6,    -1,     4,     2,    -3,     0,     3,     3,     2,    -1,    -1,    -6,    -2,    -2,    -4,     2,     7,    -2,     5,     5,    -5,     3,    -1,     1,     1,     5,    -2,    -8,    -3,    -3,    -3,    -7,     1,     6,     4,    -1,     1,     4,     3,     2,     0,     1,    -1,     4,     2,    -6,    -3,    -2,    -3,    -2,     2,     5,    -2,    -2,    -6,    -8,     0,    -1,    -5,     2,     2,     2,     1,     5,     1,     1,    -6,   -14,     1,    -1,    -2,    -4,     0,    -6,    -4,    -7,     1,     4,     5,     1,    -1,    -5,    -5,    -5,     1,     5,    -2,    -2,    -2,    -2,     0,     3,     0,    -9,    -5,   -11,     0,    -1,    -4,    -5,    -5,    -3,    -2,     1,    -3,     3,     0,     6,     5,    -1,    -2,    -4,     0,    -3,    -2,    -8,    -4,   -10,    -5,     5,     9,     1,     8,    -6,     0,     1,    -6,     7,    -3,     6,     1,     2,    -6,    -3,     0,    -4,     3,     5,    -1,    -3,    -4,     0,     1,     4,    -6,    -1,     5,    11,    10,     3,     2,   -11,     0,     0,    -5,     5,    -2,    -3,   -10,    -4,    -5,    -5,    -1,    -1,     1,     3,     1,    -1,    -7,     2,    -1,     3,     4,     8,    12,    11,     5,    -3,    -3,     2,    -2,     0,     0,    -9,     0,    -9,    -4,    -4,    -7,    -9,     0,    -4,     0,     5,     2,     1,    -6,     5,    -6,     3,     0,     6,     1,     9,     5,    -3,    -7,     0,     0,     1,    -1,     3,    -1,     2,     1,    -3,     0,    -8,    -2,     1,     3,     2,     0,    -2,     4,   -11,    -4,     2,    -4,    -8,    -2,     6,     7,     0,    -9,    -6,     0,    -1,    -3,     4,    -6,     6,    -2,     1,    -5,    -6,    -3,    -1,     5,     1,    -1,     1,    -5,    -2,    -2,    -7,    -9,    -7,    -5,     3,     1,     2,    -7,    -5,     0,    -1,    -3,     3,    -9,    -1,    -1,     4,    -3,    -5,     1,     4,     5,    -3,     5,     5,    -2,    -2,    -9,    -7,    -4,    -7,    -4,     0,    -1,     1,    -1,    -3,    -2,    -1,    -1,    -4,    -6,    -3,    -2,    -4,    -5,     5,     4,     7,    -3,   -11,    -2,     5,     0,    -1,    -2,     3,    -2,   -11,    -3,     0,    -7,     1,    -1,    -3,     0,    -1,    -3,    -2,    -7,    -3,    -3,    -6,     5,     2,     6,     6,    -5,   -10,    -5,     2,     1,     4,    -5,    -1,    -3,    -7,     0,    -4,    -5,     0,    -4,    -2,     0,     1,    -1,    -3,   -11,    -1,    -5,     4,     3,     3,     5,     6,     1,    -3,    -1,     1,     0,    -3,     0,     1,    -3,    -3,    -4,    -5,     0,     1,    -5,     0,    -1,    -4,    -3,     0,   -10,   -11,     1,     2,     2,     2,     0,    -1,     2,    -5,    -4,     2,    -5,    -3,     2,    -3,   -11,    -6,    -1,    -4,    -2,     3,    -6,     0,    -1,    -1,    -2,    -4,    -7,   -14,    -7,     2,    -2,     1,     0,     3,    -1,     3,    -4,    -1,   -10,     0,     1,    -9,   -15,    -7,    -4,    -4,     1,     3,    -9,     0,     0,     0,    -4,    -6,    -8,   -10,    -3,     0,     6,    -4,    -6,     1,     3,     1,     2,    -5,    -2,     6,    -7,   -14,   -13,    -6,    -6,    -2,     3,     3,    -8,     1,    -1,     0,    -1,    -1,    -9,   -12,    -6,     0,     3,     0,    -1,     1,     5,     5,     3,    -1,     3,    -5,    -7,    -8,    -4,    -3,    -4,    -1,    -3,    -7,    -7,     0,     0,     0,    -4,    -3,    -4,    -6,    -2,    -1,    -5,    -5,     5,    -6,    -7,    -3,    -1,     4,    -2,     0,     2,     4,     4,    -2,    -4,    -2,    -6,    -3,    -3,     0,    -1,     0,     1,    -1,    -2,    -4,    -7,    -1,     1,    -4,    -9,    -6,    -5,    -7,   -10,    -9,    -4,    -2,     0,    -2,    -3,    -4,    -3,    -1,     0,     1,     1,     0,     0,     0,    -1,     1,    -2,    -1,     0,    -3,    -4,    -2,    -2,    -2,    -1,    -2,    -2,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     1,     0),
		    19 => (    0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,    -1,    -1,    -1,     1,     0,     1,     1,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,     1,     0,     1,    -1,     0,     1,     0,     1,    -1,    -1,    -1,     0,     1,    -1,    -2,     0,    -3,    -3,    -4,    -2,    -1,     0,    -2,     0,     0,     1,     1,    -1,     0,    -1,     1,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     1,     0,    -3,    -1,     0,    -1,    -3,    -1,    -2,     1,    -1,    -1,    -1,    -1,    -1,     1,     0,     1,    -1,     0,    -1,    -5,     0,    -1,    -4,     0,    -1,     0,    -1,     0,    -3,    -8,    -4,     2,     8,     3,    -5,    -2,    -3,     0,    -1,    -2,    -1,     1,    -1,     0,    -1,    -2,     0,    -3,    -3,     0,    -1,     0,     1,    -1,    -4,    -6,    -7,   -12,   -13,   -13,    -8,   -10,   -11,    -6,    -6,    -7,    -4,    -6,    -3,    -1,     1,     0,    -2,    -1,    -1,    -1,    -1,     0,    -5,    -1,    -2,    -5,   -11,   -12,   -16,   -16,   -13,   -11,    -3,    -3,     1,    -1,    -5,    -9,    -7,    -5,    -6,     1,    -1,    -2,    -4,    -4,     3,     0,    -3,    -4,    -4,    -9,    -7,   -15,   -17,    -9,    -1,    -2,    -1,     5,     4,    -4,    -1,    -2,    -5,    -8,    -5,    -4,    -5,    -6,     0,    -3,    -5,    -2,    -3,    -2,    -4,    -5,    -2,   -12,   -17,   -10,    -3,     3,     3,     7,     6,    -3,     3,    -1,     5,    -4,    -2,     2,    -7,    -5,    -4,    -3,    -5,    -4,    -4,     1,    -1,     0,     8,    -3,    -1,    -5,    -7,    -3,     2,     3,    -3,    -5,     0,     1,     2,     4,    -7,     0,     6,     4,    -8,    -8,    -4,    -2,     0,    -4,     4,     4,     5,     1,    -2,    -4,    -9,    -3,     1,     3,     4,     0,    -7,     0,    -7,   -12,    -4,     0,    -4,    -4,    10,    -4,    -4,    -9,    -2,    -4,     0,    -5,    -9,     4,     5,     1,    -4,    -8,    -3,     2,     3,     5,     2,     1,     1,    -1,    -6,    -7,     0,     0,    -2,     1,     0,    -4,    -2,    -7,    -5,    -3,     0,    -2,    -4,     1,    -1,    -1,    -2,    -1,    -3,    -3,    -1,     4,     1,     3,     0,    -1,     2,    -3,     4,     0,    -2,     1,     1,    -3,    -2,    -3,    -6,    -3,     0,     0,     2,     1,     2,    -4,    -5,     0,    -1,    -3,     2,     1,     1,     0,    11,     7,     5,    -1,     1,    -7,   -12,    -2,    -7,    -2,    -5,    -8,    -7,    -7,     1,    -2,    -2,    -2,    -1,    -3,     1,    -5,     1,    -2,     5,     8,     4,     3,     3,     4,    -2,     0,    -2,   -16,   -15,    -5,    -7,    -2,     1,    -4,    -3,     0,    -2,    -1,    -4,    -2,    -2,    -1,    -2,     1,    -4,    -4,     1,     1,     0,     1,     5,     2,    -1,    -1,     0,   -13,    -9,    -6,    -4,    -3,     1,     0,     0,    -1,    -1,    -1,    -5,    -1,    -2,    -5,    -1,     0,     1,    -3,     3,     1,     2,     2,     4,     2,     6,     2,     4,   -17,   -12,    -4,    -5,     2,     2,    -2,     7,     1,     0,    -1,    -4,     0,    -1,   -11,    -8,    -3,     0,     0,    10,     4,     4,    -4,    -3,    -1,     1,     1,   -15,   -20,    -6,     5,     2,     0,     8,    -5,    -2,     0,     1,    -2,    -3,    -1,    -2,    -9,    -9,    -5,    -6,    -3,     4,     2,    -6,     0,     5,     0,    -3,    -4,    -9,    -9,     3,     7,    -6,    -4,     6,    -2,    -5,     0,     4,    -1,    -3,    -2,    -4,    -4,    -3,   -12,   -13,    -5,    -1,    -3,    -7,     2,     3,     2,    -6,    -5,    -8,    -8,     6,     6,     1,    -2,     0,     0,    -6,    -4,     0,    -3,    -4,    -2,    -5,    -7,    -6,    -9,   -16,   -13,   -10,    -9,    -1,     1,    -2,    -1,    -7,    -3,    -9,    -2,     3,     8,     1,    -3,    -2,     0,    -2,    -3,     0,     0,    -3,    -3,    -5,    -1,    -4,   -11,    -8,    -4,    -6,     0,     0,    -3,     0,    -7,    -5,    -5,    -7,     5,     1,    -2,    -1,    -2,     5,     3,    -1,    -1,    -1,     0,    -4,    -4,    -5,    -2,     2,    -2,     1,    -1,    -1,    -3,     1,    -1,    -2,     0,    -2,    -7,    -4,     5,     5,    -1,     0,     6,    -8,     5,    -4,    -1,     0,     1,    -3,    -6,     0,     2,    -4,     1,     2,     0,    -3,     1,    -5,    -7,    -3,    -3,    -3,   -10,    -4,     4,     8,     0,    -2,     5,     8,     0,     1,    -1,    -1,    -1,    -2,    -2,    -6,     1,    -2,     5,     1,     2,     1,    -5,    -2,    -4,    -5,    -7,    -4,    -6,    -5,     3,     9,     1,     0,    -2,     5,    -4,     1,     0,     0,     0,    -1,    -4,    -3,     2,     0,     4,    -1,     1,    -1,    -5,     0,    -3,    -4,    -5,    -3,    -2,    -8,    -5,     3,    -1,     0,     1,    -5,    -3,    -4,    -1,    -1,     0,     3,    -1,     6,    -2,     0,     5,     0,    -6,    -4,     4,    -2,     2,    -5,    -3,    11,     3,    -5,    -3,     2,     2,    -1,     2,    -6,    -5,    -4,     0,    -1,     0,     1,     7,     8,     1,    -1,     5,    -1,     3,    -3,     4,     8,     3,     7,     2,    13,    12,     0,    -8,     1,     3,    -2,    -2,     0,    -1,     0,    -1,    -1,     1,     0,    -1,     0,    -1,     1,     1,     0,     0,     4,     8,     7,     7,     9,     5,     3,    -2,    -2,    -2,    -3,    -2,     0,    -1,     1,     0,     0,     1),
		    20 => (    0,    -1,    -1,     0,    -1,    -1,     1,     1,     0,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,     1,     1,     1,    -1,     0,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,     0,     1,     1,     0,    -2,    -4,    -5,    -5,     1,     1,     0,    -1,     5,     3,     3,    -1,     0,     0,     0,    -1,    -1,    -1,     1,    -1,     0,     0,     1,     0,     2,     3,    -1,    -2,     0,    -3,    -5,    -3,    -1,     1,    -2,    -5,    -4,     0,     0,     1,    -1,     0,    -1,    -5,    -4,    -2,    -2,     0,     1,     0,     1,    -1,     2,     0,    -5,    -3,    -1,    -5,   -10,    -3,    -4,    -3,    -8,    -6,    -2,    -2,     1,    -2,    -2,    -7,    -6,    -5,    -8,    -3,    -4,    -5,     0,     1,     0,    -2,    -4,    -3,    -9,    -3,    -2,    -3,    -2,     0,     0,    -5,    -4,    -3,    -2,     3,     4,     3,     3,    -2,    -5,    -4,    -5,     1,   -10,    -4,     1,     0,     0,    -3,    -1,     2,    -4,    -2,    -5,    -5,     0,     1,     1,    -2,    -3,     1,     2,     6,     5,     6,     3,    -2,    -1,    -7,    -6,    -1,    -9,    -4,     0,     0,    -1,    -3,     0,    -1,     0,    -1,    -2,    -5,    -4,    -1,    -1,    -3,     1,    -1,     3,     4,     4,     5,     3,     5,     2,     0,    -1,    -3,    -5,    -1,     3,    -1,    -4,    -6,    -4,    -3,    -2,     0,     1,    -6,    -3,    -2,    -1,    -1,     0,     2,     0,     1,     3,     1,     2,     3,    -2,     2,     0,     0,     2,    -5,     1,     2,    -7,     1,    -3,    -4,    -2,    -5,    -3,    -5,    -4,    -3,     0,     0,    -1,    -2,    -4,    -2,     0,     3,    -1,     1,     3,     1,     1,    -1,    -3,    -5,    -1,    -1,    -2,     1,    -1,    -4,    -4,    -7,    -2,    -5,    -4,    -5,     0,    -2,    -2,    -6,    -5,    -3,    -4,    -6,    -6,    -4,    -4,    -3,    -3,    -1,    -7,    -7,     0,    -1,     1,     4,     0,    -5,    -7,    -3,     0,    -5,    -5,    -6,    -7,    -8,    -8,    -4,    -5,    -3,    -2,    -5,    -5,    -9,   -10,    -3,    -2,    -4,    -3,    -5,    -1,    -1,     6,    -6,     1,    -4,    -2,     2,    -3,    -8,    -6,    -6,    -6,    -6,    -4,    -4,    -2,    -4,    -3,    -2,    -1,    -4,    -5,    -1,    -2,    -2,    -3,    -2,    -1,     0,     1,    -8,     2,    -3,     0,    -1,    -3,    -3,    -1,    -2,     0,     1,     1,     1,    -1,     0,    -1,     2,     1,     1,    -1,     1,    -1,    -2,    -4,    -3,    -2,     0,     2,     0,     1,     0,    -1,     1,    -2,    -4,     0,    -3,    -2,    -1,     1,     0,    -4,    -2,     0,     4,     0,    -4,     0,     1,     2,    -1,    -1,    -5,    -4,     0,     0,    -2,    -5,     1,     0,    -1,     1,     1,    -1,    -7,    -4,    -3,    -2,    -7,    -6,    -4,    -1,    -1,    -5,    -2,    -1,     0,    -4,    -2,     3,    -6,    -1,     1,     1,    -1,    -7,     2,     2,    -4,     1,     1,    -5,    -7,    -8,    -5,   -11,   -12,    -5,    -4,     0,    -1,    -1,     2,     0,    -3,    -5,    -1,     1,    -7,    -2,     1,     0,    -4,    -1,     5,     0,    -4,    -5,    -1,    -7,    -9,    -6,    -9,   -11,    -7,     0,     0,     3,     1,     0,     3,    -2,    -3,    -1,     2,     2,    -9,     1,     0,    -1,    -4,    -1,     1,     0,     1,     1,    -1,     0,    -6,    -5,    -3,    -3,    -2,     3,     1,     4,    -1,     2,    -1,    -3,    -2,     3,     2,     1,    -9,     2,    -2,    -1,    -3,    -1,     2,    -2,     1,     1,     1,     1,    -1,    -4,    -6,    -4,     0,     5,     3,     3,     0,    -2,    -3,    -2,     1,     2,     1,     0,    -5,    -4,     0,     1,     0,     0,     1,     1,    -1,     4,     2,     2,    -1,    -1,     0,    -5,     0,     3,     0,    -5,    -8,    -5,    -1,     5,     2,     1,     4,    -8,    -3,    -3,    -1,     2,     2,     1,     0,     1,    -2,    -1,    -1,    -2,     0,    -2,    -2,    -4,    -1,     0,    -3,    -6,    -3,    -1,     0,    -1,    -1,     3,     2,    -2,    -1,    -1,     1,     1,    -2,     0,    -1,    -1,    -2,    -1,     0,     0,    -2,    -6,    -4,    -7,    -3,     1,    -3,    -3,     0,     1,     1,    -4,    -1,     3,     2,     0,     2,     1,     0,    -1,    -5,     0,     2,     0,     0,    -1,    -1,    -1,    -5,    -2,    -3,    -2,     0,    -5,    -1,    -4,     0,     0,    -3,     0,     2,     1,     1,    -1,     0,     0,    -1,     0,    -4,    -4,    -3,    -2,    -1,    -1,    -6,    -4,    -1,     1,     1,     0,    -3,    -2,    -1,     1,     2,     1,    -2,     2,     3,     1,    -7,    -5,    -3,     0,    -1,     1,     0,    -3,    -4,     2,    -5,    -2,    -2,    -4,    -9,    -7,    -5,    -5,    -6,    -4,    -3,     2,    -1,     0,    -2,    -2,    -2,    -3,    -2,    -1,    -1,     1,    -1,     0,     0,    -4,    -6,    -4,    -4,    -3,    -3,    -3,    -4,    -7,    -7,    -9,    -8,    -6,    -6,    -2,    -2,    -8,    -5,    -5,    -5,    -3,     0,     0,     1,     0,     0,    -1,    -1,     1,    -5,    -6,    -8,    -4,    -2,    -4,    -5,    -1,    -2,    -4,    -4,    -6,    -5,    -8,    -8,    -9,    -6,    -6,    -5,    -2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -4,    -4,    -3,    -1,     0,    -1,    -3,     1,    -1,    -2,    -3,    -2,    -3,    -1,    -2,    -3,    -2,    -1,     0,     1,    -1),
		    21 => (    1,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     1,     1,     1,     0,     1,     0,    -1,     1,     0,     1,     0,     0,     0,     1,     0,    -1,    -1,     1,     1,     1,     1,    -1,     0,     1,     0,     1,    -1,    -1,     1,     0,    -3,     5,     6,    -1,    -5,    -2,    -3,     0,    -1,    -1,     1,     1,     1,    -1,    -1,     1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -6,    -6,    -4,   -10,    -3,    -6,    -5,    -1,    -5,    -3,    -1,    -2,    -7,    -9,    -5,    -4,    -2,     0,     0,     0,    -1,     9,     6,    -1,    -5,    -1,     5,     5,     6,     2,    -8,    -5,     7,    -1,    -7,    -6,    -2,    -2,    -4,    -1,   -12,    -8,    -5,    -5,    -2,     1,     1,    -1,    -1,     8,     8,     1,    -3,     0,     7,     7,     7,     4,    -2,    -1,     3,    -1,     0,    -6,    -6,    -2,     1,    -3,    -8,    -4,    -4,    -4,    -9,   -10,    -7,    -1,     0,     7,     1,     2,     4,     4,     7,     2,     6,     9,    10,     5,     5,     1,    -3,    -3,    -2,    -3,     1,    -3,    -6,    -5,     3,     1,   -15,    -7,    -6,     0,     0,    -3,     0,     3,     1,     5,     9,     2,     3,    11,     5,     2,     4,     1,     0,    -2,     0,     0,     0,    -1,    -5,    -3,     4,     0,    -7,    -8,    -4,     0,    -6,    -9,    -7,   -11,     4,     7,    10,    -3,    -4,     5,     2,     5,    -2,     5,     0,     2,     2,    -5,    -4,     3,    -3,     4,     3,    -2,    -5,   -14,    -9,    -2,    -6,    -8,   -11,   -11,    -1,     7,     8,    -4,    -9,     4,    -4,     2,     6,     4,     3,     1,     4,     6,     2,    -2,    -1,     3,    -1,    -7,    -6,   -14,    -6,     1,    -2,    -8,   -11,    -8,    -4,     0,     5,    -2,    -3,    -5,    -7,    -3,     7,     1,     2,    -1,     5,     7,    -2,     1,     2,     1,    -4,    -6,    -6,    -6,    -8,     0,    -4,    -7,   -10,    -8,    -5,    -5,     0,     4,    -4,    -6,    -7,    -1,     4,     0,     0,     7,     8,     2,    -2,     0,    -4,    -5,    -7,    -8,    -5,    -9,     1,     0,     0,    -3,    -6,     0,    -2,    -3,     7,     3,     1,    -3,    -5,    -1,     2,     0,     1,     9,    13,     4,     0,     5,    -6,    -8,    -7,    -8,    -7,    -9,     7,     0,     1,   -11,    -4,    -1,     1,     6,     6,     1,    -3,    -3,     0,     2,     0,     3,     6,     6,     8,     5,    -1,     1,    -7,    -8,    -2,    -8,    -3,     1,     7,     0,    -1,    -5,     0,    -3,     3,     6,     3,    -3,    -6,    -2,    -3,    -1,    -2,     0,    -2,     1,     9,    -5,     1,     0,    -6,    -6,   -12,    -9,     2,     6,     1,     0,    -1,     1,     2,    -4,     1,    -4,    -5,     0,    -4,    -5,     1,    -1,    -1,     5,    -1,    -3,    -1,   -10,    -4,     2,    -2,    -2,    -5,    -8,     3,    10,     0,     0,    -1,     1,    -3,    -8,    -6,    -3,     0,    -2,    -1,     2,    -4,     0,     1,     3,     1,    -3,    -6,   -10,    -7,    -2,     2,    -8,    -8,   -11,    -4,     0,    -2,     0,     0,     1,    -7,    -7,     1,     1,    -5,    -5,     3,     0,    -3,     0,     4,     3,    -6,   -10,   -10,    -3,    -4,     0,     0,    -2,    -1,     4,     0,    -3,    -2,     0,    -1,    -2,   -11,    -6,     3,    -1,    -4,    -4,    -6,    -5,     4,     4,     3,     4,   -10,    -8,   -11,    -7,    -1,     2,     4,     7,     7,     6,     0,    -5,    -7,    -1,    -1,    -3,   -11,    -7,    -7,   -12,    -8,    -6,    -4,    -3,     0,    -1,     1,     1,    -3,    -6,    -6,     6,     7,     7,     6,     1,    -1,     3,     4,    -4,     2,     1,     0,     2,   -13,   -10,    -3,    -2,    -1,    -1,     1,     4,     4,    -3,    -4,     3,    -2,    -2,     0,     1,     4,    12,     6,     1,     5,     7,     6,    -2,     1,    -1,     0,    -6,   -11,    -2,    -1,     3,    -1,     2,     5,     8,     3,    -1,    -3,    -2,     1,     0,     3,     8,     7,    11,     4,     1,    -1,     3,     2,    -1,     0,     3,     2,    -9,     0,    -2,     2,    -1,     1,    -1,     3,     5,    -3,    -6,    -4,    -2,     4,     3,    -2,     9,     9,    11,     9,    -1,    -2,     4,     3,    -4,     0,     1,     1,    -8,    -6,    -3,     2,    -1,    -2,     5,     2,     2,    -2,    -5,     0,    -5,     5,    -1,     3,    15,    10,     6,     9,     2,     0,     3,     5,    -1,     0,    -1,     1,    -3,    -1,    -6,    -2,     1,     1,    -6,    -1,    -3,     0,     6,     2,     3,    10,     4,     6,     7,     5,     7,     2,    -1,    -6,    -8,    -4,     4,    -1,     0,    -1,     0,    -1,    -6,    -6,    -6,    -1,    -8,    -9,     2,    -5,     1,     1,     1,     5,     3,     8,     2,     3,     1,     5,     2,    -6,    -5,     2,     1,     0,     0,     0,    -1,    -3,    -6,   -11,   -12,   -13,    -8,   -19,   -18,   -15,    -2,     0,    -3,     1,    -7,   -14,   -13,   -16,   -13,   -10,    -4,    -4,    -4,    -4,    -3,     1,     1,     0,     0,    -3,    -8,   -16,   -14,   -10,   -19,   -19,   -10,    -7,   -10,   -12,    -1,    -1,     2,    -7,    -6,    -2,    -3,    -7,    -1,    -1,     1,     1,     0,     0,     1,     1,     0,    -1,    -2,    -2,    -2,     0,    -1,    -2,    -8,    -5,    -2,    -3,    -4,    -2,    -1,    -1,     2,    -1,    -1,     1,    -1,     0,     0,     1,     1,    -1),
		    22 => (    0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     0,    -2,    -3,     2,     2,     0,    -1,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,     1,     1,     1,     0,    -3,    -3,    -7,    -5,    -3,    -4,    -3,    -7,    -2,     0,     0,    -1,    -3,   -12,    -7,    -4,    -4,    -3,     1,     0,     0,     1,     0,    -1,    -1,    -2,    -4,    -2,    -1,    -4,     3,     5,     6,     6,     5,     3,    -3,    -2,    -1,    -4,    -6,    -7,    -7,    -4,    -3,    -1,     1,     5,     1,     0,     1,     1,    -2,    -7,    -7,     6,     5,    -4,    -1,    10,     4,     7,     7,     2,     1,    -2,     0,    -1,    -7,    -5,    -3,     4,     0,    -7,     1,     2,    -1,     0,    -1,     0,     0,    -3,     5,    -2,     2,     5,     3,     8,     5,     4,     5,     4,     0,     1,     2,     4,     2,    -1,    -1,    -5,    -2,    -4,    -3,    -4,    -3,    -3,    -1,     1,     2,     1,     4,     3,    -1,     2,     3,     1,    -1,     0,     0,     1,     2,     2,     7,     2,     5,    -3,    -2,    -1,     2,    -3,    -4,    -3,    -3,    -3,     0,     0,     1,     0,     0,     2,    -2,     1,     5,     2,     1,    -1,     3,     0,     5,    10,     6,     0,     1,     1,    -6,    -4,    -3,    -7,   -12,    -1,    -2,    -2,    -1,     0,     1,    -4,     1,    -1,     4,     4,     3,     4,     0,     1,     0,     2,     1,    -5,     0,    -1,    -2,    -2,    -5,    -6,    -4,   -11,    -4,     1,    -3,    -1,    -4,     3,    -5,    -5,    -1,    -3,    -1,     0,    -2,     0,     5,     2,    -4,    -2,    -1,    -2,    -2,     1,     3,     3,     1,     0,    -7,    -7,    -4,    -4,    -1,    -3,     1,     0,    -1,    -6,    -6,    -8,    -7,    -6,    -9,    -9,    -1,    -1,    -1,    -4,    -5,    -6,     0,    -2,    -1,    -3,     0,    -2,    -3,    -8,    -9,    -7,     1,    -1,     0,     0,    -1,    -8,    -5,    -2,     1,    -4,    -8,    -9,    -6,    -8,    -5,   -11,    -8,    -8,    -3,     2,     3,     3,     2,    -4,   -11,    -4,    -1,    -2,    -1,    -3,    -1,    -4,    -3,    -7,    -5,    -8,    -8,   -15,   -13,   -14,   -13,   -13,   -11,    -8,    -8,   -11,    -6,    -1,    -4,     3,    -1,    -3,    -2,     3,     3,     0,    -8,    -2,     0,    -5,    -6,    -5,   -11,   -10,   -10,   -15,   -12,    -8,    -7,   -10,    -3,     0,    -2,    -4,    -2,    -3,    -2,     3,    -2,    -1,    -2,    -4,   -10,     2,    -6,    -2,    -1,    -5,    -2,    -4,    -8,    -9,    -5,    -1,    -2,    -5,    -5,     4,     9,     7,     4,    -3,    -2,     0,     5,    -1,    -1,    -6,    -3,     0,     4,     4,     4,     2,    -1,    -6,    -5,     6,    -1,    -2,     2,     3,     4,     6,     8,    10,    11,     2,     5,     2,     3,     0,     3,    -1,     0,    -4,     0,     1,     6,     1,     5,     6,     0,    -2,     0,     5,     4,     8,     5,     1,     3,     7,     7,     5,    -1,    -1,     2,     4,     0,    -1,     1,    -1,    -4,     2,    -1,    -2,    -1,     6,     5,     9,    -1,     1,     4,     1,     7,     2,     4,     3,     1,     2,    -1,     3,     0,    -2,     2,     2,     3,     5,     4,     3,     5,     7,     3,     1,    -2,    10,     8,     2,     1,     0,     4,    -2,     2,     3,     6,     0,     6,     0,     4,    -2,     0,    -6,     2,     4,    -2,     4,     3,     1,     0,    -4,     2,    -2,   -10,     6,    -1,     5,    -1,     0,    -3,    -8,    -4,     6,     4,     5,     8,     4,     1,    -5,    -6,     0,     1,     2,     3,    -1,    -4,     1,     4,    -4,     5,     1,     3,     0,    -2,    11,     0,    -3,    -1,   -10,    -2,    -8,     1,     2,     3,     0,    -1,    -7,    -6,    -6,     1,     7,     2,     2,     2,    -4,     0,    -1,     2,    -3,     0,    -3,     7,     9,     0,    -5,     4,    -1,     2,     1,    -7,     0,     7,    -1,    -5,    -2,    -3,    -1,    -3,    -4,    -3,    -4,     3,    -2,     0,    -4,    -2,    -5,     6,    -5,     5,     0,     1,     1,     3,     5,     3,    -1,     0,     0,     2,     0,     4,     0,    -3,    -2,    -3,    -9,   -10,    -5,    -4,     1,    -4,     3,     0,     1,    -6,    -5,   -12,    -1,     1,     1,     3,     9,     4,     1,     1,    -5,    -3,     0,    -2,    -1,    -7,    -4,   -11,   -17,    -3,    -7,     1,     0,    -6,    -5,     3,     1,    -1,    -8,   -13,     0,     1,     0,     1,     2,    -2,    -2,    -7,    -5,    -3,    -2,     0,    -3,    -4,   -12,    -7,   -10,    -8,    -8,    -5,   -13,    -8,    -6,     1,    -5,    -5,    -7,   -13,     0,    -1,    -1,    -7,    -3,    -8,    -5,   -15,    -7,    -8,   -11,   -12,    -8,   -13,   -16,   -14,   -14,   -10,    -5,   -16,   -16,   -10,    -4,    -2,    -9,     1,     2,     0,    -1,     1,     1,     0,    -1,     0,    -3,    -3,    -6,   -10,   -12,    -7,    -5,    -7,    -9,    -8,    -9,   -12,   -13,    -9,   -11,    -9,    -4,    -3,     0,     3,     5,     5,    -1,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -2,    -2,     0,    -1,     0,    -2,    -1,    -3,    -4,    -5,    -4,    -2,    -2,     1,    -4,    -1,    -2,     1,    -1,    -1,    -1,    -1,     1,     0,    -1,     1,    -1,    -1,     0,     1,    -1,    -1,     0,     0,    -2,     0,     0,    -1,    -1,     1,    -1,    -2,    -1,     0,     1,     0,     1,     0),
		    23 => (    0,     0,    -1,     0,     1,    -1,     0,     0,    -1,     0,     0,     1,     0,    -2,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     1,    -1,     1,     0,     0,     1,    -1,     0,     1,     0,     0,     0,     1,    -1,    -1,    -3,    -3,    -4,    -2,    -3,    -3,    -3,    -5,    -4,    -2,    -2,    -1,    -1,    -1,     1,     1,     0,     0,     1,    -1,     1,     1,    -1,    -1,     0,    -1,    -6,    -5,     1,     0,    -4,    -3,    -4,    -6,   -10,    -7,    -5,    -6,    -3,    -2,    -2,    -5,     0,     1,    -1,     0,     1,     0,    -2,     2,    -2,     4,     7,    10,     5,     3,    -4,    -1,     0,     1,    -3,     1,     4,    -2,   -12,    -7,    -3,    -8,    -5,    -8,    -3,    -2,     1,     0,    -1,     2,     1,     1,     5,     5,     1,     3,     8,     6,     0,    -2,     1,     2,     2,    -1,     0,     1,    -7,   -10,   -14,    -5,    -7,   -12,    -7,    -2,    -2,     0,     1,     0,     4,     1,     1,     5,     4,     0,     1,     0,     3,     3,     1,     5,     1,     2,     2,    -4,    -5,    -3,   -12,   -11,   -13,   -11,    -5,    -5,    -3,    -1,     1,     1,     2,     4,     1,     7,     6,     2,     4,     6,     7,    -2,     0,     3,     0,     2,     2,     1,     3,    -2,    -4,   -11,   -12,   -11,    -3,    -3,    -6,    -1,     0,     1,     0,     5,     8,     8,     3,     1,    -1,    -1,     0,    -2,    -3,     3,     1,     0,     5,     3,    -2,    -2,    -9,   -11,   -12,   -13,    -7,    -1,    -6,    -3,    -2,    -1,     2,     3,     0,     6,     6,     4,    -1,    -9,    -4,   -16,   -10,    -3,    -2,     2,     4,     1,     1,     5,    -7,    -9,   -12,   -13,    -9,    -3,    -6,     0,     1,    -2,    -1,    -2,    -2,    -2,    -3,   -12,   -19,   -17,   -10,   -11,    -3,    -2,     4,     5,     3,     2,     0,    -8,   -16,   -12,   -11,    -6,    -5,    -3,    -6,     1,     0,    -3,     2,     0,    -7,   -12,   -21,   -22,   -14,    -5,     5,     0,     1,     4,     6,    -1,     0,     2,    -7,   -13,   -17,   -13,    -3,     0,    -5,    -2,    -4,    -2,     1,    -2,    -1,    -2,   -13,   -14,   -13,   -10,     6,     4,     5,     9,     5,     6,     3,     0,    -8,    -8,    -6,   -10,    -8,    -8,    -5,     0,    -7,    -1,    -3,    -1,     1,    -2,    -3,    -5,    -4,    -1,    -2,     6,     6,     9,     4,     1,     0,     1,    -1,     2,    -6,    -8,    -4,    -6,    -5,    -5,    -3,    -3,    -6,    -1,    -3,    -1,     1,    -1,    -2,    -4,     0,     2,     6,    14,     9,     3,     0,    -4,     0,    -1,     6,     1,     0,    -7,    -3,    -2,     0,    -1,    -4,    -1,    -7,    -6,    -4,    -3,     0,     1,     0,    -5,     1,    -3,    -2,     0,     3,    -1,    -1,    -4,    -4,     0,     0,    -4,    -2,    -3,    -3,     3,     0,     6,     1,     3,     0,   -13,    -1,    -3,    -2,     3,     0,    -3,    -1,    -1,    -2,   -10,    -4,    -7,    -4,    -7,    -3,     0,     0,    -8,     0,     3,    -1,    -1,    -1,     6,     2,     3,     5,    -7,    -1,    -1,     0,     0,     1,    -4,    -4,    -3,    -7,   -12,    -3,    -7,    -8,   -13,   -18,   -11,    -4,    -5,    -1,     3,     0,     3,     1,     6,     7,     5,     3,   -13,   -11,    -3,    -1,     2,     3,     3,    -4,    -3,    -2,     1,     6,     1,    -2,   -12,   -16,   -11,   -12,    -6,     0,     2,    -5,    -6,    -1,     2,     3,    -5,    -3,   -13,    -2,    -3,    -1,     2,    -1,     6,     3,     4,     9,    -4,    10,     2,    -2,    -1,    -2,    -5,    -4,    -3,     4,    -3,    -3,     0,     1,     1,    -1,    -6,    -5,    -7,    -4,    -3,    -1,     0,    -7,     2,     3,     3,    -2,    -2,     3,    -2,    -2,     3,     6,     5,    -2,    -1,    -6,    -2,    -1,     0,    -3,    -5,     0,    -2,     1,    -4,    -6,    -3,     1,    -1,    -6,     2,    -4,     1,     3,    -1,     2,     3,     0,    -4,    -3,    -4,     0,    -3,     0,     0,     1,    -4,     1,    -7,    -5,    -2,     2,    -2,    -5,    -1,    -1,     0,     2,     0,     0,     0,     1,     2,     2,     3,     0,     2,     4,     1,    -4,    -4,     1,    -4,    -1,     1,    -2,    -5,    -2,    -2,    -4,    -1,    -3,     0,     0,     0,     0,     4,     8,     2,     5,     1,     0,     2,     2,     1,     0,     0,     0,     0,    -5,    -2,    -2,     0,    -2,    -1,     2,     2,     2,    -5,     0,    -1,     0,     1,     2,    10,    10,     2,     1,     5,     2,     1,     1,     0,    -3,     4,    -2,     0,    -1,    -3,     2,     0,     1,     1,    -4,     1,     4,     1,    -1,     0,     0,     0,    -3,     2,    -1,    -1,    -7,     4,    -3,    -3,    -3,     2,     0,    -1,    -1,    -3,    -3,    -3,    -1,    -4,    -3,    -6,    -7,    -5,    -3,    -1,     0,    -1,    -1,     0,     1,    -2,    -1,    -2,     4,     6,     6,    -1,    -2,    -5,   -12,    -5,    -6,    -4,     3,     1,     0,     5,    -1,    -7,    -9,    -6,     0,    -2,    -1,    -1,     0,    -1,     1,    -2,    -3,    -4,    -3,    -1,    -3,    -5,    -3,    -4,    -7,    -7,    -9,     0,     2,    -2,    -1,     1,    -3,    -4,    -6,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,    -1,     0,     0,    -1,    -2,    -7,    -4,    -8,     0,    -2,    -1,     1,    -1,     1,    -2,    -1,    -2,    -1,     1,    -1,     1,     0),
		    24 => (    0,     0,    -1,     1,     1,    -1,     1,     0,    -1,     0,    -1,     0,    -4,    -3,    -2,    -2,    -1,     1,     0,     0,     1,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,    -3,    -4,    -2,    -5,    -7,    -3,   -10,    -2,     3,    -4,    -7,    -4,    -5,    -2,    -4,    -1,    -2,    -4,    -1,     0,     0,    -1,    -1,     0,    -1,   -11,   -12,    -3,    -4,    -9,    -9,    -6,    -8,   -11,   -11,    -4,    -1,    -8,    -7,    -6,    -4,    -8,    -4,    -2,    -1,     0,     0,    -1,     1,     0,     1,     0,    -1,   -10,    -9,     0,    -4,    -9,    -8,   -11,    -1,    -6,   -12,    -7,     0,     0,     4,     3,     3,     0,    -3,     0,     4,     3,     5,    -3,     0,    -1,    -1,     1,     0,    -2,     2,    -7,    -1,    -3,    -3,    -1,    -1,     1,    -3,     3,    -5,    -1,     2,    -1,    -4,    -6,     5,     4,     9,    11,     6,     1,    -5,    -1,    -1,     0,    -2,     3,    -4,    -1,    -3,    -5,    -5,    -3,     0,     3,     1,    -3,    -4,    -4,    -8,    -9,    -5,    -2,     3,     0,     0,     2,     1,     0,     1,     1,    -1,    -1,     1,    -2,    -3,     2,    -4,    -7,    -2,     3,     2,    -4,    -5,    -1,    -4,    -3,   -18,   -23,   -10,    -1,     6,     2,     4,     1,    -6,    -2,     1,    -5,     0,    -1,    -1,    -4,    -2,    -3,    -4,    -3,     2,     1,     0,    -1,     1,     1,    -1,   -12,   -21,   -19,    -5,     3,     3,     5,    10,     7,    -4,    -7,     6,    -4,    -2,    -4,     3,    -2,    -6,    -5,    -3,    -2,    -2,    -6,    -1,    -3,    -2,     3,    -4,   -10,   -18,   -14,    -3,     3,     1,     1,     6,     5,    -3,    -1,     3,    -6,     0,    -2,     4,    -4,    -4,    -3,    -2,    -4,     1,     1,    -1,    -3,     2,     2,    -7,   -16,   -19,   -11,    -2,     8,     4,    -1,     5,     3,     1,    -1,    -4,    -2,     1,     0,     3,     5,    -3,    -3,    -5,    -3,     1,     0,    -1,     2,     3,    -1,   -14,   -18,   -12,    -6,     7,     6,     1,    -1,     0,     2,     1,    -2,    -2,    -3,    -1,    -2,    -2,     1,    -3,    -3,    -2,    -3,     0,    -3,     2,     2,    -1,    -2,    -6,   -11,    -8,    -1,     2,     7,    -3,     0,     0,     2,    -1,    -3,    -4,    -6,     0,     0,     3,    -4,    -3,    -5,    -3,     1,     1,    -1,     0,     0,     2,    -4,   -12,    -7,    -8,    -2,     6,     3,     1,    -3,    -1,     1,    -5,    -6,    -4,    -6,    -1,    -2,    -2,    -4,    -2,     0,    -1,    -1,     3,    -1,    -1,    -3,     0,    -5,    -6,    -5,    -5,     0,    -3,    -2,    -1,     3,     3,    -1,    -9,    -1,    -4,     0,     0,     0,    -5,     8,     1,    10,    -2,     2,    -6,     3,     1,     0,    -4,    -6,    -3,    -4,    -3,     0,    -5,     2,    -1,    -2,    -1,    -3,    -3,    -7,     0,    -1,     0,     1,    13,     7,     2,     3,    -3,    -1,    -1,     6,     5,     1,    -4,    -2,    -5,    -5,    -5,     3,    -1,     0,    -1,    -5,     3,    -2,   -12,    -7,    -5,    -2,     1,     1,     4,     0,   -10,    -2,     4,     6,    10,     6,    11,    -1,    -3,     0,    -4,    -1,     1,    -1,     0,     0,     1,     0,     4,    -7,    -7,    -7,    -3,    -4,    -1,    -1,    -1,    -6,    -6,    -3,     2,     7,     9,     5,     7,     3,    -4,    -1,     1,     0,    -1,     1,     8,     5,     3,     5,     3,     0,    -8,    -5,     3,    -4,    -1,     1,     0,   -13,     2,     1,    -1,     2,     1,     1,     1,     1,     5,    -1,     2,     4,     2,     4,     5,     4,     2,     3,     2,    -5,    -9,    -5,     0,    -1,     0,     0,    -1,    -8,    -2,     4,     5,     1,    -1,     1,    -2,    -3,    -5,    -2,     0,     4,     0,     0,     2,     5,    -1,    -6,    -3,    -5,    -1,    -9,    -3,    -1,    -1,    -1,     1,    -9,    -8,    -2,    -5,    -4,    -5,    -8,    -9,    -8,    -2,    -4,     2,    -1,    -4,    -2,    -5,     6,     2,    -3,     1,     1,     2,    -7,    -3,     0,     0,     0,    -2,    -8,    -2,    -3,    -4,    -2,    -7,   -14,   -14,    -5,    -4,    -2,     0,    -3,    -1,    -1,    -1,     3,    -1,    -3,     4,     4,    -1,    -8,    -4,    -1,    -1,     0,    -1,    -6,    -7,    -4,    -6,    -9,   -11,   -10,   -11,     5,    -1,    -3,    -4,    -2,     0,    -3,    -3,     1,    -4,     4,     4,     6,    -3,     1,    -2,    -1,    -1,    -1,    -1,    -2,    -5,    -3,    -6,    -8,    -3,    -3,     0,     4,     2,    -2,    -1,    -4,     2,    -1,    -1,    -2,    -7,     4,     1,     1,    -5,    -3,    -2,    -1,     0,     1,     0,    -1,    -3,     1,    -1,    -5,    -2,     0,    -1,    -2,    -1,     0,    -4,    -1,     3,     3,    -6,    -3,    -8,     0,     5,     3,    -6,    -4,    -1,     0,    -1,     1,    -3,     1,    -1,    -1,    -2,     0,     1,    -2,     0,    -3,     0,     1,    -8,     0,    -3,    -6,     1,    -1,    -7,    -8,    -2,     1,    -4,    -1,    -1,    -1,     1,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     3,     3,     2,     3,     2,   -13,    -9,    -3,    -4,    -6,    -1,    -8,    -9,    -8,    -3,    -2,     0,     0,     1,     1,     1,    -1,    -1,     0,     0,    -3,    -3,    -4,    -2,    -3,    -3,    -1,     0,     0,    -1,    -5,    -7,    -1,    -3,    -2,    -5,    -5,     0,     0,    -1,    -1,     0),
		    25 => (   -1,     1,     1,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     1,    -1,    -1,    -1,     1,    -1,    -1,     0,     0,    -1,     1,     1,    -1,     1,     0,     0,     0,     1,    -1,    -2,    -1,    -2,    -1,    -3,    -3,    -4,    -4,    -2,     0,     0,     0,     0,     1,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -2,     0,    -3,    -3,    -2,    -1,    -4,    -1,    -3,     5,     4,    -4,     2,    -1,    -1,    -1,    -2,    -3,    -1,     1,     0,    -1,    -1,     1,     3,    -4,    -2,    -3,    -1,    -1,    -2,    -4,    -5,    -8,    -2,     2,     1,     4,     4,    -3,     2,     4,     2,    -5,    -4,    -2,     4,     1,     1,     0,    -2,     2,    -1,     1,    -1,    -1,    -1,    -1,    -4,   -11,    -8,    -9,     0,     4,    -3,     2,     4,     0,    -3,    -1,    -3,     2,     3,     2,     1,    -7,     0,     0,    -3,     1,    -1,    -1,    -2,    -2,    -2,    -4,    -9,   -11,    -5,    -4,    -3,    -2,     1,    -1,    -2,     0,     0,    -5,    -2,     5,     2,     7,    -2,    -4,     0,     1,     1,    -1,    -2,    -4,     1,    -3,    -2,    -4,    -5,   -15,    -2,    -2,     5,     0,    -1,    -4,     0,     4,     2,    -1,     6,     5,     6,     6,     0,     0,     0,     0,     0,    -2,    -2,    -2,     1,     0,    -3,   -11,    -2,   -11,    -4,    -1,    -1,     1,     2,     1,    -3,     0,    -1,     2,     5,     5,     4,     9,     2,     1,    -1,    -4,    -4,    -2,    -1,    -1,     3,    -3,    -4,    -3,    -1,     0,     6,    -1,    -2,    -1,    -3,    -3,     1,     1,    -3,     3,     5,     8,     7,     8,     0,     4,    -1,     0,    -5,    -3,    -1,     2,    -3,    -3,     0,    -1,     3,    -2,     3,    -4,     0,    -1,    -3,     1,    -1,    -2,    -1,    -1,     5,     8,    13,     8,     0,     6,     0,    -2,    -1,     0,    -2,     0,     0,     0,    -2,    -7,     3,    -3,     2,     3,     6,     0,    -2,    -4,     3,     3,     4,    -4,     2,     2,     8,     5,     5,     5,    -1,     0,    -2,    -1,    -1,     0,     2,    -1,     0,    -2,     3,    -1,     0,    -1,    -3,    -3,    -9,    -7,    -7,     1,    -9,    -4,    -1,     1,    -1,     2,     7,     2,     1,     1,     1,    -1,    -3,    -1,     2,     1,     4,     0,     1,    -2,     1,     4,    -3,    -9,   -16,   -18,   -16,   -17,   -16,   -16,   -11,    -5,    -5,     0,     4,    -7,    -1,    -2,     1,     0,    -3,    -1,     4,     3,    -1,     1,     2,    -3,     2,     1,     1,    -7,   -10,   -13,   -17,   -13,   -15,   -14,   -14,    -8,     0,     0,     6,    -3,     2,     0,    -2,     0,    -2,    -3,    -1,     0,    -1,    -3,     3,    -4,    -1,     0,    -2,    -3,    -6,   -13,   -16,   -13,   -11,    -9,    -7,    -6,     1,     1,     0,    -3,     1,    -2,    -3,     0,    -2,    -7,    -6,    -6,    -1,    -1,    -1,    -1,     4,    -3,     1,     2,    -1,     0,    -7,   -10,   -12,    -9,    -7,    -4,    -2,     0,    -1,    -2,     1,    -2,    -3,     4,    -2,    -5,    -9,   -10,    -4,    -5,    -3,    -2,     0,     1,     2,     0,     2,     1,    -6,    -9,   -13,    -9,    -6,    -6,    -2,    -2,    -4,    -1,     1,    -1,    -7,     8,     2,    -5,    -9,   -10,    -4,    -7,    -8,    -1,     3,    -1,     1,    -1,     3,     6,    -6,    -7,   -10,    -7,    -5,    -7,    -6,    -2,    -4,    -4,     0,    -1,     0,     9,     7,     4,     0,    -1,    -7,    -8,    -6,    -6,    -3,     1,    -1,    -2,    -3,    -3,    -5,    -3,   -10,    -5,    -4,    -4,    -2,    -2,    -4,    -1,     0,    -1,     2,     1,     6,     5,     6,     8,    -1,    -5,     0,    -4,    -5,     3,    -4,     0,     0,     5,    -6,    -4,    -5,    -3,    -3,    -4,    -1,    -6,    -3,    -3,    -1,    -1,     0,     1,    -2,     4,     5,     8,     4,     1,    -1,     1,     2,     3,     1,     1,     5,     0,    -2,    -6,    -4,    -3,    -2,     0,    -1,     0,    -2,     0,     0,    -1,     0,    -2,    -4,    -4,    -5,     4,     5,     2,    -1,     3,     3,     1,     5,     3,     1,    -2,    -1,    -3,    -4,    -1,    -1,    -2,     0,     0,    -1,     0,     0,     1,    -3,     4,    -1,    -4,     1,     2,     0,     0,     0,     6,     4,    -1,     0,     1,    -4,     0,    -1,    -4,    -4,     0,     0,    -1,     1,    -2,    -1,    -1,    -1,    -1,     3,     3,     3,    -2,     0,     7,     7,     6,     3,     7,     4,     1,     3,     0,     0,     4,     0,    -1,    -2,     0,     0,    -1,     1,    -2,    -5,     0,     0,     0,    -2,    -1,     0,    -4,     1,     5,     1,     8,     6,     5,     5,     2,     1,    -3,    -4,     2,    -2,     1,     0,    -1,     0,    -1,    -1,    -7,    -2,     1,    -1,     0,     1,     0,    -6,    -5,    -1,    -4,    -3,     4,    -1,    -2,    -3,     0,    -7,    -6,    -4,    -3,     5,     2,     0,    -2,    -1,    -1,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -3,    -9,    -9,    -4,    -2,     2,     4,     6,     2,    -7,    -9,    -2,     0,    -2,     0,     1,     1,     1,    -3,     1,     0,     0,     0,     1,     1,     0,     0,    -2,     0,    -2,     0,    -1,    -1,     0,     1,     1,    -1,    -2,     0,     0,     1,     0,    -1,     0,    -1,    -4,     0,     0,    -1,    -1,     0),
		    26 => (    0,     0,     1,     0,    -1,    -1,     0,     1,     0,     0,     0,    -1,     5,     4,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     1,     0,     1,    -1,    -1,     1,     0,     0,    -1,    -1,     3,     5,     6,     3,    11,    10,     2,     4,    -5,     1,    -2,     1,     4,     4,    13,     5,     3,     5,     1,     0,     1,    -1,    -1,     0,     2,     3,     7,     9,     4,     6,    12,    10,     5,     5,    -9,    -6,     0,    -1,    -1,     6,     3,     0,     4,     4,     7,     4,     1,    -5,    -1,     0,     1,     0,   -10,    -2,     0,     9,     8,     2,     1,     1,    -1,    -7,    -9,    -2,     4,     3,    -1,     4,     4,     3,     0,    -3,     1,     9,     5,    -7,    -6,     1,     0,     1,    -9,     0,     0,     7,    -1,    -2,     5,     7,    -2,    -5,   -15,    -4,     0,    -4,     2,    -1,    -5,     0,    -2,     4,     5,     8,    -1,   -10,     5,     9,     1,    -1,    -8,    -6,     3,    -3,    -9,     5,     3,     1,    -6,   -13,    -5,    -3,     0,     0,    -7,    -1,    -7,    -4,     0,     0,     1,     6,     1,    -5,    12,     8,     0,    -1,     3,    -2,     2,    -3,    -6,     3,    -2,    -9,    -5,    -6,     1,    -7,    -6,    -1,    -3,    -2,    -1,     1,    -2,    -4,     5,     0,     3,    -4,     3,     5,     0,     0,     0,    -4,     2,    -1,    -3,    -1,    -4,    -7,    -7,    -1,    -1,    -3,    -2,    -4,    -1,    -2,    -5,    -2,    -2,    -1,     0,     1,     1,     0,     2,     4,    -1,     1,    -5,    -4,     3,    -4,    -6,    -6,    -4,    -8,    -1,    -2,    -4,    -3,    -5,    -6,    -4,    -5,   -11,     0,    -9,     0,    -2,    -2,     3,   -13,    -2,    -9,     1,     0,    -6,     2,     1,   -10,    -3,    -7,    -6,     0,    -1,     1,    -4,    -3,    -2,    -8,   -13,   -12,   -13,    -7,    -7,    -7,   -18,    -6,     2,    -1,    -3,    -9,    -1,    -1,    -7,    -6,    -4,    -7,   -10,   -10,    -6,     3,    -4,    -2,     1,    -1,    -5,    -6,    -9,    -7,    -5,    -3,    -4,    -3,    -6,     5,     5,     9,    -5,   -11,     1,    -1,     0,    -4,    -3,    -3,    -6,    -1,    -1,     1,     4,     3,     1,     6,     2,    -2,    -1,    -3,    -7,    -9,     2,    -5,    -4,     1,     1,    -2,    -6,    -3,     1,     0,    -1,    -5,    -4,    -7,     0,     3,     6,     8,     8,     3,     1,     2,    -1,    -2,     2,    -1,    -6,   -12,    -9,    -2,     4,     9,     6,    -1,   -10,    -2,     1,     0,    -2,    -4,    -4,    -1,     8,     4,     1,     5,     8,     2,     1,    -3,    -2,     0,     0,     1,    -5,    -4,    -6,    -4,     2,     9,     6,     3,    -3,     1,     0,     1,    -1,    -8,    -6,     5,     2,     3,     6,     8,     2,     5,    -1,    -5,    -1,    -1,     2,    -2,    -2,    -1,    -2,     3,     7,     5,     2,     3,    -8,    -5,     0,     0,    -3,    -9,    -8,     6,     7,     8,    11,    10,     6,     5,     5,     1,    -2,    -4,    -1,     0,    -1,     2,     1,    -2,     7,     6,    -7,    -3,   -10,    -5,     0,     0,     0,    -8,    -1,     5,     4,     8,    13,    12,     9,     8,     8,     1,     1,    -1,     3,    -2,    -2,     6,     3,     1,     5,     7,    -4,    -7,   -10,    -6,    -1,    -1,     0,    -7,    -7,     3,     3,     6,     4,     4,    10,     3,     8,    10,     1,    -1,    -1,    -3,    -1,     3,     2,     5,    -1,    -1,    -2,    -7,   -11,    -9,     1,     0,    -1,    -1,    -4,    -3,    -1,     4,    -3,     3,     3,     0,     7,    10,     3,    -6,     0,     0,    -4,    -6,     0,    -2,    -3,    -4,   -12,    -8,    -6,    -6,     1,     0,    -6,     1,     0,    -9,    -6,    -2,    -5,     0,    -2,     4,     3,     1,     0,    -2,    -2,     3,    -3,    -3,    -2,    -1,    -1,    -1,    -5,     2,    -4,    -7,     1,    -2,     0,    -9,     2,    -6,    -6,    -5,    -4,     1,    -2,    -1,    -2,    -5,     4,    -1,    -6,    -4,    -1,    -3,    -1,    -3,     5,     0,     4,     8,    -2,     0,    -1,     0,    -3,    -4,    -4,    -3,    -6,    -2,    -1,     2,     1,    -5,     7,     7,     1,    -4,    -1,     0,     1,     4,    -1,     0,     5,     6,     5,     2,    -1,    -2,     1,    -1,     0,    -3,    -4,   -11,   -11,    -7,     3,    -4,     0,    -3,     5,     6,     2,     3,     5,     1,     1,     2,    -2,     4,    -2,     0,    -4,    -9,    -1,    -2,     1,     0,     1,    -1,    -5,    -9,   -10,    -8,    -5,    -2,    -3,     0,    -3,     1,    -1,     2,    -4,     0,     5,     7,     0,    -6,    -9,    -8,    -7,    -7,   -10,     0,     1,     0,     0,     0,    -3,    -3,    -1,    -7,    -7,   -10,   -11,    -8,    -3,    -5,     1,     3,     5,     5,     1,   -12,    -5,   -12,    -7,    -6,    -4,    -5,     0,     0,     1,     0,     0,    -1,     0,    -2,    -2,    -6,    -3,    -4,    -6,     0,     6,     0,    -5,    -2,    -6,    -5,    -2,    -5,    -9,    -3,    -3,    -3,    -2,     0,     0,    -1,     1,     0,     1,    -1,     0,    -2,    -3,    -1,     0,    -2,    -4,    -3,    -1,    -1,     0,    -2,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     1,     0,     1,    -1,     0,    -1,     1,    -1,    -1,     1,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -2,     0,    -1,     0,    -1,     0,     0),
		    27 => (    1,     0,     1,     0,     1,     1,     0,     1,     0,    -1,    -1,     1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,     0,     0,    -1,     0,    -1,     1,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,    -6,    -4,    -5,     0,    -1,    -2,    -1,     1,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     1,     1,    -2,    -2,     0,     0,    -2,    -1,    -1,    -2,    -3,    -6,    -4,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,    -2,     0,     1,    -1,     0,     1,     1,    -1,     0,    -3,    -3,    -2,    -2,    -3,    -5,    -5,    -3,    -6,    -5,    -2,    -1,    -2,    -3,    -3,     0,    -3,     0,    -4,    -3,    -2,    -1,     0,     1,     1,    -1,     1,     0,     0,    -7,     0,    -2,    -6,    -6,    -8,   -11,   -10,    -9,   -11,    -8,    -9,    -7,    -3,    -3,    -2,     0,    -5,    -7,    -5,    -4,    -3,    -2,     1,     0,     1,     1,    -4,     1,     2,    -2,    -6,     5,     4,    -5,    -4,    -7,    -6,    -5,    -7,   -10,   -20,   -24,   -16,   -11,    -4,     0,   -11,    -8,    -8,    -4,     0,    -1,     1,     1,    11,     8,     7,    -3,    -6,     7,    -1,    -4,    -1,     3,     4,     0,    -7,    -1,     1,     4,    -1,     3,    10,     0,   -14,   -10,   -10,    -7,     0,    -1,     8,     0,     8,     8,    -3,     0,     1,     1,     3,     6,     5,     4,     0,    -1,    -1,     2,     2,     1,     6,     4,     5,     8,     9,    -1,    -4,    -8,    -4,    -6,    10,     2,     6,     3,    -5,    -4,     2,     3,     1,     1,     2,     2,     2,     0,     2,     3,    -1,     2,     2,     2,     4,     3,     2,     3,    -5,   -11,    -2,    -1,     6,    -3,     1,     3,     3,     0,     4,     5,     6,     6,     4,     6,     0,    -2,    -1,    -2,     1,     0,     5,     2,     9,     2,     0,    -1,    -2,   -10,     0,     0,     4,     0,    -4,     7,     5,     1,     2,     3,     3,     1,     7,     1,    -2,    -9,    -5,     1,     7,    -1,     4,     5,     3,     2,    -3,    -5,    -6,    -6,     1,     0,    -3,     8,    -1,     6,     2,     2,     5,     0,     1,     8,    10,    -1,   -13,   -19,    -3,     2,     4,    -1,    -1,     5,    -2,    -1,    -2,     2,    -9,    -2,     1,     0,     4,     1,     1,     1,     5,    -4,     3,     1,     0,     5,    -1,   -11,   -29,   -19,    -2,     2,    -1,     2,    -8,    -1,     1,    -1,   -10,    -1,    -3,    -3,     1,    -1,     5,     0,    -1,    -4,    -1,     2,     4,     5,     4,     3,     0,   -18,   -30,   -11,    -4,     1,     0,    -6,    -8,     0,     1,    -8,   -10,    -4,    -2,    -3,    -2,     0,     1,     4,     1,    -1,    -3,     5,     3,     2,     2,     6,    -9,   -25,   -26,     0,    -1,     1,    -2,    -7,    -1,     0,    -4,    -4,     1,     4,    -3,    -2,     0,     0,    -1,     4,    -1,    -4,     1,     0,     5,     0,    -1,     0,   -17,   -28,    -7,    -3,    -6,    -1,    -3,    -2,    -1,     2,    -2,    -1,     2,     4,    -1,     0,    -1,     1,     0,     4,    -4,    -5,     0,    -3,     0,    -1,    -7,    -8,   -16,    -9,    -3,    -4,    -3,    -5,    -2,    -4,    -2,     1,    -1,    -3,    -8,    -9,    -4,     0,    -3,     1,     0,     0,    -3,    -4,    -3,   -11,    -6,    -5,    -4,    -3,    -2,    -9,    -7,    -4,    -3,     1,     0,     4,     2,    -1,     1,     0,    -8,   -11,    -5,     0,    -5,     1,    -1,     6,    -7,    -8,    -1,    -5,    -5,    -6,    -1,    -2,    -6,    -8,    -5,    -1,    -5,     1,     3,     3,     2,     0,    -7,    -3,    -5,   -12,    -9,     0,    -3,     1,     3,     1,    -8,     1,     4,    -1,    -9,     5,     5,    -3,     0,    -3,    -2,     2,    -2,    -2,    -4,    -4,    -1,    -1,    -5,     2,    -5,    -6,    -3,    -1,    -1,     0,     6,    -2,    -2,    -3,    -9,    -7,    -2,    -1,     1,     1,    -2,     6,    -3,    -1,    -1,    -6,    -4,    -5,     0,    -5,   -13,   -10,    -9,    -8,    -1,    -3,     1,     0,     1,    -1,    -5,    -8,    -7,    -7,   -10,    -2,    -4,     1,     5,     2,    -1,     1,    -2,    -2,    -5,    -2,     1,    -1,     3,     2,    -4,     1,    -1,    -3,     0,     0,     0,    -1,    -4,    -6,     2,    -7,    -5,    -2,     1,     0,    -3,    -2,     1,    -1,     1,    -3,    -3,     2,     2,    -5,    -2,    -3,    -4,    -2,     0,   -10,     0,     0,     1,    -2,    -5,     1,     6,     2,     1,    -4,     2,     4,    -3,    -7,     1,    -3,     0,     1,     1,    -3,    -1,    -5,     0,    -6,    -4,    -2,    -1,    -5,    -1,     0,    -1,     3,     7,    14,     8,    -1,    -2,     0,    -4,     5,    -3,    -2,    -8,   -10,     1,    -2,    -1,    -3,    -1,    -4,     1,    -3,    -2,     0,    -2,     0,     1,     1,     1,    -6,     5,     1,    -8,    -6,    -1,     2,     0,    -6,    -3,     5,    -1,     4,     2,     0,     1,     1,    -2,     1,     8,     4,    -5,    -1,     0,     1,     0,     0,     0,    -1,    -4,    -6,    -9,    -4,     5,     7,    -1,    -7,    -6,    -4,     2,     0,     4,     2,    -3,     0,     6,     4,    -1,    -1,    -2,    -2,    -1,     0,    -1,     0,    -1,     0,     0,     5,     6,     2,     0,     3,     3,     2,     1,     1,     6,     6,    -1,     0,     6,     2,     5,     4,     1,     1,     8,    -1,    -1,    -1,     0),
		    28 => (    0,    -1,    -1,     0,     0,     1,    -1,     0,     0,    -1,     1,    -1,    -1,    -1,     0,    -1,     1,     1,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     1,     0,     1,     0,     0,     1,    -1,    -1,    -4,    -4,    -5,    -5,   -10,    -8,   -10,    -1,    -2,    -1,     2,     0,     1,     1,     0,     0,    -1,     1,     0,     0,    -1,    -2,    -1,    -2,     0,    -4,    -8,   -14,   -13,    -6,    -5,    -2,   -11,   -11,   -10,    -4,    -8,    -5,    -5,    -7,    -5,    -2,    -2,     1,     0,     1,    -1,    -4,    -3,    -2,    -8,   -14,   -17,   -20,   -22,   -14,   -12,    -3,     6,    -4,    -1,    -3,    -7,   -14,   -13,    -3,     2,     5,     6,     4,     0,    -3,     0,     0,    -5,    -3,    -8,   -10,   -17,    -8,    -7,    -2,    -3,     0,    -6,    -5,     3,     3,     0,    -2,    -4,    -5,     2,     4,    -5,    -4,    -4,     3,    -5,     6,    -1,     1,    -1,    -7,    -6,    -5,   -14,     0,    -1,     2,     0,    -5,    -1,    -2,     0,     3,    -4,    -2,    -1,    -7,    -1,    -1,     5,     4,    -2,     9,     8,    -6,     2,     0,     0,    -2,   -11,    -4,    -6,     4,     0,     0,    -1,    -1,     2,     2,    -4,    -3,    -2,     2,    -1,     4,    -3,     2,     4,     5,     7,     2,    -5,    -6,     0,    -1,    -4,    -3,   -10,     1,     2,    -1,     4,     1,    -1,     3,    -1,    -2,    -4,    -6,     1,     1,     0,     1,     0,    -5,     5,     8,     3,    -2,    -4,    -8,     1,    -4,    -5,    -9,    -1,    -1,    -3,     2,     3,    -1,     4,    -1,    -5,    -3,     2,    -3,    -9,    -6,     2,     4,     0,     0,    -1,     6,     3,     6,    -5,     4,     4,    -1,    -4,    -9,    -1,    -8,    -2,    -1,    -3,     4,    -1,    -3,    -2,    -4,    -2,    -6,    -7,    -3,     3,    -6,     5,    -2,    -3,    -1,     5,     7,     0,     3,    -4,    -1,    -1,   -13,   -11,     2,    -1,    -2,     3,     0,     4,    -3,    -1,    -2,    -4,     8,     2,    -2,    -3,    -2,     2,     1,     0,     1,    10,     6,    -6,     2,    -2,     0,    -1,    -8,     8,     3,     2,    -2,    -1,     3,    -1,     1,     0,     2,     4,     8,     9,     1,    -1,    -2,    -2,     3,     3,    -1,     3,    13,    12,     7,    -5,     0,     0,    -5,     9,     6,     4,    -3,     1,     0,    -6,    -6,     5,     9,     9,     5,     6,     3,     7,    -2,     8,     2,     0,    -8,    -2,     3,     9,     4,    -6,     0,     0,    -3,    11,     1,     1,    -2,     3,    -4,     1,     2,     8,     5,     8,     7,     7,     4,     4,     5,     6,    -2,    -8,     1,    -4,    -8,    -1,    -3,     0,    -1,    -1,    -1,     8,     2,     1,     2,    -4,    -6,    -1,    10,     6,     5,     8,     4,     0,     4,     3,     4,     3,    -8,   -10,    -6,    -4,    -7,     8,    -8,     0,    -1,     0,    -3,     0,   -11,    -8,    -3,     2,     1,     6,     7,     5,     4,     8,     5,     3,     5,     4,    -1,    -4,    -6,    -8,     1,     2,    -9,     9,   -18,    -6,    -1,    -1,    -2,    -1,    -2,    -2,     2,     1,     2,     3,    10,     3,     9,    -1,     2,     2,     8,    -5,    -4,     1,    -7,    -3,    -1,     8,   -10,     4,   -15,    -7,    -1,    -1,    -2,    -6,     6,     3,    10,    -2,    -4,     4,     7,    10,     9,    10,     7,     0,     9,     0,    -6,    -3,    -5,    -3,     2,    12,     4,    -7,    -4,    -9,    -1,    -2,    -3,    -8,     7,    -1,    -2,     1,    -2,     1,     4,     6,    12,    15,     7,     5,    -2,    -4,    -3,    -7,    -2,    -4,    -2,     3,    -2,    -9,    -5,    -3,    -1,    -1,    -9,    -4,    -4,     0,     3,    -2,     3,     2,     2,    -5,     1,     7,     2,    -4,    -9,    -5,     0,    -2,     1,    -2,     3,    -4,    -2,   -11,   -14,    -3,     0,     0,    -4,     0,    -1,     1,     3,     1,    -7,    -2,    -3,    -5,    -4,    -4,    -2,    -3,    -2,    -5,     0,    -2,     3,    -3,     5,    -5,    -4,    -8,    -8,     0,    -4,    -1,    -6,     1,    -2,     1,    -1,    -4,    -6,     0,    -7,   -10,    -8,    -6,    -5,    -6,    -6,     5,     6,    -3,     0,    -2,    -1,    -5,   -13,    -8,   -14,    -2,    -3,    -2,    -3,    -1,     2,    -6,    -2,     0,     1,    -1,    -3,    -6,    -4,    -7,    -6,    -1,    -5,    -7,    -2,    -3,    -1,     5,    -5,    -7,   -10,     2,    -6,    -1,    -1,     0,    -4,     2,     1,     0,    -7,     0,     2,     4,    -5,    -4,    -5,    -1,    -6,    -1,    -1,     0,     0,     4,     7,    -5,     2,     4,    -5,     2,    -8,    -1,     1,     1,    -4,    -3,   -14,   -11,    -9,   -13,    -7,    -1,     0,    -2,     0,    -1,    -5,    -3,    -7,    -9,    -5,     6,    -2,    -8,    -3,     1,    -3,    -5,    -2,    -1,     0,    -1,    -4,    -3,    -3,    -1,     6,     5,    -2,    -1,     8,     1,    -8,    -4,    -1,     3,     5,     0,     2,    -6,    -3,    -5,    -8,    -6,    -9,    -6,    -4,     0,     0,     0,     1,    -4,    -4,    -8,   -10,   -10,   -12,   -17,   -14,    -7,    -6,    -6,    -7,   -17,    -9,    -6,    -7,   -14,   -10,    -6,    -4,    -4,     0,    -1,     0,    -1,     0,     1,     1,    -1,     0,    -1,    -1,    -4,    -8,    -8,    -5,    -1,    -3,    -6,    -7,    -9,    -6,    -6,    -4,    -5,     0,    -1,    -1,     0,     0,     0,     1,    -1),
		    29 => (    1,     0,     0,    -1,     0,     0,    -1,     1,     0,     1,    -1,     0,     1,     1,    -1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,     1,     0,     0,     1,    -1,     0,    -2,    -3,    -2,     0,    -1,    -4,    -5,    -4,    -3,     1,    -2,     0,     0,     1,    -1,     0,    -1,     0,     1,    -1,    -2,    -2,     0,     0,    -2,    -1,    -2,    -2,    -4,     0,     0,    -7,    -5,    -4,    -1,    -1,    -1,    -9,    -3,    -6,    -4,    -2,    -1,     0,     1,     0,     0,     1,    -2,    -3,    -8,    -7,    -7,    -9,    -8,   -15,   -15,   -10,   -12,   -22,    -9,   -11,   -16,   -12,    -8,   -13,   -14,    -9,    -5,    -3,    -2,    -1,     0,     1,    -1,    -3,    -3,    -4,   -13,   -18,    -7,    -8,   -10,    -5,    -3,    -2,    -2,    -4,     2,    -2,    -7,    -2,   -18,   -16,    -5,    -7,    -4,    -3,    -9,    -6,    -1,     0,    -1,    -1,    -2,    -1,    -5,    -6,    -6,    -3,     1,     1,     5,     1,     4,     3,    -1,     1,     3,     6,     6,     2,    -8,    -8,    -8,    -3,    -6,    -4,     1,    -1,     1,    -1,    -5,    -5,    -9,    -3,    -6,     0,     6,     3,    -3,    -5,     1,     1,     3,     2,     0,     7,     5,     6,    -2,    -3,     3,     1,    -2,    -4,    -7,     0,    -1,    -6,    -4,    -6,    -7,    -9,    -7,     0,     2,     1,    -3,     0,    -5,    -1,    -3,    -2,    -1,     0,     2,    -3,    -5,    -6,    -2,     1,     3,    -5,    -3,    -4,    -5,    -2,    -2,    -2,    -6,     2,    -1,     3,     6,     4,    -2,    -2,    -1,    -3,    -1,    -1,    -2,     1,    -3,    -8,    -7,    -8,    -4,     2,    -1,    -6,    -2,    -1,    -5,     2,     7,     7,     3,     3,     0,     3,     7,    -1,    -1,    -2,    -3,    -3,    -4,     2,     5,     5,    -2,    -1,    -2,    -7,   -10,    -6,    -8,   -13,    -5,     1,    -6,    -5,     4,    15,     8,     9,     6,     1,     1,    -2,    -3,     2,    -3,    -3,     2,    11,     9,     1,    -3,    -3,    -2,    -5,    -3,    -4,     2,    -4,    -2,     1,   -12,    -1,     0,     8,     9,     8,     1,    -4,    -1,    -1,     1,    -1,     4,     5,     3,    12,     8,     1,    -6,    -3,    -1,     3,     3,     1,     7,    -2,    -3,     1,    -3,     2,    -3,     6,     5,     7,    -2,    -1,    -2,    -2,    -1,    -1,     2,    13,     9,     5,     1,     2,    -2,     2,    -1,     2,     2,    -3,    -4,    -5,    -3,     0,    -3,    -2,    -3,     5,     7,    -1,     0,    -3,    -3,    -2,     1,     0,     9,    12,    12,     6,     1,     2,    -3,     0,     2,     3,     1,     0,    -2,    -4,    -2,     0,    -4,    -5,    -4,     1,     1,     4,     1,     1,     2,    -1,     1,     4,    11,    13,     9,     9,     3,     3,     4,     3,     0,    -3,    -5,    -4,    -4,     0,     0,     1,     1,    -9,    -3,    -2,    -2,     3,    -1,    -5,    -2,    -2,     0,     4,    12,    12,     7,     7,     2,     7,     4,     6,     2,    -4,    -8,    -8,    -3,    -1,    -2,     1,    -2,    -8,    -7,    -2,    -4,     5,     2,     4,    -3,     4,     3,     6,     6,    10,     7,     1,     4,     7,     6,     9,     0,    -2,    -4,   -11,    -8,    -2,    -3,    -1,     0,    -7,    -1,    -3,    -7,     5,     7,    -1,     2,     1,     8,     6,     4,     9,     3,     2,     4,     6,     4,     6,     0,    -2,    -4,   -10,    -4,    -6,    -2,     3,    -1,    -8,    -3,    -8,    -8,     6,     7,     7,     5,     3,     1,    -1,     2,     1,     2,     1,    10,     4,     7,     4,    -3,    -1,    -6,   -12,    -6,    -6,    -6,     0,     0,   -10,    -3,    -9,    -8,     4,     7,     5,     6,     3,     2,    -2,     1,    -4,     1,     8,     6,     3,     1,     0,     0,     3,    -1,    -3,    -2,    -3,    -2,     0,    -1,   -10,    -4,    -9,    -6,    -4,     2,     6,     1,    -3,     0,     2,    -2,    -5,    -1,     4,     2,     0,     0,    -1,    -3,    -3,     0,    -1,     3,    -3,     1,     0,     1,    -9,    -4,    -7,    -1,    -3,     1,    -5,    -2,    -4,     1,     2,    -4,    -4,     4,     0,     0,    -5,    -4,    -2,    -2,    -4,    -2,     2,     0,    -8,     0,    -1,     0,    -6,     5,    -5,    -7,    -2,    -4,    -4,    -2,    -1,     1,     1,    -7,    -2,     1,    -6,    -6,    -7,    -4,    -3,    -7,    -5,    -4,     2,    -6,    -2,     0,     0,     1,    -4,     1,    -3,    -5,    -1,    -6,    -7,    -6,    -6,    -1,     2,    -1,     1,    -4,    -7,    -6,    -5,    -4,     5,    -5,    -5,    -7,     1,    -2,    -4,    -1,    -1,     1,    -5,    -7,    -2,     2,    -6,    -6,    -3,    -3,    -2,    -2,     1,     0,    -3,    -9,    -7,    -4,    -6,    -5,    -3,    -3,     0,    -3,     0,    -1,    -1,    -1,     0,     1,     4,    -3,    -1,    -2,    -7,   -10,    -6,     0,    -4,    -3,     0,    -2,    -2,    -8,     1,    -2,    -2,    -5,    -3,    -3,     0,     4,    -2,     0,    -2,     0,    -1,    -1,     0,     7,    -3,    -7,    -5,    -6,    -5,    -4,    -4,     0,     1,     0,     0,    -2,     6,     4,     3,    -7,     0,     1,    -1,     1,     1,     1,     1,    -1,     1,    -1,    -1,    -1,    -1,    -2,     3,     4,     2,     3,     2,     1,     0,     5,     2,    -2,    -1,    -4,     0,     0,    -2,    -4,    -2,    -4,     0,     0,     0,    -1),
		    30 => (    1,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     0,     0,    -1,     1,     0,    -2,     0,     0,     0,    -1,     0,    -1,     0,    -1,     1,     0,     1,    -1,     1,    -1,    -1,     0,     0,     1,     0,    -1,    -5,    -5,    -8,    -5,     4,     2,     1,    -3,     5,     7,     5,    -3,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     7,     6,     0,    -1,    -1,    -5,    -6,    -9,   -12,    -7,   -10,    -9,   -15,   -13,   -14,    -9,    -8,    -7,    -6,    -9,    -5,    -3,    -3,     0,    -1,     1,     1,     0,     4,    -2,    -5,    -4,    -7,    -7,    -2,    -8,     1,     4,     6,    -3,   -10,    -4,    -2,    -9,   -13,    -3,    -5,    -5,    -5,    -7,    -1,    -4,     0,     1,     0,    -4,    -9,    -2,   -11,     1,     0,    -1,     1,     2,    -1,     2,     1,    -4,    -4,    -9,     0,     0,     4,     0,     0,    -3,    -6,   -10,   -12,    -5,    -1,    -1,    -1,    -2,    -6,    -1,    -2,     4,     2,     0,    -3,     2,    -2,    -7,    -7,    -2,    -5,    -6,    -1,     3,     3,    -4,    -4,     1,    -7,    -1,   -15,    -9,    -1,    -1,     0,    -2,     0,    -2,     0,     1,     4,     2,   -11,     0,    -4,    -8,     1,    -2,    -2,    -2,     0,     0,     1,    -3,     0,     2,     0,     3,   -13,    -4,    -1,     1,    -3,     0,    -4,    -1,    -1,     0,     0,    -5,     0,    -1,     6,    -2,     5,    -1,    -4,     2,     0,     3,     5,     2,     6,     3,     8,     2,     0,    -8,     0,    11,    -8,     5,     1,    -3,    -9,    -7,    -3,    -2,     0,     6,     0,     2,    -1,     1,     7,     6,     8,     2,     6,     7,     6,     6,     0,     1,    -7,   -11,    -4,    -1,    -1,     9,    -6,    -6,    -4,    -5,    -6,     0,     3,     2,     0,     0,    -1,     4,     3,     4,     3,    -3,     1,     8,     4,    -1,     0,     2,    -9,    -5,    -2,    -2,    -1,     8,     4,    -8,    -4,     3,     0,    -1,    -1,     1,    -2,    -3,    -2,     0,     6,     3,     6,     1,     0,     3,     3,     1,    -5,    -4,   -10,   -12,    -1,    -1,     8,    -6,    -2,   -14,     0,     2,     2,     2,    -4,    -3,    -6,    -5,     1,    -3,    -5,    -3,    -2,    -3,    -4,     0,     7,     2,    -8,   -10,   -10,    -8,    -1,     0,     2,    -6,    -2,    -3,     2,     5,     3,     0,     2,    -1,    -8,    -3,    -2,    -8,    -4,    -1,    -3,    -4,    -2,     0,     5,     6,     0,    -5,    -3,    -4,    -3,    -1,     2,     0,     4,     6,     2,     9,     5,     0,     4,     0,    -5,    -2,    -7,    -3,    -7,    -2,     3,     1,     2,    -7,     3,     0,     0,    -6,    -3,    -5,    -5,     1,     0,     0,    -1,    11,    12,    12,     6,     4,     6,     6,     2,     0,    -5,    -6,    -1,    -6,    -1,     1,     3,    -2,    -8,     0,    -4,     3,    -8,   -11,     0,     0,     0,    -5,    -4,     8,    14,     4,     8,     9,    13,     8,    -3,     6,    -4,    -5,    -2,    -4,     0,    -1,    -3,    -1,    -6,     1,     2,     0,    -6,   -12,    -6,    -1,     0,    -3,    -9,     8,     9,     5,     6,    11,    12,     5,     9,     7,    -4,     1,     3,    -3,    -2,     0,    -4,    -3,    -7,    -8,     4,    -9,   -13,   -17,     9,     1,    -1,    -3,   -12,     3,     3,    -2,     5,     3,     5,     7,     8,     0,    -4,    -2,    -1,    -1,     1,     1,     0,     0,    -8,     2,    -3,    -9,   -10,    -9,    12,    -1,    -1,    -2,   -13,     0,    -2,    -2,     0,     6,     3,     4,     1,     3,    -1,    -1,     0,    -2,    -4,    -4,    -3,    -3,    -3,     0,    -3,    -4,    -8,    -9,    -3,     0,     3,    -3,    -9,    -4,    -1,    -2,    -1,    -2,    -7,    -4,    -1,     5,     1,    -1,     0,    -3,    -5,    -1,     0,    -4,     0,     1,    -4,    -4,   -13,    -7,    -3,     0,     4,    -3,   -11,    -3,    -1,    -2,    -4,    -6,    -8,    -3,     2,    -1,     2,     5,     2,    -1,    -4,     0,    -4,    -3,    -2,    -2,    -3,    -5,   -12,     0,    -1,    -1,     1,   -10,    -7,    -7,    -2,     4,     1,    -3,    -3,    -2,    -2,     3,     7,     5,     6,     6,     2,    -3,    -8,    -7,    -3,     1,    -3,    -4,    -3,     8,     3,     0,     1,   -13,    -4,   -12,    -4,     0,     2,     8,    -1,     3,     3,    10,     4,     8,     7,     1,    -1,    -4,    -4,     0,     3,     4,     5,    -5,    -3,     5,     2,     0,    -1,    -3,   -13,   -11,    -3,     3,    -2,     0,    -3,     2,     2,     3,     3,     5,     1,     4,    -4,    -3,    -3,    -3,     3,    -2,    -4,    -5,    -4,   -10,     0,    -1,     0,    -1,    -3,    -2,     4,    -3,    -6,    -7,   -12,   -11,    -7,     3,     9,     8,     7,     7,    -1,    -3,   -12,    -8,    -4,    -6,    -7,    -4,     0,    -1,     1,     1,     1,     0,    -4,   -20,   -16,    -4,    -1,    -2,   -13,   -10,    -7,    -1,    -3,    -4,    -6,    -2,    -1,    -8,   -13,   -10,    -9,    -5,    -2,     0,     0,     1,     0,     0,     0,     1,    -1,   -10,    -9,   -13,    -4,    -6,   -10,   -10,    -5,    -6,    -6,   -11,    -9,    -6,   -14,   -14,    -7,    -9,   -10,    -4,    -6,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -4,    -2,     1,     1,     1,    -3,     0,     0,    -2,    -2,    -3,    -3,    -1,    -5,    -5,    -4,     0,     1,    -1,     1),
		    31 => (    1,    -1,     0,    -1,     0,    -1,     0,     1,    -1,    -1,     0,    -1,     1,     1,    -1,     1,    -1,    -1,     1,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,     0,     1,     1,     1,    -1,    -1,    -1,    -1,     0,    -2,    -2,    -1,    -5,     2,     3,     0,    -3,    -1,     1,    -1,     1,     0,     0,     1,     1,     1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     1,    -4,    -6,    -4,    -4,    -8,     3,    -2,    -1,     3,     1,     2,     7,     6,   -11,    -9,    -5,    -2,    -2,     1,    -1,     0,     0,     5,     4,     0,    -5,    -7,     4,     6,     6,    -1,    -7,    -3,    -4,     0,     5,     1,     0,     0,     6,     5,    -3,    -1,    -3,    -5,    -1,    -1,     0,    -1,    -1,     6,     5,     4,     6,     0,     0,     4,     1,     4,    -1,     0,     3,    -1,    -1,     0,     6,     9,     6,    -1,    -1,     1,    -1,    -3,    -6,    -8,    -6,     1,     1,     3,     2,     7,     8,     6,     6,    -3,    -6,    -2,    -3,     0,    -1,    -4,     0,    -2,    -2,     0,     6,     3,    -2,    -2,     4,    -2,    -9,    -6,    -6,     0,    -1,    -5,     2,     7,     6,     7,     5,    -3,    -3,     0,    -2,    -5,    -3,    -3,    -4,     1,     0,     1,     3,     2,    -4,    -4,     0,    -1,    -4,    -9,    -1,     0,    -3,    -8,    -3,   -12,     1,     6,     7,    -5,    -3,    -4,    -2,     0,     2,     2,     1,     1,    -6,    -1,     2,     3,    -2,     0,     4,    -1,    -7,   -16,    -9,     0,    -8,    -9,   -12,   -11,    -5,     2,     0,    -6,    -4,    -1,    -1,     6,     5,     7,    -1,    -1,    -3,     2,     1,    -5,    -3,     3,     1,    -1,    -6,   -22,    -4,     1,    -2,    -7,   -13,   -10,    -5,    -6,    -3,    -6,    -4,    -1,     2,     7,     8,     5,    -2,     0,    -3,     0,     1,    -4,    -7,     0,    -3,    -6,    -6,   -10,    -6,     0,    -2,    -7,    -4,   -10,    -7,    -7,    -4,    -5,    -9,    -5,    -2,     9,     8,     5,    -1,    -2,     2,    -3,    -4,    -5,    -5,    -7,    -7,    -6,    -4,    -3,    -1,    -1,     2,    -1,    -6,    -6,    -8,   -10,    -9,    -9,    -6,    -7,    -6,     0,     7,     2,     4,    -3,    -2,    -2,    -5,     1,    -4,    -2,    -8,    -9,    -5,    -5,     7,     0,    -1,   -11,    -3,    -1,    -7,    -6,   -13,    -9,    -7,    -4,    -4,     1,     7,    -1,     0,     5,     1,    -2,    -2,     2,    -6,    -6,    -3,    -6,    -2,     1,     6,     1,     0,    -9,     3,    -3,    -8,    -4,    -7,    -6,    -5,    -4,    -6,     0,    -1,     3,     3,     8,     5,    -1,    -2,    -2,   -11,    -9,    -9,    -8,     1,     1,    -1,    -1,     0,     2,     1,    -4,    -5,    -6,    -4,    -6,    -3,    -6,    -6,     2,    -1,     1,     2,     2,     1,    -3,    -7,    -2,    -8,    -6,    -5,    -6,    -6,    -2,    -1,     0,     0,     1,    -4,    -8,    -7,    -7,    -8,    -6,    -1,    -1,    -1,     0,     3,     2,     1,     3,     3,     2,    -3,    -7,   -13,   -11,    -8,   -21,   -10,    -6,    -4,    -1,     0,     2,    -9,    -8,    -1,    -3,    -6,    -3,     2,    -2,    -3,    -2,     1,     1,    -1,     3,     0,    -1,    -2,    -5,    -9,    -5,    -4,     2,    -7,    -4,    -5,     1,     0,    -3,   -10,    -4,    -3,    -5,   -10,     2,     0,     3,     4,    -3,    -3,     6,     5,     4,     2,    -1,     0,    -2,     3,     3,    -2,     2,    -4,    -6,    -5,    -1,     1,     1,   -11,    -7,    -7,   -15,   -10,     0,     4,     5,    -2,    -6,    -3,     2,     7,     6,    -2,     2,    -7,    -4,    -2,    -2,     2,     2,    -1,    -5,     0,    -1,     0,    -2,   -11,   -13,     1,     0,    -1,     4,     5,     5,    -2,    -3,     2,     3,     3,     3,    -3,    -4,    -9,    -6,     0,     5,     5,     6,     3,    -6,    -1,    -1,     1,    -4,   -11,    -2,     6,     8,    10,     2,     7,     6,     1,     3,     4,     3,     2,     2,    -4,     2,    -2,     2,     3,     6,     5,     6,     1,    -2,     0,     4,     2,    -1,    -1,    -2,     4,     5,     7,     9,     9,     4,     0,     4,     8,     0,    -4,     1,    -3,     1,    -1,     3,     4,     5,     1,     1,     3,    -4,     1,     2,     2,    -3,    -1,    -1,     6,     7,     7,     6,     9,     4,     4,     4,     8,    -8,    -5,    -1,    -2,     1,     3,     6,     5,    -5,    -2,     4,     0,     1,     0,     0,     1,    -2,    -2,    -3,     2,     2,     0,     2,     9,     5,     5,     6,     0,    -7,    -4,    -6,     2,    -2,    -2,     3,     0,    -2,    -6,    -6,    -5,     8,    -1,     0,    -1,     1,    -1,    -5,     1,    -3,     1,    -2,     3,     3,    -6,    -2,    -1,    -7,    -7,    -7,     1,    -1,    -7,    -2,     3,    -1,    -8,    -8,     1,     1,     1,    -1,     0,     0,    -2,    -6,    -9,    -5,   -13,     1,    -5,    -1,    -5,     4,     0,    -6,    -8,    -9,   -13,   -15,   -11,   -20,    -7,    -5,    -4,    -2,    -2,    -2,     0,     0,    -1,     0,    -2,    -6,   -13,   -19,   -21,   -14,   -13,     2,     0,    -8,    -8,    -8,    -8,    -5,   -11,    -5,    -2,    -4,    -4,    -1,    -1,     0,     0,    -1,     1,    -1,     0,     0,     1,    -1,    -2,     0,     1,     1,    -1,    -8,    -6,     1,    -2,    -6,    -2,    -2,    -1,     0,     0,     1,    -1,    -1,     1,     0,    -1,     1,     1),
		    32 => (    0,     1,     0,    -1,    -1,     0,     0,     1,     0,    -1,     0,    -1,    -3,    -2,     1,     0,     0,    -1,     0,     0,    -1,     1,     1,     0,     0,     1,     1,     0,     0,    -1,     0,     1,     0,     0,     1,     0,    -5,    -3,    -3,    -1,    -2,    -2,    -8,     0,     1,    -2,    -1,    -6,    -3,    -2,    -3,     0,     1,    -1,     0,     0,     1,    -1,     0,    -1,    -2,    -1,    -1,    -4,    -2,     1,     2,    -2,     1,    -2,    -1,    -3,    -4,    -5,     2,     0,    -5,    -2,    -2,     0,     0,     2,     1,     0,    -1,    -1,    -1,    -2,    -4,     3,     2,     2,    -4,    -4,    -7,    -4,    -7,    -9,    -5,    -3,    -9,   -11,    -8,    -2,    -7,    -8,    -3,    -1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,     5,     6,     8,     6,     6,     4,     0,     2,     3,    -3,    -4,    -2,    -2,    -7,    -2,    -1,    -6,    -5,    -8,    -4,    -3,    -2,    -4,     0,    -1,    -1,     2,     1,     2,     0,     2,     1,     3,     5,     3,     3,    -1,    -4,    -6,    -8,    -2,    -1,    -5,    -4,    -3,    -2,    -5,    -4,    -1,     0,    -3,    -2,     1,     0,    -3,     5,     4,     5,     7,     0,    -2,     0,     0,     1,    -3,    -2,    -3,    -3,    -1,     0,    -1,     0,    -4,    -2,    -1,    -5,    -2,    -4,    -2,     0,     1,     0,     1,     7,     7,     3,     7,     3,     7,    -1,    -3,     0,     3,    -1,    -5,    -2,    -1,    -5,     0,    -2,    -2,    -2,    -4,   -11,    -7,    -3,    -4,    -2,    -3,     2,     0,     3,     4,     2,     6,     5,     4,     4,     1,    -1,     3,    -2,     3,    -2,    -8,    -3,    -5,    -2,    -2,    -7,     0,    -4,    -8,    -4,    -6,    -2,     1,    -1,    -1,    -2,     1,     4,     1,     1,    -1,    -2,    -8,    -5,    -3,    -4,     1,     0,    -2,    -5,    -2,    -1,     0,    -2,     2,    -2,    -7,    -3,     2,    -1,     0,    -1,     1,    -7,    -4,     0,     3,     0,    -2,    -7,    -6,   -13,   -13,    -6,    -1,     0,    -2,    -3,    -2,    -2,     2,    -4,    -5,     0,    -3,    -3,    -3,    -1,     1,    -1,    -3,    -4,    -5,    -4,    -1,    -2,    -3,    -7,    -2,    -4,   -12,    -6,    -3,    -2,     0,    -4,    -3,    -1,    -2,    -4,     0,    -2,     0,     1,    -8,    -2,     1,     0,    -1,     0,    -7,   -12,    -9,    -8,    -7,    -7,    -4,    -2,    -4,    -6,    -3,    -6,    -3,    -1,    -4,     0,    -3,    -3,     4,     1,     7,     2,    -1,    -1,    -1,     0,     0,    -2,    -2,   -11,   -14,   -12,    -8,    -8,    -5,     1,     0,    -1,    -3,    -7,    -4,    -5,    -3,     0,     3,    -2,     5,     7,    10,     6,     1,    -2,     1,    -2,    -2,    -1,    -5,    -9,   -14,    -9,    -7,    -4,     4,     2,    -3,    -6,    -1,    -4,    -5,    -8,    -2,     6,     1,     2,     5,     3,     2,     1,     3,     5,     1,    -3,     4,     3,    -4,    -9,    -8,    -1,     0,     2,     4,    -1,     2,     4,     4,     0,    -2,     1,     1,    10,     8,     4,     1,     5,     6,     6,     4,     7,    -1,    -2,     5,     1,    -3,    -9,    -1,     1,     0,     0,     2,     1,     1,     1,     0,    -2,    -7,     1,     6,     8,     1,     5,     6,     6,     2,    10,     3,     4,     1,    -1,     7,    -2,    -5,    -2,     2,     5,     3,     6,    -1,     0,    -4,    -4,     2,    -1,    -8,     5,     8,    -2,    -1,     4,    -1,    -1,    -7,     6,    -1,     4,     0,     1,     1,     5,    -7,     1,     3,     3,     3,    -1,    -4,    -3,     1,    -4,     0,    -3,     2,     6,     4,    -4,    -6,    -2,    -3,    -3,     3,     8,     1,    11,    -1,    -5,    -3,    -2,    -7,     0,     2,     5,     2,    -3,    -4,    -1,    -2,     0,    -2,     0,     4,     5,     1,    -4,    -6,    -8,     1,    -5,    -7,     0,     7,     8,    -1,    -5,     0,    -1,    -5,     0,     3,     3,     2,    -4,    -5,     0,     1,     3,    -3,     0,     1,    -1,    -1,    -4,    -6,    -6,    -5,    -6,    -8,    -1,     1,     1,     0,     1,     2,     1,    -8,    -5,    -1,    -5,     3,    -1,    -2,     2,     0,     2,     0,     3,     5,     0,     1,    -3,     0,     1,    -3,     1,    -5,    -1,     2,    -1,     0,     1,    -1,     3,    -6,    -9,    -5,    -5,    -4,    -4,    -2,     5,     1,     6,     5,     0,     0,     2,     0,    -3,     1,     0,    -6,     1,     0,    -1,    -3,     0,     0,     0,    -1,     4,    -6,    -8,    -6,    -4,    -4,     0,     3,     2,     7,     4,     1,     1,     2,     3,    -3,    -2,    -3,    -1,     1,     3,     1,     2,    -4,     0,     0,     1,    -6,    -5,   -10,    -6,    -9,    -3,    -6,    -8,    -7,    -6,    -5,    -6,    -2,    -3,    -7,    -2,     1,     2,     1,    -3,     0,     2,     4,    -1,     1,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -4,    -9,   -12,    -9,    -9,   -15,    -1,    -1,    -4,     0,    -3,     3,     4,     3,    -4,    -1,     1,     1,     1,     0,     0,    -1,     1,    -1,     0,    -4,    -4,    -4,    -3,    -7,    -1,    -2,    -4,    -4,    -5,    -3,    -7,    -8,    -7,    -4,    -4,    -3,    -4,     0,     0,     0,    -1,     0,    -1,     0,     1,    -1,    -1,     0,     1,     0,    -1,     0,    -3,    -2,    -3,    -5,    -4,     1,     0,    -2,    -1,    -1,    -2,    -4,    -3,     0,     1,     0,    -1,     1),
		    33 => (   -1,     0,     0,     1,     1,     1,     0,     1,     1,    -1,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     1,     1,     1,    -1,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     1,     0,     0,     0,     1,    -1,    -1,     1,     0,    -1,     0,     0,     0,     0,     1,    -1,     0,    -3,    -4,    -2,    -2,    -5,    -4,    -7,     0,    -2,    -1,    -3,    -2,    -4,    -2,    -2,    -3,     0,     1,    -1,    -1,     0,     1,     0,    -1,     0,     0,     1,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -3,    -2,    -1,    -3,    -1,    -1,    -1,    -3,    -4,    -3,     0,     0,    -1,     0,     0,     4,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -2,    -2,    -1,    -1,     0,    -1,    -3,    -2,    -3,    -2,     0,     0,    -8,    -4,    -2,     0,     0,     0,     0,     2,     4,    -1,     1,    -1,    -3,    -4,    -3,    -4,    -5,    -2,    -4,    -1,     0,     3,     4,     3,     0,    -2,    -3,    -2,    -2,    -7,    -2,     0,     0,    -1,     3,    -1,     3,     3,     1,     1,     0,     1,     2,     1,     2,    -1,    -2,    -2,    -4,    -5,     1,     1,    -2,    -5,    -4,    -3,     0,     0,    -5,    -1,     0,     1,     5,     0,    -1,     3,     0,     3,     3,     3,     1,     3,     0,    -3,    -3,    -5,    -4,    -2,    -4,    -9,    -5,    -3,    -4,    -3,    -3,    -1,    -7,    -2,    -1,     2,     5,     4,     3,    -1,     3,     4,     3,    -2,     1,    -2,    -4,    -1,     1,     2,     0,     2,     0,     0,    -4,    -2,    -1,    -1,    -1,    -4,    -6,     0,     1,    -5,    11,     3,     3,     0,     6,     2,     0,     3,     3,    -5,    -3,     1,     4,    -1,    -7,     1,     3,    -1,     0,     2,    -3,     0,    -6,    -7,    -3,     0,     1,    -4,    10,     3,    -1,    -3,     3,     0,    -3,    -6,    -4,    -4,     0,     1,     5,    -5,    -6,    -1,     1,    -1,     1,     2,    -1,    -1,    -5,    -3,    -1,    -1,     0,    -1,    -4,    -3,    -2,    -4,    -6,    -5,    -6,    -7,    -3,     0,     2,    -3,    -5,    -5,    -1,     0,     1,     0,     1,     2,     2,    -1,    -3,    -6,    -2,     0,     1,     0,    -5,    -2,    -2,    -6,    -7,     0,    -2,    -2,    -1,     0,    -3,    -9,    -4,     0,     0,     3,     3,    -1,     0,     0,     0,    -2,    -2,     1,     0,    -1,     1,     1,    -3,    -2,    -1,    -3,    -4,     0,     1,     1,    -3,     0,    -3,     2,    -1,    -1,    -2,     3,    -2,    -2,    -4,     0,     1,    -2,    -3,    -3,    -3,    -2,     0,     3,    -1,    -2,     0,    -1,    -2,    -5,    -2,    -3,     0,    -1,    -3,     1,     3,     2,     1,    -4,    -6,    -3,    -5,    -2,    -2,    -1,    -2,    -7,    -3,    -2,    -1,     2,    -1,    -3,     2,    -3,    -3,    -1,     0,    -2,     0,     0,     1,     2,     2,    -2,     0,     0,    -3,    -5,    -3,    -3,     2,     0,    -2,     0,    -1,     0,    -1,     0,    -2,    -2,     0,    -3,    -1,    -3,    -1,     5,     1,    -1,    -1,     1,     0,    -2,     0,    -5,    -1,     0,    -1,     0,     2,     0,    -1,     1,    -5,    -3,    -1,     2,    -1,     4,     1,    -1,     0,    -2,     0,     4,    -1,     2,     2,    -1,    -2,     0,    -1,    -6,    -5,    -3,    -2,     0,     2,     0,    -3,    -1,    -1,    -2,    -2,     0,     0,     3,     3,     2,     0,    -4,     0,     3,     6,    -1,     1,     5,    -1,    -2,    -2,    -5,    -5,    -3,    -1,     3,     4,     1,    -3,    -2,    -1,    -3,    -1,     0,     1,     1,     4,     3,     1,    -2,    -1,     0,     2,    -2,     2,     1,    -3,    -2,    -4,    -3,    -3,    -3,     2,     1,     5,     4,    -3,    -1,    -2,    -2,     0,     0,    -1,     1,     1,     2,     2,    -2,    -3,     1,     0,    -7,    -1,     3,     0,    -3,    -1,    -2,    -3,     1,    -1,     2,     5,     4,    -4,    -4,     0,    -1,     0,     0,     1,     2,     3,     1,    -1,    -4,    -6,    -1,    -3,    -6,    -6,    -4,    -6,    -1,     2,    -3,    -1,     0,     0,     0,     0,     4,    -3,    -3,     0,     1,    -2,     0,     0,     2,     5,     1,     0,    -3,    -6,    -3,    -2,    -7,    -9,    -5,    -9,    -6,    -2,    -2,     5,     6,     2,    -2,     0,     4,    -1,    -3,    -1,     1,     0,     1,     3,    -1,    -1,    -2,    -1,    -1,    -4,    -7,    -2,    -2,    -5,    -4,    -6,    -1,     4,     2,     3,    -2,     0,     1,     2,     0,    -2,    -3,     1,    -1,     0,     0,    -2,     0,    -2,    -2,    -1,     2,    -4,    -5,    -6,    -1,    -7,    -2,     3,     8,     5,     0,    -2,    -1,     0,    -1,    -3,     2,    -5,    -3,    -1,    -1,     0,     0,     2,    -2,    -6,    -6,    -2,     1,     3,     0,    -2,    -2,     1,     8,    11,     2,     3,    -3,     0,     0,     3,     0,    -5,   -12,    -1,     0,     0,     0,     0,     1,    -1,    -4,    -4,    -4,    -7,    -5,    -5,    -7,    -4,    -3,     4,     8,     5,    -1,    -3,    -2,    -2,    -3,    -4,    -3,    -6,     1,     1,     0,     0,     1,     0,     1,     0,     1,     0,     0,    -1,     1,     1,    -4,    -4,    -2,    -2,    -2,    -2,    -4,     0,     0,    -2,    -1,    -2,    -2,     0,     0,     0,     0,     1,     0),
		    34 => (   -1,    -1,    -1,     0,     0,     0,    -1,     1,     0,     1,    -1,    -1,     0,    -1,     0,     1,     0,     1,     0,     0,    -1,    -1,     0,     0,     1,    -1,    -1,     1,    -1,    -1,     1,     1,     1,     0,    -1,    -3,    -2,     1,    -1,     0,     1,    -5,    -4,    -1,    -1,    -2,     0,     1,     0,    -1,    -2,    -1,     0,    -1,    -1,     0,     1,    -1,    -1,    -1,    -3,     0,    -2,    -4,    -2,    -1,    -2,    -2,    -1,    -3,    -4,    -2,    -1,    -3,    -1,     0,    -4,    -1,    -1,    -1,     1,     0,     0,     1,     1,    -1,     0,    -1,    -2,    -1,    -6,    -3,    -5,    -2,    -1,    -2,    -2,    -4,    -7,    -7,    -4,     2,     0,    -3,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     1,     0,     0,    -2,    -2,    -1,    -3,    -2,    -1,    -2,    -2,    -2,    -3,    -6,    -8,    -4,    -2,    -3,    -7,    -5,    -1,    -4,    -5,    -1,     1,    -1,    -1,    -1,     1,     1,     1,    -1,    -2,     0,    -2,    -1,    -3,    -4,    -1,    -5,    -8,    -5,     0,     3,    -2,   -10,    -9,     0,    -3,    -1,    -2,     4,     4,     0,    -4,    -1,    -1,     0,     1,    -3,    -2,     4,    -3,    -1,    -3,    -3,    -5,    -3,    -1,     0,     7,     0,   -15,   -18,    -6,     1,     7,     0,     4,    -4,     2,    -2,     4,    -6,    -1,    -7,     0,    -1,    -1,     6,    -1,    -1,     1,    -3,    -8,    -5,     3,     3,     3,   -12,   -17,   -13,    -2,     3,     2,    -1,     4,     3,     2,     2,     0,    -3,    -2,    -6,     2,    -1,    -1,     1,     1,     3,     0,    -2,    -8,     1,     4,     5,    -6,    -7,   -14,    -4,     1,     0,     2,    -1,     4,     1,     3,    -1,    -2,    -5,     1,    -5,     2,    -1,     1,    -2,    -4,    -2,    -4,    -6,    -5,     6,     1,     0,    -4,   -12,    -9,    -1,     2,     3,     2,     0,     1,     1,     1,    -3,     0,    -3,    -1,    -1,    -4,     0,     0,    -6,    -5,    -1,    -5,    -6,    -1,     6,     0,    -4,    -8,    -4,    -3,    -2,    -1,     0,    -1,    -6,    -9,     1,    -6,     0,    -2,    -2,    -1,    -1,    -4,    -2,    -4,    -4,    -3,    -5,    -1,    -2,     2,     3,     0,    -3,     0,     4,    -2,     0,     0,     5,    -2,    -3,    -5,    -6,    -4,    -2,    -4,    -6,     1,     0,    -7,    -5,    -7,    -4,    -5,    -3,    -4,     0,     3,    -2,     0,     0,     2,    -2,     0,    -2,    -2,     1,    -1,     2,    -3,    -5,    -4,    -3,   -10,    -6,    -1,    -1,    -5,    -5,    -8,    -4,     0,    -2,     0,     0,     7,     2,    -2,     2,     3,     3,     4,    -1,    -4,     3,     3,     1,    -5,    -6,    -6,    -8,    -9,    -1,    -1,    -1,    -3,    -7,    -8,    -3,    -3,    -1,    -3,     1,     3,    -1,    -2,     1,    -1,     4,     4,    -4,     0,     3,     6,     2,    -5,    -2,    -4,    -4,    -4,    -1,     0,     0,    -2,    -1,     1,    -3,    -5,     1,    -1,     1,    -1,    -2,    -1,    -1,     0,     6,    -3,     0,    -3,     5,    -4,     1,     0,     2,    -4,    -3,    -1,     2,    -1,     1,    -2,     0,     0,     2,    -3,     0,     3,     3,    -3,    -3,    -2,     2,     0,    -1,    -3,    -5,    -9,    -3,    -5,    -4,    -3,     1,     1,     0,    -2,    -1,     1,     0,    -4,    -1,    -3,    -3,     1,    -3,     3,    -1,    -5,    -1,    -3,    -4,    -3,    -1,     3,    -6,    -7,    -6,    -4,    -1,    -2,     2,    -1,     0,     0,    -2,    -1,     1,    -4,     2,     3,     0,    -1,     0,    -7,    -7,    -5,     0,    -3,    -2,    -1,    -1,     0,    -6,     0,    -1,     1,     0,    -2,     0,    -1,    -1,     1,    -1,     1,    -5,    -5,     1,     5,    -2,    -6,    -6,    -7,    -4,    -7,     0,     0,    -2,    -1,    -1,     0,    -4,    -1,     2,     0,    -3,    -4,     0,    -1,     1,     0,    -2,     0,    -1,    -1,    -2,     1,    -4,    -9,    -6,    -9,    -3,    -2,     2,    -3,    -3,    -5,    -7,    -3,    -6,    -3,    -2,    -3,    -3,    -1,     2,     1,    -3,    -1,     1,     0,     1,    -3,    -4,     0,    -3,   -12,    -7,    -1,     0,     0,    -2,     0,    -2,    -4,    -5,    -9,    -5,     1,     1,    -3,    -4,     2,     2,     2,    -7,    -2,     0,    -1,     1,     1,    -3,    -4,     0,    -4,    -6,     1,     0,     2,     4,     1,    -2,    -6,    -2,    -4,    -3,     2,    -4,    -3,     0,     1,     0,     1,     0,     0,    -1,    -1,     1,    -3,    -2,    -2,    -5,    -3,    -4,     1,    -2,     1,     0,    -4,    -7,    -4,    -1,    -2,    -2,     5,     3,    -6,     0,     1,     4,     2,     1,     1,     0,     1,     1,     0,    -1,    -5,    -3,    -1,    -1,     1,     2,     4,     2,    -6,    -1,    -1,     2,     0,    -2,     6,     6,     4,     2,     3,     3,    -1,     6,     0,     1,     0,     0,    -3,     1,    -5,    -1,    -5,    -3,    -5,    -4,     1,     1,     2,     1,     1,    -3,    -5,     0,     5,     5,     2,     1,     5,     2,     2,    -1,    -1,     1,     0,     0,     0,    -1,    -4,    -1,    -3,    -4,    -4,    -5,     1,    -2,     2,    -2,    -6,    -3,    -1,    -3,    -6,    -3,    -3,    -9,    -9,     0,    -2,     0,     0,    -1,     1,    -1,     0,     1,     1,     0,    -2,    -1,     0,    -2,    -8,    -8,    -5,    -5,    -6,    -1,    -3,    -7,    -2,    -4,    -3,    -3,    -2,    -2,    -1,     1,     1,     0),
		    35 => (    1,     0,     1,     1,     0,     0,    -1,     0,     0,     1,    -1,     0,    -1,    -1,     1,     0,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,     1,     1,     0,    -1,     0,     1,     0,     1,     0,    -1,     0,    -1,    -1,     1,    -2,    -2,    -1,    -1,    -2,    -4,    -3,    -1,    -3,    -1,    -2,    -1,    -1,     0,     0,    -1,    -1,     1,    -1,    -1,    -2,    -2,     1,    -3,    -3,    -3,    -5,    -6,    -5,    -7,    -6,   -15,   -10,    -6,    -3,    -2,     2,     0,    -7,    -3,     1,    -3,    -2,     0,     0,     1,     1,    -1,     1,    -1,    -6,    -5,    -4,   -10,   -11,    -8,    -2,    -2,    -1,    -2,    -3,    -4,     3,     7,     3,    -4,    -2,    -3,    -4,    -4,    -1,     1,    -1,     0,     0,    -2,     2,    -4,    -2,    -6,     0,    -2,    -1,     3,    -2,    -7,    -2,     3,     4,    -1,    -3,     0,    -4,    -5,    -2,    -5,    -8,    -9,    -6,    -2,    -1,     0,     0,    -1,    -1,    -4,     0,    -4,    -9,    -6,    -3,    -4,    -1,    -6,    -6,    -3,    -6,    -6,   -10,   -11,    -2,     2,    -5,    -5,    -1,    -6,    -8,     2,     1,    -1,     0,     4,    -6,    -6,     3,    -3,    -5,    -2,    -5,     1,    -2,    -6,    -2,     0,    -3,    -5,    -4,    -2,    -1,    -1,    -1,     0,    -1,     0,    -7,    -1,     0,     1,    -2,     4,    -3,    -7,     3,    -7,    -3,    -1,    -1,     9,     2,    -3,     0,    -1,     2,    -5,    -6,   -10,   -10,    -3,    -1,     1,     1,    -3,    -2,     0,     5,    -1,     0,    -5,     1,    -2,    -2,    -4,    -1,     0,     1,     2,     3,    -2,    -2,     3,     3,     4,     3,     0,     4,     4,     4,     6,     7,     6,     4,    -4,     3,     0,     0,    -5,    -4,    -3,    -9,     2,     3,    -1,    -1,    -1,    -5,    -2,    -1,     3,     3,     7,    11,     8,     9,     6,     7,     6,     5,    11,     8,    -6,     1,     0,    -1,    -1,    -4,     0,    -2,     2,     2,    -2,     0,     1,     5,    -3,    -1,     1,     2,     1,     4,     9,     8,     8,    10,     7,     3,    11,     8,     4,     6,     1,    -1,    -1,    -1,     2,     0,    -2,    -6,    -2,    -4,     2,    -1,    -2,    -4,    -9,    -8,    -6,    -7,    -5,    -8,    -6,     2,     1,     4,     1,    10,     9,     1,     0,    -1,    -1,     1,    -2,    -3,    -4,    -1,     0,     3,     4,     6,     3,     0,    -4,    -6,   -10,    -8,   -17,   -28,   -18,   -12,   -12,    -7,    -6,     6,     9,    -3,     0,     0,    -1,     2,    -2,    -6,    -7,     3,     0,    -1,     7,     2,     4,     1,     1,     0,    -5,     0,    -6,   -12,   -15,   -10,   -13,   -14,    -5,    -2,     6,    -3,     2,     1,    -2,    -2,     3,    -1,     3,     2,     5,     5,     0,     0,    -1,    -1,    -1,     0,    -3,     2,     0,    -9,   -10,    -8,    -7,    -5,    -5,    -6,    -2,    -1,     1,     0,    -5,     5,     8,     4,     1,     6,     4,     5,    -1,     1,     2,    -1,    -4,    -5,    -8,    -2,     3,     0,    -4,    -4,    -7,    -3,    -5,     3,    -2,    -4,     0,     0,    -5,     1,     3,     9,    -1,     5,     0,     3,     0,    -3,    -3,    -1,    -7,    -3,    -4,    -2,     2,     0,     0,    -4,    -3,    -4,    -2,     3,    -5,    -5,     1,    -1,    -9,     1,     2,     2,     2,    -3,    -2,     2,     1,    -1,    -6,    -6,    -5,     0,    -3,     0,    -3,     0,    -3,    -5,    -2,    -2,    -8,    -9,    -9,    -9,    -2,    -1,    -5,    -9,    -4,    -3,     0,    -2,    -3,    -5,   -10,     4,     5,    -3,    -5,     1,    -4,     1,    -2,     0,     3,    -5,    -1,     5,     1,    -3,   -10,    -6,     0,     0,    -1,    -8,     4,     5,    -2,    -3,    -2,    -7,    -8,    -8,     0,     3,    -6,    -4,    -2,     2,     1,     4,     0,    -6,     2,     8,     8,     9,    -8,    -7,     0,     0,    -1,    -5,     4,     0,    -4,    -1,    -4,    -3,    -5,     0,     2,     3,   -10,    -3,     1,     0,     0,     3,     2,    -4,     2,     1,     9,    10,    -7,     0,     0,     1,    -2,    -4,    -2,     3,    -4,    -5,    -1,    -1,     1,     1,     2,     2,    -3,     5,    -2,    -1,    -1,    -1,     2,    -3,    -5,     0,     7,    12,     6,    -1,     0,    -1,    -4,    -1,    -2,     3,     3,    -4,    -6,    -1,     1,     2,     5,     1,     0,     4,     2,     4,     0,    -4,     1,    -1,    -4,     8,    14,    14,    13,     1,    -1,     0,     4,    -1,     0,     0,    -2,    -6,    -5,     3,     6,    -3,     0,    -4,     1,     2,    -2,    -1,     0,    -5,     0,    -4,    -1,    13,    14,    12,    16,    -1,     1,    -1,    -1,     0,    -6,    -9,    -6,    -4,    -2,    -3,     1,     2,     4,    -2,     4,    -2,    -1,    -2,    -3,    -3,     1,     4,     9,     5,     3,    -9,    -3,     1,     0,     1,     0,     0,    -9,   -10,    -6,    -8,    -6,    -3,    -5,     1,     9,     5,    -1,    -5,    -4,    -3,     2,     0,    -5,     4,     5,     7,     7,    -1,    -1,    -1,    -1,     0,    -1,     0,    -5,   -10,   -14,   -13,   -13,   -12,   -11,    -7,    -7,   -11,   -18,    -5,    -1,    -3,    -1,     1,     0,     2,     0,    -6,    -3,     1,     1,     0,     1,     1,     1,     1,     0,    -2,    -1,    -3,    -3,    -1,    -1,    -2,    -3,    -2,   -10,    -5,    -2,    -4,    -6,    -4,    -2,    -4,    -9,    -7,    -1,     1,    -1,     0),
		    36 => (    0,     1,     0,     1,     0,     0,     1,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,     1,    -1,     0,     1,     1,     1,     1,    -1,    -1,     0,    -1,     0,    -1,    -1,     1,    -1,     1,     1,     4,     4,     4,     3,     6,     1,     0,     3,    -4,     0,     1,     3,     5,     4,    11,     4,     4,     4,     1,     1,     0,     1,    -1,     0,     3,     2,     5,     5,     5,     7,     4,    -2,    -3,    -4,    -6,    -6,     1,     3,     5,     9,     5,     2,     2,    10,     9,     7,     4,     6,    -1,    -1,     0,     0,    -7,     1,    -3,     3,     7,     6,     0,    -3,    -3,   -10,   -13,     0,     6,     4,    -5,    -3,     2,    -3,    -3,     0,    -5,     2,    -7,    -4,    -6,    -1,     0,     1,   -10,    -1,     3,     8,     6,    -3,    -7,    -5,    -7,   -12,   -16,    -7,    -9,    -5,     0,    -3,    -2,    11,     7,     1,    -8,   -10,   -15,   -11,    -4,     3,     0,     0,    -5,    -6,     3,     6,     3,    -2,    -3,    -3,    -4,   -14,    -9,     0,     1,    -5,    -3,     0,     3,     3,     6,     4,    -3,     0,    -7,   -11,     1,     1,    -1,    -1,     5,     2,     2,     6,     6,    -1,    -2,    -7,    -8,    -5,    -3,    -5,    -4,     5,     4,     1,     0,    -1,     0,     0,     2,    -4,    -3,    -8,    -4,    -1,     0,    -1,    -1,    -2,    -2,     1,    -3,     0,    -5,    -9,   -15,   -11,    -4,    -4,     2,     4,    -4,    -6,    -2,   -10,     1,    -1,     4,    -5,   -12,   -12,    -2,    -5,     0,     0,    -5,    -4,    -2,     1,     4,    -5,    -7,   -14,   -14,    -2,     0,    -1,    -2,     2,     0,    -5,   -12,     0,    -4,    -5,    -5,   -13,   -11,    -5,    -5,    -6,     0,     0,    -5,    -3,     7,    -2,    -1,    -1,    -7,    -7,    -4,    -1,    -2,     1,     4,     2,    -5,    -9,   -12,   -15,   -19,   -17,   -16,   -15,   -12,    -6,    -7,    -2,     1,     1,    -4,    -2,    -4,    -5,    -6,    -6,   -12,    -3,     1,     0,     1,     2,     0,    -1,    -5,    -2,    -2,   -10,   -11,   -10,   -13,   -15,   -10,    -9,    -6,    -5,     0,     0,     1,    -7,    -3,    -1,    -2,    -3,     1,     0,     1,     2,     3,     3,    -1,    -7,    -6,    -3,    -5,    -2,    -3,    -5,     0,   -13,   -13,   -12,    -8,    -7,     1,    -1,    -2,    -5,    -5,    -2,    -1,    -5,    -1,     1,     5,     3,     2,     8,    -3,     1,    -5,     3,    -1,     0,    -2,    -4,     2,     2,    -5,   -12,   -12,    -6,    -1,     1,    -1,    -6,    -5,    -3,    -5,    -6,     1,     1,     2,     8,     2,     4,     0,     1,    -2,     2,     8,     0,     1,     0,     8,     7,    -7,   -14,    -7,     0,    -1,     1,    -1,    -8,    -5,     1,    -7,     0,    -2,     3,     5,     2,     0,    -3,    -2,     0,     0,   -10,     2,     4,     0,     7,     5,     0,     2,    -5,    -6,     0,     0,     1,     0,    -7,    -1,     2,    -4,     0,     3,     3,     3,    -6,    -2,    -2,     0,    -7,    -6,    -8,     2,     6,     3,     9,     3,     1,    -6,    -9,   -11,    -6,     0,     1,     0,    -2,    -2,     3,    -1,     5,    -1,     3,     0,     3,     6,     4,     3,     0,     2,     0,     0,    -1,     4,     8,     4,    -1,    -9,   -10,   -10,    -8,     0,     0,    -1,     0,     1,     2,     1,     1,     6,     0,     2,     3,    -3,     0,    -2,    -3,    -3,    -1,     0,     0,     3,     7,    -2,    -2,    -8,    -7,     0,    -8,     0,    -1,     1,     0,     6,    -2,    -4,    -2,    -1,     6,     4,    -3,    -2,    -3,    -1,     7,    -1,     3,     5,     3,     2,    -1,   -12,    -9,    -7,    -6,    -1,    -3,     0,    -3,    -3,     1,     4,    -4,    -2,     0,    -4,     1,     3,     5,     0,   -10,    -3,     3,    -1,    -1,     4,    -3,    -2,    -5,   -13,    -5,    -3,    -3,    -4,    -1,    -1,    -3,    -2,    -8,     5,     2,    -2,    -2,    -1,    -3,     1,     5,     5,    -3,    -1,    -2,    -7,    -5,    -7,    -2,     0,    -1,    -2,    -6,    -3,    -4,    -5,     1,     0,    -1,    -4,    -4,    -3,    -5,     0,    -1,    -1,     0,    -2,     5,    -3,    -1,    -3,    -6,    -2,    -4,    -2,    -4,    -2,     1,    -5,    -4,    -4,    -4,    -4,    -1,    -1,     0,    -1,    -3,    -5,    -7,    -8,    -4,    -5,    -3,     0,     1,     3,     4,     0,     1,    -2,    -5,    -3,    -5,    -8,    -7,    -2,    -5,   -10,    -4,     1,    -1,     0,     1,     1,    -1,    -3,    -4,    -5,    -8,    -6,    -7,     0,     3,     2,    -1,     2,     4,    -5,   -10,     5,     7,     4,    -1,    -1,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     1,     1,    -2,    -1,    -1,    -3,    -5,    -8,    -9,    -9,    -4,    -2,     2,     6,     7,     0,    -1,    -9,    -6,    -2,    -2,     0,    -1,    -1,     1,     1,     1,     0,     1,     1,     1,    -1,    -3,    -4,    -3,    -1,    -4,     2,     5,     1,    -1,     0,    -1,    -1,     0,    -2,    -4,    -1,     1,     0,    -1,     1,    -1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,    -1,     0,    -2,    -2,     0,     0,     1,     0,    -2,     0,    -1,     0,    -1,     1,     0,     1,    -1,     1,     0,     0,     0,     1,    -1,     0,     1,    -1,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     1,     0,     0,     1,     0,     1,     0,     1,     0),
		    37 => (    0,    -1,     0,     1,     0,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,     1,     0,     0,     0,    -1,    -1,     1,     0,    -1,     0,     1,     1,    -1,    -1,     0,    -1,     0,     1,     0,     0,     1,    -1,    -1,    -1,    -1,    -4,    -5,    -3,    -2,    -4,    -5,    -4,    -1,     0,     0,     0,     1,    -1,     0,     1,    -1,     1,    -1,     1,     0,    -3,    -3,     0,    -1,    -4,    -6,    -2,    -1,    -5,    -2,    -1,     0,    -1,     0,    -2,    -1,     1,     0,     0,     0,    -1,     1,     0,     1,     0,    -1,     1,    -1,    -2,    -2,    -1,    -3,    -9,    -9,    -3,    -5,    -4,    -3,    -4,    -2,    -2,    -2,    -6,    -3,    -4,    -1,    -2,    -2,     0,    -1,     0,    -1,     0,    -1,     0,     1,    -2,    -6,    -5,    -3,    -5,   -10,    -9,    -9,   -11,   -10,    -5,    -9,    -7,    -5,    -5,    -5,    -2,    -3,    -3,    -4,    -4,    -4,    -2,     0,     1,    -1,     1,     1,    -7,   -12,     2,    -4,     3,    10,     3,    -6,    -9,    -5,     4,    -3,    -2,   -11,   -13,    -9,   -14,   -12,    -6,    -6,    -6,    -2,    -5,    -1,    -1,     0,     0,     2,     2,    -1,     0,    -1,    -5,     0,    -2,    -8,    -5,    -6,    -7,    -3,    -5,   -11,    -1,     3,    -1,     0,     6,     1,    -5,    -8,    -1,    -9,    -3,     0,     2,     2,     4,     3,     1,     3,     4,     1,     0,     1,    -6,    -4,    -2,    -3,    -8,    -6,    -1,     0,   -12,    -7,    -2,    -2,    -3,    -8,    -4,    -4,    -2,    -3,     2,    -4,     1,     4,     5,     8,     3,     1,     7,    -1,     1,     3,     1,    -6,    -3,    -4,    -3,     3,    -6,    -2,     0,    -3,     1,     0,    -4,    -7,    -2,     0,     2,     0,     2,    11,     0,     1,     0,    -1,     1,    -5,     2,     7,     4,     5,     3,    -4,    -4,    -1,    -2,     1,     5,     4,     9,     2,    -6,    -4,     5,     0,     6,     3,     4,    11,     5,     5,    -4,     1,     4,     0,     4,     1,     0,     4,     5,    -1,     0,    -1,     0,    -2,    -2,    10,     4,    -7,    -1,    -4,     5,    -1,     4,    10,     8,    10,     2,    -4,    -1,    -3,     0,     2,     4,     0,     1,     2,     2,    -4,    -3,    -2,     1,    -5,     3,     3,    -3,   -11,    -9,    -2,     8,     1,     1,     1,    11,     5,     2,    -2,    -2,    -2,    -2,    -1,     1,     1,    -2,     2,     2,     1,    -4,     3,     2,    -1,     4,     6,    -6,    -6,     3,    -2,     6,     1,     4,     5,    10,     4,     3,    -3,    -3,    -6,    -4,     3,     3,    -1,    -7,     2,    -5,     0,    -2,    -2,    -3,     8,     5,     2,    -2,    -1,     7,    -3,    -3,    -2,     2,    10,    10,    -1,     4,    -3,    -6,    -4,    -1,     4,     3,    -5,   -13,    -2,    -3,     0,     4,     0,     6,     4,     5,     3,     9,     9,    -4,    -5,    -1,    -1,     1,     6,     5,    -4,     1,     1,     0,    -2,     1,     5,     0,    -7,    -8,    -1,    -5,    -5,     1,     1,     9,     3,     2,     5,     4,     3,    -6,    -3,    -2,     0,     0,     3,     2,     7,     2,    -3,     3,     3,     7,     1,    -2,   -12,    -6,    -4,     0,    -2,     1,     1,     3,     0,     7,    10,     9,     4,   -15,    -6,     1,    -1,     0,    -2,    -1,     4,     2,    -4,     0,     3,     3,    -5,    -6,   -10,    -9,     3,     2,     1,    -2,    -1,    -2,     3,     4,    10,     5,     0,   -14,    -4,    -9,     4,     1,     3,   -11,     0,     1,    -4,     2,     3,     1,    -4,    -9,   -20,    -7,     6,     4,     1,     0,    -1,    -4,     1,     3,     5,    -1,    -8,    -3,     0,    -3,     0,     4,    -1,   -10,    -2,     1,     4,     1,     0,    -2,   -12,   -22,   -18,    -6,     7,     0,    -3,     1,    -4,    -2,    -3,    -9,   -14,    -7,    -6,    -6,     0,    -1,    -1,     3,    -1,    -2,     2,     7,     5,     5,     1,   -12,   -17,   -23,    -6,    -2,     0,     0,    -1,    -3,    -4,    -5,    -6,    -7,   -10,    -9,    -1,    -5,     0,     1,     0,    -1,    -1,    -2,    -5,     4,     1,     2,    -6,   -11,   -14,   -11,     0,    -5,     1,     3,     4,    -4,    -4,    -4,    -7,    -3,    -5,    -9,    -9,    -3,    -1,     0,     0,     0,    -1,    -2,     0,     0,     1,    -3,    -8,    -7,   -12,    -6,    -2,    -3,     3,     0,     0,     1,     1,     2,     2,    -3,    -5,    -6,    -4,    -3,    -6,     1,    -1,     0,    -3,    -2,     1,     2,    -1,    -3,    -8,    -7,   -10,    -6,     1,    -1,     5,     3,    -1,     1,     6,     0,    -1,    -5,    -5,    -8,     0,    -2,    -4,    -1,    -1,     1,    -2,     0,     1,    -1,     0,    -4,    -6,    -7,    -9,    -4,     1,    -3,     0,    -1,    -1,     2,     1,     4,    -1,    -1,    -2,    -8,     0,     0,    -1,     1,     0,     1,    -2,     0,     0,    -1,     1,    -1,    -5,    -6,   -11,    -5,    -6,    -3,     4,    -1,     5,     4,     3,     5,     1,     1,     2,   -10,    -1,    -3,     1,    -1,     1,     0,    -1,     0,     0,    -1,     0,     1,     2,     1,    -2,   -10,    -7,    -3,   -10,    -4,     4,     3,     4,     7,     1,     2,     2,    -2,    -2,     1,     0,    -1,     0,    -1,    -1,     1,     1,     3,    -4,    -4,     0,     5,     4,     0,    -2,    -6,    -8,    -4,     4,     5,     1,    -6,     1,     6,     4,     5,     1,     1,    -1,     0),
		    38 => (    0,     0,     0,     1,     1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,    -1,     0,    -1,    -1,    -1,     0,     0,     1,     1,     1,    -1,     1,     0,     1,    -1,     1,    -1,     1,    -1,     1,     1,    -1,     1,    -1,    -2,    -5,    -6,    -3,    -3,     0,    -2,    -1,    -2,    -1,    -1,     0,    -1,     1,     0,     1,    -2,    -1,     0,    -1,     0,     0,    -2,    -3,    -5,    -4,     1,    -1,     0,    -3,    -2,    -3,    -1,    -1,    -4,    -5,    -6,    -3,    -1,    -2,     0,    -1,     1,     1,    -2,    -1,     0,    -4,    -2,    -6,    -6,     1,    -1,    -4,    -4,    -5,     1,     4,     4,     3,     1,    -2,    -3,    -1,    -1,     1,    -1,     0,    -3,    -1,    -1,    -1,     1,    -3,    -7,    -3,    -1,     0,     1,    -1,    -2,    -1,    -3,    -4,    -1,     2,     2,     1,     1,     1,     5,     3,    -4,    -2,    -7,    -3,    -1,    -3,    -1,     0,    -2,    -6,    -7,    -2,    -1,    -2,    -4,    -5,    -4,    -5,    -6,    -6,    -4,     2,    -2,    -1,     2,     3,     4,     1,     0,    -5,    -3,     0,     0,    -4,     0,     0,    -3,    -3,     0,     2,    -3,    -2,    -2,    -5,    -8,    -8,    -6,    -4,     1,     1,     0,     0,    -2,     4,    -3,     4,     1,     0,    -5,    -1,    -1,     0,     1,    -5,    -3,    -2,     1,    -1,    -1,     0,     2,    -1,     1,    -2,    -2,     3,     1,     2,    -1,    -4,    -2,    -1,     0,    -4,     0,    -1,    -3,     3,     5,     2,    -2,    -3,    -2,     1,     1,     1,     0,     1,    -2,     3,     3,     0,     0,    -1,     7,     6,     1,     1,    -3,     0,    -4,    -2,    -4,    -1,     5,     9,     6,     3,     1,    -2,    -1,     1,    -2,    -2,    -2,    -1,    -5,    -5,    -1,    -3,    -2,     0,     2,     5,     1,    -4,    -5,     0,    -3,    -1,     1,     6,     6,     6,     2,    -8,     1,    -1,     0,     0,    -2,    -3,    -4,    -3,    -3,     1,    -3,    -6,    -5,    -3,     1,    -1,    -2,    -3,    -6,    -3,    -1,     6,     5,     2,     0,    -8,    -4,    -8,     0,    -1,    -1,    -1,    -2,    -3,    -4,    -3,    -5,    -1,    -1,    -6,    -3,    -3,     2,    -2,     2,    -4,    -1,     1,    -4,    -1,     6,     0,    -3,    -5,     3,    -5,     1,     1,    -1,    -4,    -2,    -4,    -3,    -6,    -7,    -1,     1,     0,     1,     1,    -1,     3,    -2,     1,     2,     1,     4,     3,     0,     0,     0,    -7,    -4,    -8,     0,    -1,    -4,    -7,    -2,    -2,    -8,    -6,    -4,    -3,    -4,    -1,    -3,     2,     0,     1,     2,     5,    -2,    -2,    -5,    -4,     1,     0,     0,    -3,    -1,     2,    -1,     0,    -1,    -8,    -3,    -5,     4,     3,    -4,   -10,    -8,     1,     0,     4,     3,     1,     3,    -4,    -4,    -9,    -2,     1,     1,     1,     0,     1,    -2,    -3,    -1,    -1,     0,    -1,    -2,    -1,     7,     3,    -4,    -4,    -1,     2,     3,     2,     0,    -1,    -1,    -5,   -10,    -5,    -3,    -1,     1,    -4,    -5,     0,    -4,    -2,     1,     0,    -2,    -2,    -2,     3,     4,     1,     2,     5,     3,     4,     2,    -4,    -7,    -5,     0,    -7,   -11,    -7,    -5,    -2,    -3,    -6,    -5,     0,    -7,    -3,     1,    -2,     0,    -2,    -1,     2,     6,    10,     8,     6,     4,     0,    -5,    -3,    -5,    -3,    -6,    -1,    -5,    -4,    -4,    -7,    -4,    -4,    -3,    -1,     1,    -2,     1,    -1,     0,    -1,    -1,     4,     7,     6,     6,     3,    -3,    -5,    -9,     0,     4,    -4,    -6,    -1,     1,    -1,    -4,    -6,    -6,    -2,    -1,    -2,     0,    -4,     0,     0,    -1,    -5,     2,     8,     4,    -1,     1,    -4,    -9,    -5,    -3,     2,     0,    -1,    -4,     1,     2,    -6,    -3,    -6,    -5,    -3,    -1,     0,    -3,    -2,    -1,    -1,    -1,    -5,    -2,     7,    -1,     2,     1,    -5,    -6,    -5,    -6,    -3,    -3,    -2,    -3,    -3,    -3,    -6,    -7,    -6,    -6,    -1,    -2,    -1,    -3,     0,    -3,    -3,    -2,    -4,    -1,     6,     1,     1,     3,    -4,    -2,     1,    -4,    -4,    -3,    -6,    -5,    -3,    -7,    -9,    -8,    -7,    -2,    -2,     0,     0,    -4,     0,    -3,    -2,    -1,    -3,     1,    -1,     1,     1,     4,    -2,    -1,     1,    -5,    -5,    -3,    -6,    -1,    -4,    -6,    -4,    -7,    -6,    -3,    -1,    -2,    -1,    -3,    -1,     0,     0,     0,    -4,    -2,    -4,    -4,     1,     0,     2,     1,     0,    -2,    -1,    -3,     0,     1,    -4,    -8,    -6,    -6,    -4,    -1,    -2,    -1,    -2,    -6,     0,     0,     0,    -2,    -1,    -5,    -2,     4,     6,     5,     8,     3,     2,     1,    -1,    -5,     1,    -3,    -4,    -4,    -3,    -2,     0,     0,     0,    -3,    -2,    -2,     0,     0,     0,    -2,    -1,    -2,    -5,    -1,     4,     3,     1,    -1,     0,     2,    -2,     3,     1,    -2,    -3,    -2,     0,     0,     0,     1,     0,     0,    -1,    -3,     0,     0,     0,     0,    -5,    -1,    -4,    -5,    -5,     2,     1,     1,     0,     1,    -2,    -3,    -4,    -1,    -2,    -1,    -1,    -5,    -2,    -3,     1,     0,     1,     1,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,     0,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,     1,    -1,     1,    -1,     0),
		    39 => (   -1,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,     0,    -1,     0,    -1,     0,     0,    -1,     1,    -1,    -1,    -1,     0,     0,    -1,    -1,     1,    -1,     0,    -5,    -4,     0,    -2,    -3,    -2,    -4,    -2,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,     1,     0,     1,    -1,     1,     1,     0,    -1,    -2,    -4,    -3,    -3,    -1,     1,    -3,     0,     0,    -1,     0,     1,    -1,    -2,    -3,     0,    -1,     1,     0,     0,    -1,     0,     0,    -3,    -2,    -1,    -2,    -2,    -6,    -8,    -5,    -8,    -4,    -5,    -3,    -4,    -2,    -2,    -2,    -2,    -6,    -5,    -2,     0,    -3,    -2,     1,    -1,     1,     1,     0,    -2,    -4,    -6,   -11,    -2,    -5,    -5,     0,    -1,    -3,    -6,    -7,    -9,    -4,    -5,    -2,    -2,    -3,    -1,    -1,     0,    -1,    -8,    -1,     0,     1,     1,     1,    -1,     0,    -1,    -4,    -4,    -7,     1,     4,     0,    -1,     3,    -4,    -7,    -4,    -6,   -11,    -5,    -4,    -6,    -1,    -2,    -1,    -3,    -2,     0,    -1,     1,     0,    -4,    -5,   -10,     1,    -3,     4,     4,     6,     2,     1,     8,     1,    -5,    -8,    -6,   -11,    -4,   -10,    -4,     3,     1,    -6,    -1,    -1,    -1,     1,    -2,    -5,    -5,    -7,    -8,    -6,    -3,     1,     6,     3,     1,     0,     2,    -2,    -8,    -3,    -8,    -4,    -7,   -11,    -4,     2,     0,    -4,    -3,    -3,    -2,    -3,    -2,    -5,    -5,    -5,    -4,    -5,    -3,    -1,    -2,    -1,    -4,     1,     3,     4,    -3,    -6,    -3,    -7,    -3,    -5,    -6,     1,     0,    -2,    -3,    -1,     0,     0,    -1,    -7,    -2,    -1,    -2,     2,     6,     3,    -3,    -5,     2,     1,     3,     2,    -2,    -3,    -2,    -4,    -7,    -4,    -8,    -4,    -5,    -6,    -6,    -2,    -1,     0,    -3,    -5,     0,     6,    -3,     4,     0,     3,    -4,    -1,    -1,    -2,    -1,    -3,     2,     1,    -2,    -1,    -6,    -5,    -2,   -12,   -12,    -6,    -5,     0,    -4,     0,    -7,    -3,     4,    -1,    -1,     8,     5,    -3,    -7,    -3,    -5,    -2,     2,     2,     4,     2,     5,    -3,     1,    -2,    -4,   -10,    -7,    -6,   -11,    -1,    -4,    -1,    -6,    -4,     3,    -1,     5,     6,    -3,    -3,    -1,    -4,    -8,    -3,    -2,     3,     3,    -1,     3,     1,    -2,    -1,     3,    -5,    -4,    -1,    -7,    -6,    -3,    -1,    -6,    -3,     0,    -4,     6,     0,    -1,     1,    -1,     2,    -6,    -3,    -2,     1,    -4,    -2,     0,     3,    -1,     3,     2,    -1,    -5,     0,    -5,    -3,    -2,    -2,    -1,    -2,     6,     0,     2,     1,    -1,    -1,     5,     5,     6,     1,     2,    -3,    -9,    -5,     1,     5,    -1,    -3,     3,     1,    -1,     2,    -7,    -3,     0,    -1,    -1,    -2,     5,     3,     4,     4,    -4,     2,     2,    -1,     2,     5,    -5,    -2,    -6,    -9,    -2,     3,     2,     2,    -1,    -1,     0,     2,    -8,    -5,    -3,    -1,    -1,    -4,     1,     7,    -5,     3,    -2,    -1,    -2,    -2,    -1,     1,    -2,    -7,    -8,    -6,     1,     6,     5,    -2,    -2,    -5,    -1,     3,     0,    -4,    -7,     1,    -1,    -4,     1,     2,    -3,     1,    -4,     0,    -2,    -1,     0,     2,     3,    -3,    -4,    -2,     2,     0,     5,    -2,    -3,    -9,    -3,    -3,    -6,    -5,    -6,    -1,     1,    -4,     2,    -3,     3,     3,     2,    -3,     0,     3,     4,    -1,    -1,     4,     5,     3,    -4,     1,     3,     3,    -8,    -5,    -3,    -3,    -6,    -7,    -4,     1,    -1,    -3,     0,    -3,    -2,     2,     4,    -1,     4,     3,     3,     7,     4,     1,     0,     0,    -7,    -5,     1,     1,    -3,    -2,     2,     0,    -8,    -5,    -2,    -1,    -2,    -2,    -1,     2,    -1,    -6,    -7,     2,    -4,     0,    -4,    -6,    -4,    -4,    -7,    -7,    -7,    -2,     6,     1,    -2,    -2,     2,     9,     1,    -8,     0,     1,    -1,    -4,    -1,     1,    -1,    -2,    -7,   -12,   -12,    -5,    -3,    -6,    -6,    -9,    -9,   -11,    -6,    -4,     5,     1,     0,    -3,     1,     5,    -4,   -10,     0,    -1,     0,    -5,     3,    -1,    -2,    -2,    -3,    -7,    -9,    -3,     4,    -1,     3,    -1,    -6,    -3,    -6,     0,     1,     3,    -1,     1,     0,     4,    -7,    -5,    -1,     1,    -1,     0,     5,     1,     1,    -2,    -3,    -4,    -5,    -3,    -3,     0,     2,     1,    -1,    -4,    -3,    -1,    -3,     2,     1,    -1,     6,     8,    -6,    -4,     0,     1,     0,    -4,     0,    -1,     0,    -2,    -3,    -3,    -7,    -4,    -5,     0,     0,     0,    -3,    -2,     0,     3,     5,     9,     2,     7,    11,     2,     3,     0,    -1,     0,     0,     4,    -2,    -3,     2,    -1,    -3,    -5,    -4,    -1,     1,     0,     2,    -7,    -8,    -9,    -7,    -1,     6,     3,     2,    -1,    -4,    -3,     1,    -2,     1,     0,     1,     1,     2,     0,     0,     3,     1,     2,     0,     0,    -3,    -2,     2,     2,    -2,    -6,    -5,    -6,    -5,     0,     1,     3,     6,     4,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,     1,     0,     1,    -1,    -1,     0,     2,     2,     3,     0,    -3,    -4,     3,     2,    -3,    -7,     0,    -3,     1,     1,     0,    -1),
		    40 => (   -1,     0,     0,    -1,    -1,     1,     0,     0,    -1,     0,     1,    -1,     1,     0,    -1,     0,     0,     1,    -1,     0,    -1,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     1,     0,     0,     1,     1,     0,     0,    -1,    -2,     1,     3,     0,    -1,     2,     3,     4,     0,     0,     1,     1,     0,     1,    -1,    -1,    -1,     0,    -1,     0,     1,     3,     2,    -1,     0,     1,    -4,    -7,    -6,    -4,    -6,   -10,    -8,   -10,    -2,    -4,    -4,    -6,    -6,    -1,    -5,    -3,    -2,    -1,    -1,     1,     0,    -1,    -1,     2,     0,    -2,    -4,    -2,    -2,     0,    -1,    -3,    -3,     0,     0,    -2,    -3,    -5,    -9,   -10,    -2,    -3,    -6,    -5,    -3,    -1,    -4,     0,     1,     0,    -1,    -2,     0,    -7,    -6,    -3,    -2,     4,    -1,    -3,    -6,     0,     0,    -2,     2,    -5,    -6,    -3,    -4,    -3,     2,    -6,    -3,    -4,    -6,     0,     0,     1,    -3,     3,    -1,    -3,    -1,     0,     4,    -3,    -1,    -4,    -3,     2,    -1,    -4,    -1,     2,     0,    -5,    -6,    -5,    -1,    -4,    -3,    -3,    -5,    -4,     1,     0,    -2,    -2,     4,     3,     1,     1,    -7,    -7,    -1,    -2,    -3,     3,    -2,    -4,     1,     2,    -4,     3,    -1,     4,     2,    -8,    -4,    -9,    -5,    -2,     1,     0,    -2,    -3,     4,     4,     1,    -3,    -9,     1,    -2,    -3,     0,    -2,    -1,     0,     2,     4,     7,     7,     2,     2,     1,     3,    -6,    -3,    -9,     3,     7,    -4,     5,     0,     3,     2,    -2,     1,    -1,     0,    -2,    -2,     6,     0,     3,     2,     3,     4,     6,    -4,     0,     3,     1,     4,    -8,   -10,    -8,    -1,     0,    -1,     6,     0,    -7,    -1,    -1,    -3,     2,     0,    -4,    -3,     0,    -2,     3,     0,    -4,     2,     3,    -2,     7,    -2,     0,    -1,     1,   -11,    -9,     0,     0,    -1,     5,     0,    -4,    -6,     0,    -3,    -1,    -1,    -4,    -7,     1,     0,     4,     0,    -1,     2,     0,    -3,     6,     3,     6,    -1,     0,    -7,    -9,     0,    -1,    12,    -4,    -1,    -5,    -6,     4,     6,     2,     2,    -1,    -1,     1,    -1,     1,    -3,    -4,     1,    -5,    -2,     3,     6,     4,    -4,    -4,    -7,    -7,    -1,     1,     2,    -2,    -2,    -5,    -4,     7,     5,     2,     3,    -1,     1,     1,    -3,    -5,    -4,    -9,    -6,    -2,    -2,     3,     6,     2,     1,    -1,    -2,    -8,     1,     0,     2,     3,     4,    -2,     2,     5,     5,     8,     3,    -1,     1,    -6,    -5,    -2,   -10,    -7,    -8,     2,     1,     1,     4,     5,     4,     1,     4,    -4,    -1,     0,     1,    -1,     2,     1,     8,     6,    11,     6,     3,     0,     1,    -2,    -1,    -5,    -7,   -10,    -5,    -1,     4,     2,     0,     0,     6,    -2,    -1,    -6,     1,     0,     0,    -2,    -3,    -1,     5,     0,     4,    10,     4,    -1,    -1,    -3,    -4,    -6,    -7,    -3,    -7,    -1,     0,     4,     6,     5,     9,     6,     1,   -10,    -3,    -1,    -1,    -2,    -4,     4,    -1,     5,     7,     3,     2,     2,    -3,    -5,    -5,    -7,    -6,    -1,    -2,     2,    -5,    -2,     5,     4,     0,     3,    -3,   -11,     7,    -1,    -1,    -3,    -8,     2,    -3,    -1,     1,     4,     5,     0,    -6,   -10,    -7,    -2,     3,     0,    -2,    -5,    -4,     2,    -5,     6,    -2,     2,    -5,    -8,     8,     1,     1,    -2,    -8,    -2,    -6,    -2,     4,    10,     6,     2,    -5,    -9,    -5,     3,     1,     0,    -2,     0,    -1,     2,     0,     4,    -4,    -1,     0,    -5,    -3,     1,     3,    -3,    -3,    -2,    -4,    -3,    -2,     9,     4,     2,    -7,    -3,    -4,    -4,    -2,     1,    -3,    -1,    -5,     6,    -1,     3,    -1,    -1,    -9,    -1,    -1,     0,     3,    -6,     0,    -1,     1,    -2,    -1,     3,     5,    10,    -4,     0,    -3,    -2,    -4,    -3,    -3,    -4,    -2,    -6,    -4,    -2,    -8,    -7,    -5,     3,     1,     0,    -1,    -8,    -4,    -2,     0,    -4,    -4,     2,    -2,     0,    -3,    -4,    -5,    -4,     0,     2,    -3,    -8,    -6,    -4,    -3,     5,    -2,    -4,    -4,     4,     2,     0,    -1,    -8,    -2,    -7,    -1,     1,     1,     5,     4,     3,    -4,    -2,    -2,    -2,    -1,    -5,    -6,    -5,    -1,    -4,     1,     1,    -3,    -3,     1,     4,     3,     0,     1,    -1,    -9,    -7,    -5,     0,     1,    -1,     2,     3,     4,    -2,     0,    -3,    -3,    -3,    -4,    -8,    -4,    -8,    -2,    -5,    -5,    -5,    -2,    -4,    -1,    -1,    -1,    -1,     1,     1,     3,    -4,    -5,    -1,     5,     4,     4,     4,    -3,    -1,     2,    -4,    -8,    -5,    -5,    -5,    -5,    -7,    -6,    -1,     2,     0,    -1,    -1,     1,    -1,    -1,    -7,   -10,    -9,    -7,    -7,    -6,    -9,    -9,   -11,    -5,    -5,   -12,   -12,   -11,   -14,    -9,    -7,    -6,    -5,    -3,    -2,     1,     0,     0,     0,     1,     0,     0,    -3,    -4,    -9,    -5,    -4,    -8,    -9,   -10,    -7,    -6,    -5,    -7,    -5,   -10,    -9,    -6,    -8,    -7,    -3,    -4,     0,     0,     1,    -1,    -1,     0,     0,    -1,     1,    -1,    -1,     1,     0,     0,     0,     0,    -1,    -4,    -2,    -2,    -2,    -2,    -1,     1,     0,    -4,    -3,    -2,     0,     0,     1,     0),
		    41 => (    1,     0,     0,     1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     1,    -1,    -1,    -1,     1,     1,     1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     1,    -1,    -1,    -1,     1,     0,    -1,    -1,    -3,    -3,     1,     3,     0,    -2,    -1,     1,     1,     0,     1,    -1,    -1,    -1,    -1,     0,     0,    -1,     1,    -1,     0,    -1,     0,     0,    -2,    -2,    -4,    -2,    -3,     6,     8,    11,     9,     5,     5,    11,     8,    -7,    -7,    -5,     1,     1,     0,     1,     1,    -1,     4,     7,    -1,    -4,    -6,     5,     3,    -1,   -10,   -10,     1,     1,     1,     4,     9,     4,     4,     5,     8,     7,    -4,    -5,    -2,    -2,     1,     1,     1,     1,     1,     5,     0,     2,    -2,    -6,    -5,    -3,     1,    -3,    -7,    -8,     1,     7,     7,     3,     5,     2,     2,     4,    -4,    -3,    -2,    -5,    -5,    -4,    -1,     0,     3,     3,     1,     6,     2,    -7,    -4,    -5,    -2,    -2,    -7,    -4,    -1,     4,     7,     2,     0,    -3,    -3,     4,    -4,    -1,    -2,    -5,    -4,    -2,    -1,     0,    -5,     0,     1,     2,    -5,    -6,    -3,    -4,    -5,    -5,    -2,     1,     1,     4,     6,    -1,    -1,    -4,    -1,    -3,    -3,     0,     1,     0,    -4,    -3,    -1,    -2,    -7,    -2,    -3,    -8,    -9,    -1,     3,     3,    -3,     1,     0,    -3,     6,     1,     1,     2,   -11,    -6,    -1,    -4,    -5,    -2,     0,     0,    -4,    -5,    -1,    -2,    -6,     0,    -3,    -9,    -5,    -4,     2,    12,    -1,    -3,    -2,    -2,     2,     4,    -1,    -3,    -1,    -6,    -1,    -3,    -3,    -2,    -2,    -1,    -4,    -2,     0,     0,    -7,    -2,    -3,    -5,     0,     2,     5,     4,     2,    -4,    -4,    -2,     2,     4,     3,    -9,    -4,    -9,    -5,    -5,    -2,    -3,    -2,    -2,    -1,    -3,     1,     0,    -8,    -1,    -5,    -8,    -4,     4,    -4,    -4,    -2,    -1,     0,    -3,     0,    -1,     0,     0,    -4,    -4,    -4,    -5,    -2,    -1,    -1,    -2,    -3,     4,     0,     2,     1,    -1,    -3,    -4,     0,    -3,    -7,     1,     5,    -1,     0,    -6,     0,    -1,    -1,    -4,    -9,    -5,    -5,    -2,    -4,    -1,    -3,    -2,    -5,     1,    -1,     1,     0,    -1,    -1,    -2,    -2,    -4,    -5,     4,     0,     5,    -3,    -9,    -1,     0,     1,    -7,    -4,    -8,    -4,    -1,    -2,    -1,    -1,    -1,     1,     1,     0,     1,     1,     0,    -4,    -2,    -2,    -4,    -2,     6,     1,    -1,    -2,   -16,     1,     3,     0,    -3,   -12,    -7,    -4,    -6,    -4,    -7,    -6,     0,     0,    -1,     0,     1,     0,    -1,    -4,    -5,    -6,    -8,     5,     3,     1,    -6,   -16,    -8,     4,     0,    -3,    -7,   -11,    -9,    -8,    -6,    -6,    -5,    -1,    -2,     2,     0,    -1,     0,     1,     1,    -6,    -7,    -8,    -6,     6,     4,    -4,   -10,   -12,     1,     2,    -1,     0,    -9,   -12,   -10,    -8,    -4,    -4,    -7,    -4,    -2,    -1,    -3,     0,     1,     0,    -3,    -4,    -6,    -5,    -3,    -3,    -2,   -15,   -11,   -17,    -1,    -4,    -5,    -7,   -12,   -15,   -10,    -7,    -5,    -4,    -9,     2,    -4,    -6,    -2,     1,     0,    -1,    -4,    -1,     2,     7,    -2,    -5,    -4,    -1,    -9,   -12,    -4,    -1,    -6,    -4,    -7,     1,     5,     2,     0,    -1,    -8,     1,   -11,    -3,    -3,    -1,     0,    -1,    -1,    -3,     7,     0,    -2,     3,    -2,    -1,   -10,   -12,    -3,     1,    -1,     2,     0,     1,     3,     6,     1,    -2,    -2,     0,    -3,    -6,    -1,     0,    -1,     1,    -2,    -5,    -2,     0,     0,     3,     3,    -2,    -2,    -7,    -2,     0,     1,     6,     1,    -2,     3,     5,    -1,     1,     3,    -1,    -5,    -6,    -4,     0,     0,     1,     5,     5,   -13,    -2,    -5,    -1,    11,     2,    -1,     0,     3,     4,     3,     6,     3,     7,     5,     4,     2,     9,     5,     0,    -2,    -2,     1,     4,     4,    -2,     8,     7,     4,    -1,     3,     4,     4,     7,    -4,    -2,     4,    -1,     0,     1,    -1,     3,     1,     4,     5,     0,    -2,     2,     3,    -3,     0,     3,     2,    -3,     5,     3,    11,     7,     1,     2,     2,     0,    -1,     1,     0,    -6,     0,     0,    -1,    -1,     0,     3,     4,     4,     5,     6,     5,     2,    -1,     1,     0,     0,    -1,     0,     3,     8,    -4,    -6,     2,     0,    -3,     0,    -1,     1,     2,     0,    -2,    -7,   -17,   -14,   -10,    -3,    -5,    -5,    -5,     3,     1,     0,    -1,     0,    -2,    -2,    -4,    -2,    -3,    -2,     2,     2,    -2,     1,     0,     2,     0,    -6,    -8,    -5,    -9,    -5,     0,    -4,    -4,    -7,    -2,     1,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     2,     2,    -1,     0,    -1,    -8,     1,     2,    -5,   -15,     0,    -2,    -4,    -6,    -5,    -3,     0,     0,     1,     1,     1,     0,     0,     1,    -2,    -4,    -1,    -1,    -3,    -4,    -1,     0,    -8,    -8,     1,     3,     4,    -5,    -1,     1,     0,    -1,    -1,     1,     1,     0,     0,    -1,     1,     1,     1,     1,     0,    -1,     0,     0,     1,    -1,    -3,    -3,    -1,    -2,     1,    -2,    -4,     0,    -1,     0,     0,     1,     1,     1,    -1,    -1,     0,     1),
		    42 => (   -1,    -1,     1,     1,    -1,    -1,     1,    -1,     1,     0,     0,     0,    -1,    -2,     1,     2,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     1,    -1,     0,     1,     0,    -1,     0,     0,     1,     0,    -3,    -3,    -2,     0,    -3,    -3,     1,     0,    -1,    -8,    -3,    -2,    -2,     0,    -1,    -1,     0,     0,     1,     0,    -1,    -3,    -2,     0,     0,    -2,    -1,     0,     6,     6,     1,     2,     3,     3,     6,     7,     2,    -1,     0,    -2,    -3,    -2,     1,     1,    -1,     0,    -1,     1,     0,    -5,    -5,    -3,    -1,    -3,     3,     3,     7,     0,    -2,    -1,    -2,    -1,     1,     6,    -5,    -1,    -1,     3,     0,    -3,    -1,    -2,     0,     1,     0,    -1,    -2,    -4,     0,    -2,    -2,    -1,     5,    11,     5,     0,     5,    -2,    -2,    -1,     4,     2,     2,    -1,    -6,    -4,    -1,    -4,    -5,    -3,    -8,    -4,    -1,     0,    -1,     0,    -1,     0,     2,     3,     0,     1,     3,     8,     3,     6,     6,     3,     6,    -2,    -2,     4,     2,     0,    -5,    -5,    -4,    -1,   -11,    -4,     1,     1,     2,    -3,    -2,     4,     4,     7,     3,     2,     3,     2,    -1,    -3,     2,     4,     5,     2,     5,     0,     2,     5,    -3,   -11,   -12,    -1,    -9,    -2,     1,     0,     4,    -2,    -1,     3,     4,     5,     2,     1,    -3,    -2,     5,     4,    -1,     4,     4,     2,     0,    -3,    -2,     1,    -5,    -7,     1,     5,   -13,    -6,    -3,     5,     5,    -2,    -1,     1,     2,     1,    -2,    -1,    -3,     2,    -3,    -3,    -2,    -5,     1,    -3,    -4,    -2,    -6,    -3,    -1,     7,     4,    -2,    -9,    -5,     1,    -6,     6,     2,     1,     1,     1,     0,     1,     3,     4,     0,    -3,    -4,    -5,    -2,    -2,    -1,    -7,    -5,    -2,     1,    -2,     5,    -1,    -7,    -3,    -2,    -1,    -2,     6,     0,     2,     1,     0,    -1,    -3,    -1,     1,     2,     7,    -1,    -2,    -1,    -1,     2,    -5,    -4,    -3,    -3,    -6,    -6,    -3,    -4,    -2,    -4,     0,    -3,    -2,    -4,     0,     2,     0,    -2,    -1,    -5,     0,     2,     4,    -5,     0,     3,     0,    -2,    -7,    -1,     2,     0,    -3,     1,    -3,     3,    -5,    -7,     1,    -3,    -8,    -2,     0,    -1,     1,    -3,     3,     8,     4,     2,     5,    -4,     1,     1,    -2,    -1,     0,     6,    -2,     3,     6,     4,    -1,    -1,     0,     0,     0,    -1,    -4,    -5,    -1,     0,     4,     4,     5,     2,     0,    -2,     0,     0,     0,    -2,     1,     2,     5,     7,     4,     5,     5,     2,    -2,    -4,     6,     1,     0,    -4,    -1,    -1,    -5,    -6,     1,     9,     6,     1,    -3,    -2,    -4,    -4,    -6,    -3,    -3,     0,     8,     6,     4,     7,     8,     9,     8,     2,     5,     5,     1,    -3,     5,     2,    -5,    -3,     0,     2,     7,     3,    -4,     2,    -2,    -9,    -8,    -3,    -2,     1,     1,     7,     8,     6,     4,     6,     1,     1,     1,     4,     0,     0,     5,    -3,    -5,    -5,    -2,     5,     3,     3,     2,     3,    -4,    -6,    -5,     5,     1,     2,     9,     9,     8,    10,     5,    12,     4,     5,     7,     3,     0,     0,     5,    -1,    -6,    -3,    -3,    -1,     5,     7,     7,     4,     3,    -2,     0,     3,    -4,     0,     7,    11,     6,     2,     2,     2,    -2,    -4,     5,     4,     0,     0,     1,    -2,    -3,    -2,    -1,     1,     2,     6,    10,     4,    -1,    -2,    -4,    -2,     0,     6,    10,    12,     9,     3,     2,     3,     3,    -5,    -2,     6,     1,    -2,    -4,    -1,    -1,     0,    -1,     1,     3,     7,     5,     3,     2,    -7,    -1,     1,     0,    15,    17,    14,     6,     3,     4,     2,     1,    -6,     0,     4,     0,    -3,     1,     2,     1,    -5,    -6,     1,     4,     1,     5,     4,     4,    -2,    -4,     2,    12,    11,    11,     8,     4,     0,    -4,     1,    -1,    -1,    -3,     0,    -1,    -1,     4,     0,     6,    -2,    -6,     1,     0,    -3,    -2,     0,     0,     2,    -1,     8,    13,    12,     9,     9,     2,    -1,    -1,    -3,    -5,    -2,     0,     1,    -1,    -1,    -2,     1,    -3,     0,    -5,    -3,     0,    -3,    -2,     0,     5,    -1,    -1,     8,    17,    11,    15,     5,     3,    -1,    -1,    -2,     0,     4,     0,    -1,     0,     1,    -1,    -1,    -3,     0,    -2,     0,     3,    -3,   -10,    -6,     0,     1,     7,    14,    19,    15,    12,     6,     0,     4,    -4,     0,     3,     3,    -4,     1,    -1,     1,    -3,    -4,   -13,   -13,    -4,    -3,    -1,    -9,    -7,    -5,    -4,     6,     9,     7,    13,    13,     9,     3,     0,     0,    -3,    -2,     3,     0,     2,     1,     1,     1,     0,    -2,    -5,    -9,     6,     2,    -1,    -3,     0,     6,    10,    12,    13,    13,     9,     4,     5,     2,    -2,    -3,    -8,    -1,     1,     3,     2,     0,    -1,     1,    -1,     0,    -2,    -6,   -10,    -9,    -9,   -10,   -10,    -5,    -7,    -7,    -9,    -7,    -7,    -7,    -6,    -8,    -3,    -3,   -10,     0,    -1,     0,     1,     1,    -1,     0,     1,     1,    -2,    -1,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -2,    -2,    -1,    -5,    -8,    -1,    -2,    -1,     1,    -1,    -1),
		    43 => (   -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,    -2,     0,     1,     0,    -1,     0,     1,     0,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -3,    -2,    -4,    -4,    -8,   -11,   -12,    -4,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,    -1,     1,     0,    -1,    -2,     1,    -3,    -4,    -8,    -8,    -2,     0,    -1,    -1,     0,     0,     2,    -1,    -4,    -3,    -5,    -6,    -6,    -7,    -3,     0,     0,     0,     0,     0,     0,    -3,    -2,     1,     0,     2,     5,    -2,     0,     2,     7,    -1,     0,     7,     8,     6,     3,    -4,     1,    -4,    -6,   -13,   -11,    -4,     1,     0,     0,     6,    -9,     2,     3,    -3,    -6,    -7,     2,     4,     6,    -2,     0,     0,    -1,     1,     4,    -2,    -3,    -6,    -5,    -1,     7,    -6,   -13,   -12,    -3,     0,     0,     0,    -2,     2,    -2,     0,     2,     2,    -1,     1,    -1,     1,    -1,     3,     1,     2,     4,    -2,    -8,    -1,     3,    -2,    -4,     7,    -2,   -14,    -5,    -1,    -1,     1,    -5,    -2,    -6,     1,     5,     4,     1,     1,    -1,    -6,    -6,     0,     3,     5,     3,     7,     4,     3,     3,     5,     2,     2,     8,   -12,   -10,    -5,     0,    -1,    -1,     1,     1,     0,     1,     2,     0,    -1,    -4,    -2,    -1,     2,     2,     1,    -3,     4,     5,     2,    -2,     2,    -2,    10,     5,   -17,   -10,    -6,    -4,    -1,     3,     4,     1,     0,    -2,     1,    -1,    -2,     2,    -1,     5,     4,    -3,    -6,    -1,     2,     3,     6,     1,    -5,     5,     5,     1,   -19,   -12,    -1,     0,    -7,     0,    -2,     3,    -1,    -5,    -7,    -6,     0,    -7,    -1,    11,     8,     3,     1,     4,     1,    -1,     2,     5,     0,     8,     5,    -9,   -15,   -13,    -5,     1,    -7,     1,     3,    -4,    -4,    -8,    -8,    -9,   -10,   -11,    -3,     7,    10,    13,     4,    -3,    -2,    -4,    -3,     0,     3,     1,     2,    -9,    -6,    -9,    -5,    -1,    -4,    -1,     5,     1,    -4,   -11,   -10,    -5,    -8,   -14,    -3,     2,    11,     7,     6,     2,     1,    -1,    -4,    -2,    -4,    -5,    -9,   -24,   -12,    -8,    -1,     0,    -2,     1,     0,    -2,     0,    -5,    -8,    -3,   -13,    -3,    -6,     2,     6,    15,     7,    -1,     3,     3,    -3,     0,    -2,   -14,   -17,   -18,    -9,    -6,    -1,     0,    -1,   -15,    -3,    -4,    -4,    -2,    -4,    -1,    -5,    -6,    -3,     1,     5,    10,     4,     9,     2,     3,     2,     1,    -4,   -10,    -4,   -10,   -10,    -7,    -1,    -2,     4,     1,    -9,    -9,    -6,    -4,    -5,    -4,    -2,    -7,    -2,     0,     5,     4,     6,     2,     0,    -6,    -4,    -5,    -7,    -3,     1,    -8,   -10,    -5,    -2,     0,     2,     0,    -6,    -1,    -1,     2,    -1,     2,    -8,    -8,     2,     8,     8,     6,     8,    -2,    -8,    -9,    -4,    -3,    -1,     4,     4,     4,    -7,     1,    -4,     0,     1,     2,     4,     1,    -3,     0,     1,     0,    -4,    -1,     4,     3,     2,     6,    -2,   -10,    -5,    -3,    -1,    -5,    -4,     6,     1,     4,   -13,    -9,    -4,     0,     2,     3,     4,     2,    -5,    -2,    -2,    -6,    -4,    -1,     6,     1,     3,    -1,    -6,    -8,    -5,    -5,    -2,    -7,    -2,     1,     1,     0,   -10,    -2,    -4,    -3,     1,     4,     6,     0,    -1,     2,     4,    -3,    -2,     5,     7,     0,     0,    -3,    -4,    -2,     1,    -3,     1,     2,     3,    -3,    -3,    -5,    -9,    -2,    -5,     0,    -4,     3,     9,     4,     7,    -3,     4,     0,     2,     6,     2,    -5,    -4,    -7,     1,     1,     3,     3,     1,     2,     2,    -4,    -2,    -3,    -7,    -9,    -5,     0,    -4,    -6,     2,     0,    -5,    -5,     3,     4,     1,     4,     2,    -7,    -2,    -2,     4,     4,     2,    -1,    -2,    -1,     2,    -3,     0,    -5,    -6,    -1,     0,    -1,    -1,    -4,     2,     0,    -7,     0,     5,     5,    -2,    -4,    -4,    -3,     1,    -2,     0,    -1,     0,    -1,     0,    -3,    -3,     0,    -5,   -11,    -7,    -3,    -1,     0,     0,    -2,     2,    -5,    -3,     5,     0,    -4,    -2,    -2,    -2,    -1,     1,     0,     0,    -1,     1,    -2,    -2,    -1,     1,     0,    -8,   -10,   -13,    -1,     0,     0,     0,     3,     8,    -2,     1,     6,     2,     4,     1,     6,     3,    -4,     3,    -4,     0,     4,     0,     4,    -1,    -3,    -4,    -5,    -7,     7,     1,    -4,     1,     1,    -1,     3,     8,    -2,     0,     2,     1,    -3,    -4,     1,    11,    -6,    -1,     7,    -2,    -2,    -3,     0,     0,    -1,    -1,    -3,    -3,    -7,    -6,    -3,     1,     1,     0,     1,    -4,    -5,    -4,    -6,     2,     3,     0,     9,     8,    13,     4,    -1,    -4,     4,     0,     2,     5,    -5,   -11,   -13,   -14,    -6,    -1,    -2,     1,     0,     1,     0,    -4,    -9,    -4,    -5,    -2,    -1,    -2,     4,     2,     5,     1,    -8,    -4,    -1,     1,     2,    -4,    -3,    -7,   -10,    -7,     0,     0,    -1,    -1,    -1,    -1,     1,     1,    -2,    -3,    -3,    -2,    -2,    -7,    -7,    -8,    -6,   -12,    -5,    -5,    -4,    -2,    -2,    -7,    -8,    -4,     0,     1,     0,     0,     0,    -1),
		    44 => (    1,     1,     1,     1,    -1,    -1,     1,     1,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     1,     0,     0,    -1,    -1,     1,     1,     0,     1,     0,     1,     1,    -1,     0,    -1,    -1,    -2,     0,    -1,    -6,    -2,    -8,    -7,    -1,    -4,    -3,     0,    -1,    -1,    -4,    -1,    -1,    -2,    -1,    -1,     0,     1,    -1,    -1,    -1,    -6,    -7,    -8,    -3,    -6,    -5,    -4,    -2,    -8,     2,     1,    -4,    -9,    -6,    -5,    -5,    -2,    -2,    -3,    -4,    -1,    -1,    -1,     1,    -1,    -1,    -1,     0,    -8,   -13,    -7,    -7,    -7,    -8,    -5,     4,    -3,    -8,   -15,    -9,    -1,    -2,    -1,    -6,    -7,    -1,    -2,    -5,    -3,     0,    -3,     0,     1,    -1,     1,    -1,    -5,    -2,     2,     2,     0,    -1,     0,    -7,   -11,    -1,     2,   -10,   -13,   -14,   -13,    -7,    -2,    -1,     0,     2,     4,     6,     2,    -4,    -2,     0,     1,    -1,    -1,    -1,     0,    -2,    -2,    -7,   -11,    -9,     1,     7,    -3,    -5,    -2,    -6,   -24,   -13,     1,     6,     2,     1,     0,     0,     0,    -3,    -2,    -1,     0,     0,    -5,     4,    12,    -2,    -8,    -5,    -3,    -6,     2,     6,     2,    -4,    -5,   -17,   -19,    -8,     6,     4,     2,     0,     4,     5,   -12,     4,   -10,     0,    -9,    -1,    -4,     2,    10,    -5,    -3,    -2,    -1,     2,     3,     0,     4,    -2,    -9,   -20,   -19,    -1,     6,     3,    -2,     0,     3,    -2,    -3,     4,   -11,    -4,    -7,     2,    -2,     0,     2,    -4,     2,    -4,     0,    -3,    -1,     4,     3,     1,   -10,   -25,    -7,     3,     3,     2,    -2,     5,    -5,     0,     7,     3,    -7,     1,    -6,     1,    -3,    -1,     2,    -3,    -2,    -3,     1,    -1,     1,     6,     6,     4,   -12,   -13,     3,     6,     2,     3,     2,     3,     2,     7,    -6,    -6,    -4,     1,    -4,    -6,     2,     4,     6,     0,    -3,    -1,     2,    -2,    -2,    -1,     8,    -3,   -14,    -9,     2,     6,     5,     1,    -1,     2,     4,     2,   -11,    -4,    -1,    -1,    -3,    -3,    -8,    -3,     3,     6,    -1,     3,    -3,     2,    -1,     6,    -3,    -9,   -13,    -8,    -3,     1,     1,    -6,     4,     0,    -1,     4,    -6,    -6,    -4,    -1,     0,    -6,    -7,   -10,    -3,     2,     5,     4,    -4,    -1,     4,     5,     3,   -11,    -6,    -2,    -1,    -2,     4,     0,     6,     1,     4,    -7,    -6,   -12,    -7,     1,    -2,    -7,    -7,    -9,    -5,    -1,    -1,     3,     3,     4,     6,     1,     2,     1,     2,     2,     4,    -3,     4,     4,     2,    -1,    -3,   -12,   -10,    -9,     0,    -1,    -1,    -2,    -8,    -6,    -1,    -1,     0,    -1,     3,     1,     4,     1,    -2,     4,     1,     0,     0,    -2,     4,     2,    -3,    -3,    -2,    -6,    -6,    -7,     0,     0,     0,    -1,     2,     0,     0,     0,    -1,     3,     1,     4,     3,     0,     1,     3,     0,    -2,    -1,     0,     7,   -12,    -4,    -2,    -1,    -6,    -9,    -6,     0,     0,    -1,    -3,     2,     0,    -2,    -8,    -1,     1,     1,     0,     0,    -1,     0,    -3,     1,    -1,    -2,    -2,    -3,    -9,    -5,    -3,    -5,    -7,   -10,   -10,    -2,    -1,     0,    -4,     2,     5,    -1,    -6,    -3,    -4,    -2,    -2,    -2,     0,     0,    -2,     1,    -3,     2,    -1,    -6,   -10,     2,    -2,    -2,    -7,     1,    -2,    -3,    -5,     1,    -5,     8,    11,    -5,    -3,    -6,    -5,    -6,   -11,     0,    -4,     1,     1,    -1,     1,    -5,     0,    -2,     1,     5,     2,     2,     0,     4,    -1,    -1,     0,    -6,    -3,     7,     4,    -5,    -7,    -4,    -2,    -6,    -6,    -1,    -5,     1,    -1,    -3,    -1,     1,    -2,    -2,    -2,     2,     1,     2,     5,     3,    -1,    -2,     1,     0,    -2,    -9,    -8,    -9,    -8,    -5,    -6,     0,    -3,    -4,    -5,     0,    -2,    -3,     1,    -1,    -3,    -3,    -8,    -7,    -5,    -3,    -8,   -11,    -2,     1,     1,     0,    -2,    -5,    -8,    10,    -1,     2,     6,     8,    -2,    -1,     0,    -1,    -2,    -2,    -1,    -9,    -7,     1,     1,    -1,     1,     3,    -4,   -15,    -5,    -1,    -1,     1,     1,    -6,   -10,     6,     6,     4,     4,     0,     4,     0,     0,     0,    -3,    -2,     0,    -4,    -7,    -3,     0,     1,     0,     4,    -5,    -5,     2,     1,     1,     0,     0,    -5,    -8,   -16,     3,     4,     3,     3,     2,     0,     2,    -2,     2,     2,     5,    -3,    -3,    -2,    -1,     3,     1,     3,    -3,     1,     3,     1,     1,     1,    -1,    -2,   -12,   -10,    -2,    -5,     0,     2,     3,    -2,     1,     0,     0,     5,     2,    -6,   -13,    -3,    -2,     4,     2,     4,    -5,     5,    -4,    -1,     1,    -1,    -2,    -1,     0,    -7,    -7,     0,    -1,    -4,     0,     1,     2,     4,     0,    -5,    -5,   -11,    -7,    -5,    -1,    -2,     3,     7,    -1,    -3,    -1,     0,     0,    -1,     0,    -6,     1,    -7,    -6,   -11,    -5,    -7,    -7,    -5,    -9,   -13,   -15,   -20,    -4,    -5,    -8,    -4,    -5,    -5,    -4,     3,     0,    -1,     0,    -1,     0,     0,     0,     1,     1,     0,    -3,    -5,    -4,    -3,    -7,    -8,    -1,    -5,    -7,    -1,    -6,    -8,    -4,    -4,     0,    -1,     1,     0,    -1,     1,     1,     0),
		    45 => (    0,    -1,     0,     0,    -1,    -1,     0,    -1,     1,    -1,     1,     1,     1,    -1,    -1,     0,    -1,    -1,     1,     1,     0,    -1,    -1,     0,    -1,    -1,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,    -2,    -2,    -2,    -3,    -5,    -6,    -4,    -6,    -6,    -6,    -5,    -1,     0,     0,     0,    -1,     1,    -1,    -1,    -2,    -2,    -3,    -1,    -1,    -1,    -7,    -2,    -3,    -2,    -5,    -6,    -6,    -6,    -2,    -3,    -4,    -4,    -3,    -5,    -5,     3,    -8,    -1,     0,    -1,     1,     0,    -1,     5,    12,    -2,    -5,    -6,    -2,     3,    -2,    -8,    -6,   -10,    -8,    -4,     3,     1,     1,    -1,     0,     2,    -8,    -7,     0,    10,     9,     1,     0,     1,    -3,     9,     0,     0,    -6,    -5,    -4,    -1,    -1,    -9,   -10,    -7,    -5,    -4,    -7,    -6,     0,     6,    -1,     0,    -6,     0,     8,     6,     1,    -3,     1,     0,    -6,    10,    -2,    -2,    -3,    -6,    -5,    -3,     0,     0,    -8,    -3,    -3,    -2,    -4,    -1,    -1,     4,     1,    -1,    -3,    -2,    -3,     2,     0,    -3,    -1,     0,    -5,    -2,    -3,    -2,    -4,    -6,    -3,    -1,    -1,    -6,     0,     1,    -1,     0,    -1,    -5,     0,    -2,    -3,    -5,     8,     6,     4,     8,     9,     0,     0,    -1,     1,    -3,    -2,    -5,    -4,    -5,     1,    -2,     0,    -1,     3,     4,     4,     2,     4,     5,    -1,    -4,     0,     3,     3,     3,     2,    -1,    10,     2,    -3,    -1,    -5,    -2,    -3,    -4,    -3,    -2,    -2,     0,     0,    -1,    -2,     0,     3,    -1,    -2,     1,     1,     9,    11,     5,     7,     6,     2,    -1,     4,     5,     1,    -2,   -10,    -7,    -3,    -4,    -5,    -3,    -2,    -3,    -4,    -1,     2,     0,     2,     0,    -1,     2,    -2,    -6,     3,     1,     3,     5,    13,    10,     2,     2,     0,    -1,    -5,    -5,    -6,     3,    -3,     0,     1,    -3,    -4,     0,     4,    -1,     0,     2,     4,    -6,   -20,   -22,   -12,   -10,   -11,    -4,     0,     3,     1,     4,     0,     1,     0,     4,     2,     3,    -2,    -2,    -5,    -9,    -2,    -6,    -7,    -4,     0,    -1,     1,    -1,   -11,   -13,   -19,   -17,   -17,   -14,   -11,    -2,     0,    -2,     1,     0,     0,     6,     3,    -1,    -6,    -9,    -8,    -6,    -2,    -6,    -8,     0,     3,    -2,    -3,     2,     0,    -2,    -8,   -14,   -13,   -23,   -15,    -7,    -1,    -4,    -1,    -1,     0,     7,    -1,    -3,    -2,    -3,    -4,     0,    -2,     0,     5,     1,     2,     2,    -1,     1,     3,     6,     4,     4,    -1,    -8,   -12,    -3,     1,    -5,     1,     0,    -2,     4,    -5,    -7,    -1,    -5,    -6,    -1,     0,     3,    -1,     1,     1,     5,     4,    -4,     0,     2,     6,    -2,     0,     5,     3,    -4,    -2,    -4,     1,     0,    -5,     1,    -4,     0,     3,    -1,    -3,    -7,    -2,    -3,    -3,     4,     0,    -5,    -3,    -1,    -3,    -2,     6,    -1,    -2,     5,     8,     0,    -1,    -1,    -1,    -3,    -9,     0,     1,    -6,     6,     1,     1,   -10,    -8,    -9,    -5,    -2,    -1,    -3,     3,     2,     0,     0,     7,     5,     0,    -4,     1,     3,    -2,    -2,    -1,    -4,   -11,    -4,     5,    -1,     6,    11,     4,     1,     1,    -6,   -11,    -5,    -6,    -5,     0,     0,    -1,    -3,     4,     0,    -9,    -7,    -2,    -1,    -4,    -2,    -1,     0,    -9,    -1,     1,     2,     3,     8,     5,     1,     2,    -3,     0,    -3,     0,     0,    -1,     1,    -3,    -4,    -3,    -2,    -5,    -9,    -6,    -3,    -7,    -6,     1,    -2,     7,    -8,    -3,    -1,     4,     7,     5,     7,     3,     5,     5,     4,     2,    -1,    -2,    -3,     2,     3,    -2,    -4,    -4,    -6,    -4,    -3,    -4,    -5,     1,    -1,     6,   -10,    -7,    -1,     0,    -4,     2,     3,     4,     3,     3,    -1,     1,     0,    -1,    -1,    -1,    -2,    -2,    -4,    -2,    -2,    -2,    -2,    -1,    -1,    -1,     0,    -3,     0,    -5,     3,    -3,    -1,    -7,    -4,    -3,     3,    -3,    -1,     2,     0,     2,     2,     2,    -3,    -5,     0,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,   -10,     3,     4,     0,    -5,     0,    -6,    -3,    -3,    -1,     0,    -2,     1,     1,     0,     0,     0,    -4,     0,     3,     1,    -1,    -1,    -1,    -1,     1,     1,    -1,     1,     2,     6,     8,     1,    -4,    -5,    -5,    -1,    -1,    -5,    -6,    -1,    -3,     0,     3,     4,     0,     0,     3,     2,     0,    -4,    -2,    -1,    -1,    -1,     0,    -5,     0,    -1,    -2,    -6,   -10,    -9,    -4,   -10,   -13,    -4,    -1,    -4,    -5,    -7,    -4,     1,     4,     3,     0,     3,     1,     2,    -6,    -2,     0,     1,     1,     0,     2,    -4,    -3,     0,    -2,    -7,    -2,   -11,   -11,     1,    -3,    -3,    -2,     0,    -2,    -1,    -1,    -1,    -4,     2,     0,     1,     1,    -1,    -1,     1,     1,     1,    -1,    -2,    -3,    -4,    -2,    -3,    -3,    -2,    -3,    -2,     4,     9,     8,     7,     4,    -1,     5,     0,    -2,     0,    -1,    -1,     1,     1,     0,     0,    -1,     1,     1,     0,    -2,    -1,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -2,    -2,    -2,    -2,    -6,    -1,     0,     0,     1,    -1),
		    46 => (   -1,     1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     0,     0,     1,    -1,     1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,     1,     0,     1,     1,    -1,     1,     0,    -1,     0,     0,     3,     5,     7,     7,     4,     2,     1,     2,     2,     1,     0,    -1,     2,     2,     9,     3,     2,     2,     0,     0,    -1,     0,     0,     0,     1,     1,     1,     0,     5,     7,     7,     4,    -2,    -2,    -2,     0,    -1,    -1,    -1,    -3,    -1,     4,     4,     1,     2,     4,     4,     1,    -1,     0,     0,    -1,    -6,    -4,     0,     1,     3,     5,     2,     4,     0,    -5,    -6,    -2,    -1,    -1,    -1,    -1,    -1,     2,     0,     4,     0,     5,     6,     0,    -2,     0,     0,    -1,    -3,    -1,     0,     1,     1,     1,     1,     1,    -4,    -3,     0,    -3,    -2,     3,     2,     0,    -1,     0,    -1,     2,     0,     2,     1,     0,     3,     4,    -1,     1,     1,    -2,     1,    -2,    -1,     1,     1,    -3,    -5,     1,     0,    -3,     2,    -2,    -4,     1,     1,     1,     2,     0,     1,     3,     3,     1,     6,     4,     0,     0,     0,    -1,    -1,    -1,    -2,     1,     0,    -2,     1,    -1,     1,    -3,    -4,    -5,    -6,    -1,     1,     2,     3,     5,     3,     2,     0,    -4,     2,     2,    -1,     0,     1,    -2,     0,    -1,    -3,    -3,     2,     1,     0,    -2,    -6,    -3,     2,     0,    -3,    -2,    -3,    -1,     0,    -1,    -2,    -1,     3,    -2,     1,     2,     1,     1,    -1,    -4,    -1,     0,    -2,    -4,     2,     2,    -1,    -6,    -4,    -1,    -1,    -4,     2,     3,    -3,    -3,    -5,    -2,    -7,    -6,    -4,    -5,    -2,    -5,     0,     1,    -1,    -1,    -2,    -5,     0,     0,     3,     1,    -2,    -4,    -4,    -4,    -1,     2,     0,    -1,    -4,    -7,    -7,    -6,    -9,    -7,    -2,    -3,     1,    -1,     0,     0,     0,    -2,    -1,    -4,     0,    -2,     3,    -4,    -4,    -6,    -3,    -4,    -1,     2,    -1,    -5,    -6,    -3,    -6,    -4,    -6,    -6,    -2,    -2,    -2,    -3,     0,     0,    -1,    -1,     0,     1,     4,     0,     1,    -3,    -7,    -4,    -2,     0,     3,     0,    -6,    -7,    -5,     0,     1,     0,    -1,    -2,     1,    -4,    -2,     0,     1,    -1,     0,    -1,    -3,     2,     1,    -2,    -1,    -3,    -6,    -3,    -2,     2,    -1,    -4,    -4,     3,     2,    -1,     1,     3,     2,     2,     2,    -5,    -6,    -1,    -1,     1,    -1,    -1,    -2,     3,    -1,     1,     3,    -5,    -6,    -3,     2,     2,    -4,    -2,     0,     0,     2,     2,    -1,    -1,     0,     3,     4,    -4,    -3,     1,    -1,    -1,     1,    -1,    -1,     5,    -1,     1,     1,    -4,    -4,     4,     2,    -1,    -4,     0,     1,     4,     4,     4,     0,    -4,    -1,     3,     3,    -1,    -2,    -3,     0,     1,    -2,    -1,    -1,     3,    -1,     0,     0,    -2,    -4,    -1,    -2,    -5,    -2,     2,     4,     3,     4,     5,    -1,    -2,    -2,     4,     4,    -2,    -3,    -5,    -1,     1,    -1,    -2,    -1,     2,    -1,    -4,     1,    -3,    -2,    -2,    -5,    -1,     1,     1,     2,     4,     0,    -3,    -1,    -1,     0,     0,     0,    -1,    -2,    -5,     0,     1,    -2,     0,     0,    -4,     0,    -5,     1,     0,    -2,    -7,    -6,    -1,     2,     1,    -1,     0,    -1,    -2,     3,     2,    -1,    -1,     0,     0,    -2,    -5,     0,    -1,    -2,     0,    -1,    -3,    -5,    -3,     3,     2,    -1,    -4,    -2,     2,     0,     1,     0,    -3,    -2,    -2,     4,     0,     0,    -3,    -2,     0,    -5,    -4,     0,    -1,     0,     0,    -1,    -4,     0,    -1,    -1,     1,    -3,     1,     0,    -2,     1,    -3,     0,    -2,     0,    -2,     2,    -1,    -1,    -1,    -1,    -2,    -2,     0,     1,     0,     0,    -3,     1,    -2,    -2,    -1,     0,    -2,     2,    -1,    -4,    -3,     1,    -1,    -5,    -2,    -1,     1,     3,     2,    -2,    -4,    -1,     1,    -2,     0,    -1,     1,     0,    -2,     0,    -3,    -3,     1,    -1,     2,    -1,     0,    -3,    -4,    -2,    -3,    -2,    -2,    -1,     1,     2,    -2,    -5,    -2,    -3,     1,    -1,     0,     0,     0,     1,    -1,     0,     0,     2,     0,     0,    -2,     0,    -3,    -1,    -2,    -3,     0,     0,    -1,    -4,    -2,    -3,    -2,    -5,    -3,    -2,    -2,     1,    -1,    -1,     0,     0,    -2,     1,     0,    -2,    -2,     2,     2,     1,     2,     3,    -3,    -2,    -3,     2,    -1,    -3,    -5,    -3,    -5,    -2,    -1,    -2,     0,    -2,     1,    -1,     0,    -1,     0,    -2,     0,    -2,    -3,    -2,    -3,    -2,     0,     0,    -3,    -2,    -4,     0,     0,    -1,    -5,    -5,    -1,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     0,    -1,     1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,    -4,    -1,    -2,    -4,    -1,    -1,     1,     0,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,    -1,     1,     0,    -1,    -1,    -1,     0,    -1,    -3,    -1,     0,     1,     1,     1,     0,     1,     1,     0,     1,     0,     0,     1,     0,     0,    -1,     0,    -1,     1,     1,    -1,    -1,     0,     1,     1,     1,     0,    -1,     0,     0,    -1,     0,     1,     1),
		    47 => (    0,     0,     1,    -1,     1,     0,    -1,     1,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     1,    -1,     0,     1,    -1,    -1,     0,     0,    -1,     1,     1,     1,     0,    -1,     1,    -1,    -7,    -5,    -6,    -2,    -1,    -3,    -2,     1,     1,     1,     0,     1,    -1,     0,    -1,     0,    -1,     1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -5,    -7,    -5,    -4,    -3,    -1,     1,     0,    -1,    -1,     0,    -2,     0,    -1,     0,    -1,     1,     0,     0,     1,    -2,    -3,    -1,    -2,    -4,    -3,    -2,     0,    -2,    -4,    -2,     0,    -5,    -5,    -3,    -2,    -1,    -2,     0,    -4,    -1,    -1,     1,    -1,    -1,     1,    -1,     1,    -1,    -1,    -4,    -4,    -4,    -6,    -3,    -4,    -6,    -7,    -5,    -4,    -5,    -4,    -5,    -3,    -1,    -3,    -2,    -6,    -4,    -3,    -2,    -1,     0,    -1,     1,    -1,    -3,    -3,    -6,    -8,    -5,    -1,    -2,    -6,    -1,     2,     0,    -5,   -10,   -11,    -7,   -10,   -13,   -11,    -7,    -7,    -6,    -5,    -2,     0,     1,    -1,     0,     1,     1,    -3,    -7,    -9,   -11,   -10,   -14,   -12,    -3,     4,     5,     1,    -4,    -7,     2,     3,     0,     2,     9,     2,     5,    -6,    -2,    -6,    -1,    -1,     5,     3,     5,     2,    -2,     5,     0,    -5,   -12,   -11,   -11,    -8,    -2,    -1,    -6,     0,     0,     3,    -4,    -8,    -4,    -3,    -2,    -1,     1,    -3,    -2,    -3,     6,    -3,     0,    -1,     0,     5,     5,    -4,   -10,   -10,    -9,    -5,    -8,    -8,    -9,    -6,    -4,     2,    -4,    -5,    -8,    -3,     5,     2,     0,    -9,    -3,    -2,     5,    -3,    -3,     0,     2,     8,    -1,     1,    -3,    -7,    -3,    -4,    -8,    -1,    -1,    -1,     0,     1,    -4,    -3,     7,     5,    10,     6,     2,    -6,     1,    -1,     3,     1,    -1,    -7,    -2,     3,     0,    -4,    -2,     0,    -1,     1,     4,     2,     0,    -2,     5,     3,     3,    -1,     5,     4,    -1,    -4,    -1,    -7,     2,    -1,     2,     1,     0,     0,     1,    -2,     6,    -2,     0,    -1,     8,     6,     4,     4,     0,    -3,    -3,     1,     3,     2,     3,     2,     3,    -2,    -4,    -1,     8,     0,     0,     2,     5,     4,     4,    -4,     5,     6,     0,     1,     6,     8,     2,    -4,    -4,     3,     5,     1,    -2,     0,    -2,     4,    -1,     7,     5,     9,     9,     1,     2,     4,     6,     4,     2,     2,    -6,    -2,     1,     4,     1,     0,    -4,    -4,    -4,     3,    -1,    -1,    -1,     6,     3,     4,    -7,     7,     6,     4,    -2,    -2,     5,     8,     6,     2,    10,     1,    -7,     3,     3,     5,    -1,   -10,   -13,    -4,    -4,    -2,    -4,     5,     1,     3,     3,     2,     1,     1,    -2,    -6,    -1,     1,    -1,     0,     8,    -6,     3,    -1,     4,     0,     5,     5,    -5,   -16,   -14,    -7,    -1,    -1,     2,     0,     6,     5,    -1,    -2,    -8,    -7,    -2,     0,     0,     1,    -1,    -1,     4,     9,     1,     1,     2,    -1,     0,    -5,   -19,   -22,    -4,    -3,     0,    -1,     0,    -5,     2,     5,     3,     1,    -5,    -8,   -11,     1,    -5,     1,     0,     5,     0,     6,     0,    -1,    -1,     0,    -5,   -13,   -16,   -13,     0,    -2,     1,    -4,    -1,    -3,    -4,     5,     4,     2,    -4,    -7,    -7,     1,    -6,     2,     1,     5,    -7,     0,    -2,     0,     4,    -1,   -11,   -16,    -7,    -4,     0,     2,     1,    -7,     0,    -2,    -2,     6,     3,     1,    -6,    -6,     0,     1,     0,     0,     6,     1,    -8,    -2,     0,     4,     1,    -4,   -12,   -14,    -5,    -3,     6,     0,    -2,    -1,     3,    -3,     3,    -1,    -3,    -3,    -6,    -6,     1,    -1,     0,    -1,     1,    -1,    -3,    -1,    -2,    -2,    -4,    -5,    -9,    -6,    -1,     2,     0,     1,    -3,    -5,     2,    -2,     0,    -3,    -1,    -2,    -5,    -4,    -1,     0,     0,     1,     1,     0,    -6,    -7,    -5,    -8,   -11,    -6,    -5,     1,     2,    -1,     0,    -1,    -4,    -4,    -1,     2,     2,     0,     2,    -2,    -6,     8,     0,    -1,     1,     0,     0,    -1,    -8,    -4,    -4,    -6,    -8,    -5,     1,    -2,     0,     2,     3,    -1,     2,    -2,    -4,     2,    -4,     6,    -2,     0,    -6,     1,     1,    -1,     0,    -1,     0,    -2,    -6,     0,     1,    -7,    -3,    -1,    -4,     3,     1,     1,     0,     0,    -4,    -1,     1,    -2,     0,     3,    -5,    -1,    -6,     2,     0,    -1,     1,     0,     0,     0,     1,     3,     0,    -4,     0,    -1,     5,     0,     3,     2,    -6,     3,    -1,    -2,     0,    -4,    -7,     3,     1,    -2,    -7,     1,    -4,     1,     0,     0,     0,     0,     1,    -2,     2,     2,     2,    -1,     0,     3,     6,     4,     1,     7,     2,     4,     0,    -2,     2,    -2,     1,     0,    -7,     2,    -1,     1,    -1,     0,     1,     0,    -2,    -1,    -3,     1,    -4,     0,     0,    -5,     0,     7,     5,    -1,    -3,     0,     2,    -3,    -5,     0,     3,     2,     1,    -1,    -1,    -1,     1,    -1,    -1,     0,     0,     1,     3,    -1,     2,     5,     4,    -1,     0,     2,     4,    -2,    -3,     2,     5,    -6,    -1,     0,     7,     7,     7,    -1,     0,    -1,     1),
		    48 => (   -1,    -1,     0,     0,     0,     1,     1,    -1,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,     1,    -1,     0,    -1,     1,     0,    -1,     1,     0,     0,     1,     1,     1,     0,     0,     1,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -2,    -1,    -3,    -2,    -2,     0,     1,     0,    -1,    -1,     1,     0,     0,    -1,     1,     1,     0,     1,     0,     0,    -1,    -1,    -4,    -5,    -7,    -5,     1,     0,     1,    -3,    -3,     0,    -2,     1,    -5,    -4,    -4,    -2,    -3,    -1,     1,    -1,    -1,    -1,    -1,     0,    -2,    -4,    -5,    -5,    -3,    -4,    -4,     1,     4,     3,     1,    -3,     0,    -1,     4,     2,     1,    -1,    -1,     8,     1,     1,    -2,     1,     1,    -1,     1,    -3,    -5,    -8,    -5,    -6,    -3,     1,    -2,    -1,    -3,    -5,     0,    -4,    -1,    -2,    -3,     4,    10,    11,     3,    -7,    -8,    -3,     3,    -1,     0,     0,    -3,    -2,    -6,    -4,    -3,    -1,    -1,    -3,    -2,     1,     0,    -4,     0,   -10,    -7,    -5,    -7,     1,     6,     8,     4,    -3,    -5,    -2,     1,    -1,    -1,     0,    -2,    -8,    -1,    -3,    -1,     1,    -5,    -2,    -2,    -1,    -2,    -2,    -3,    -5,    -2,    -1,     1,    -2,    -2,    -1,    -1,    -3,    -6,    -4,     0,     1,     0,    -2,    -2,    -5,     0,     0,     0,    -1,     0,    -3,    -3,    -5,    -6,     0,     0,     2,     1,    -3,     0,     7,     1,     0,     2,    -2,    -6,    -3,     2,     3,     0,    -4,    -2,     2,     2,     2,     2,     0,    -1,    -4,    -5,    -8,    -7,    -6,    -2,     2,    -3,     3,    -1,    -3,     1,     7,     6,    -1,    -4,     1,     3,     6,     0,    -3,    -4,    -2,     2,     0,     2,     3,    -1,     1,    -1,    -5,    -7,   -11,    -5,    -3,    -3,    -1,     0,    -1,     1,     3,    -1,    -2,    -2,    -3,    -1,    -1,     1,    -3,    -5,    -5,     0,     3,     0,     0,    -3,     3,    -2,    -2,    -6,    -8,    -4,    -1,     3,     2,    -2,     4,     5,     0,    -1,    -2,    -2,    -6,     0,    -3,     0,     0,    -3,     4,    -3,     0,     2,    -2,     1,     3,     3,    -2,    -1,     0,    -2,    -8,    -2,     5,    -1,     1,     2,    -1,    -5,    -4,    -6,    -4,    -1,    -2,     0,     1,    -3,    -3,    -2,    -1,    -3,    -3,    -6,    -2,     2,     6,     1,    -4,    -6,    -6,    -1,     3,    -3,    -2,     1,     0,    -3,     0,     1,    -2,    -3,    -3,     0,     0,    -4,    -4,    -6,    -2,    -2,    -1,     0,     3,     1,     6,     3,     2,    -6,    -5,     1,    -2,    -9,    -3,    -3,    -2,     0,    -1,    -5,    -4,     1,    -1,    -1,    -1,    -2,    -5,    -4,    -5,    -8,    -6,     2,    -4,    -1,     2,     1,     3,    -2,    -4,     1,    -5,    -6,    -7,    -6,    -2,    -5,    -3,    -6,    -2,    -8,    -3,    -1,     0,    -2,     2,     0,     0,    -7,    -6,    -5,    -4,    -8,    -1,    -2,     4,     3,     3,     2,     0,    -7,    -8,    -6,    -1,    -4,    -3,    -2,    -1,    -6,    -5,    -1,    -2,    -2,     3,    -1,    -3,    -4,    -5,    -1,    -5,    -3,    -1,    -3,     2,    -4,    -2,    -1,     0,    -6,    -3,    -4,     2,    -4,    -4,    -3,    -3,    -6,    -5,    -1,    -2,    -4,     3,    -1,    -4,    -6,    -5,   -10,   -10,    -2,     0,     3,     4,    -4,    -3,    -6,     0,     0,    -4,     3,     3,     6,    -1,    -4,    -1,    -1,    -3,    -2,    -1,    -2,    -1,    -2,    -3,    -7,    -7,    -7,    -4,    -1,     2,     7,    -2,     0,     3,    -2,     4,     1,     1,    -1,     0,     2,    -2,    -3,    -2,    -2,    -2,     1,     1,    -1,    -2,    -1,    -3,    -7,    -5,    -5,    -2,    -2,     0,     6,    -4,    -1,     3,    -5,     5,     5,     1,    -2,    -2,     1,     2,    -4,    -2,    -5,    -2,     1,     1,    -2,    -1,    -4,    -3,    -8,    -7,    -4,     0,     4,     5,     4,    -3,    -3,     1,    -8,     6,    -3,     4,     1,     0,    -1,     1,    -2,    -2,    -6,     0,    -2,    -1,    -1,    -1,    -4,    -5,    -9,    -8,    -4,    -2,     3,     4,     1,    -5,    -2,    -1,     0,     0,     0,     3,    -1,     1,     2,     1,    -7,    -1,    -5,     1,    -1,     0,    -2,    -1,    -2,    -5,   -12,    -9,    -9,    -6,     0,     1,    -2,     2,    -3,     1,    -2,    -6,    -2,    -1,     1,     5,     1,    -5,    -4,     0,    -3,    -1,     1,     1,    -3,    -3,    -1,    -3,    -5,    -4,    -7,    -5,    -1,    -5,     0,    -1,     0,     1,    -1,     2,    -3,    -1,     6,     2,     5,    -1,     1,    -1,    -3,     0,     0,     0,    -1,     0,    -1,    -3,    -7,    -7,    -7,    -3,    -1,    -3,    -5,    -7,    -5,    -3,     5,    -4,     1,     1,     7,    -1,    -3,    -2,    -4,    -2,    -1,    -1,    -1,     0,    -3,    -1,    -3,    -4,    -3,    -7,    -6,    -6,    -4,    -5,    -4,    -5,    -1,     6,     7,     4,     4,     2,     2,    -3,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,     0,    -4,     0,    -2,    -4,    -2,    -1,    -4,    -7,    -4,    -4,    -5,    -9,    -7,    -5,    -2,    -1,    -8,    -9,    -3,    -4,    -1,    -1,     0,     1,    -1,    -1,    -1,     1,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -2,     1,     0,    -3,    -2,    -4,    -4,     0,     0,     0,    -1,     0,    -1,     1,     1,     1,     0),
		    49 => (   -1,    -1,     0,     0,     0,     0,     1,    -1,     0,     1,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     1,    -1,     0,     1,    -1,     1,     0,     1,     1,     0,     0,     1,     0,     0,     1,     0,    -1,    -1,    -2,    -3,    -3,    -3,     0,    -9,    -8,    -7,    -3,    -1,     1,    -2,     0,    -1,     1,     0,    -1,    -1,    -1,     1,    -1,    -2,    -2,     0,    -1,    -4,    -4,    -2,    -2,    -6,    -3,    -3,    -7,    -3,    -6,    -2,     0,    -2,    -5,    -1,    -1,    -3,    -1,     1,     0,     0,    -1,     1,    -1,   -10,    -3,    -3,    -1,    -5,    -6,    -8,    -7,    -7,   -14,   -10,   -12,   -11,   -11,    -5,     1,    -5,    -6,    -4,    -2,    -1,    -2,    -2,    -1,     1,     0,     1,    -3,    -3,    -3,    -7,   -10,    -7,    -6,   -10,    -7,   -14,   -16,    -4,    -9,    -6,    -4,     1,     3,   -17,    -9,   -11,    -6,    -2,    -1,    -7,    -6,    -2,    -1,     1,    -2,    -3,    -1,    -4,    -8,    -6,    -7,    -7,    -4,     1,    -2,     4,    -4,    -2,    -6,    -5,    -5,    -5,    -3,    -3,   -11,    -9,    -6,    -5,    -5,     0,    -1,    -2,    -2,    -9,   -11,   -22,   -11,    -1,     0,     9,     2,     4,    -1,     7,    -1,     1,     2,     3,     4,     0,     3,     2,    -7,    -7,   -10,   -10,    -6,    -4,     1,    -6,    -8,   -10,   -17,   -21,    -1,    -7,    -3,     1,     3,     4,     7,     2,    -2,     5,    -1,     3,     2,     0,    -1,     0,    -4,   -10,   -10,    -8,    -6,    -2,    -9,    -7,    -6,    -6,   -11,     0,    -1,    -6,     1,    -3,    -2,     0,     0,    -4,     0,    -3,     0,    -1,     3,    -3,     0,     3,    -4,    -4,    -6,    -9,    -9,    -4,    -2,    -4,    -1,    -3,   -10,    -1,    -1,     0,    -3,    -4,     0,     2,     0,    -2,    -3,     6,    -2,    -3,    -3,     1,     0,     3,     0,    -2,    -3,    -9,    -9,    -3,    -1,    -7,   -10,    -1,     2,     1,    -4,    -4,    -2,     2,    -2,     2,     2,    -4,    -5,    -5,    -2,     3,    -2,     2,     4,     1,     3,    -2,    -5,    12,    -9,    -6,     1,   -15,     5,    -2,     5,    -2,    -3,    -2,     3,    -1,     6,     1,     1,     1,    -4,    -2,     1,     6,     2,     2,     4,     4,     9,    -4,     1,    12,    -7,    -7,    -1,    -4,     3,     3,     9,     2,     1,     3,     1,     6,     0,     3,    -7,    -8,     1,     0,     2,     6,     8,     8,     3,     6,     6,     9,   -10,   -19,   -11,    -2,     1,    -7,    -6,     1,    12,     9,     3,     7,     7,     4,     5,     0,     2,     2,     4,     3,     7,     0,     3,     5,     7,     5,    14,     3,   -16,   -10,    -7,     0,    -3,    -6,    -3,     2,     9,     8,     2,     3,     8,     2,     5,    -3,    -3,     2,    -2,     0,     5,     1,     4,     6,    -1,     3,    15,    -1,   -22,   -15,    -1,    -1,    -1,    -1,   -12,     3,     9,     1,    -4,     4,    10,     5,     1,    -5,    -4,     2,    -3,     5,     5,     8,     6,     5,    -3,    -5,    -1,    -5,   -20,   -11,     5,    -2,     1,    -1,   -11,    -7,     2,    -6,    -1,    -1,    -1,    -5,     6,    -5,    -3,    -3,    -3,     0,    -1,     1,    -1,    -3,    -2,    -9,    -3,    -5,   -17,    -9,    -2,    -6,     1,     0,   -13,     0,    -4,    -5,    -5,     1,    -1,    -3,    -3,    -8,    -2,    -4,    -4,     2,     1,     2,    -4,    -5,    -5,    -5,    -5,    -4,   -13,    -1,    -2,    -4,     5,     0,   -12,     1,    -5,    -7,    -3,    -1,     1,    -1,     1,    -2,    -4,    -8,     0,    -2,    -1,     0,     2,    -1,    -6,     1,    -1,   -11,   -23,    -2,    -6,    -4,     1,    -1,    -6,     8,    -4,    -9,    -7,    -8,    -5,    -6,    -6,    -4,    -7,   -14,    -2,    -1,    -4,    -3,    -2,     3,    -1,    -4,     4,    -5,   -10,    -1,    -5,    -2,     1,     0,   -11,     6,    -3,     7,    -4,   -17,   -13,    -8,   -10,    -2,    -8,    -9,     2,    -3,     1,     1,    -4,     2,    -7,    -5,    -3,    -2,     1,     4,    -3,    -1,    -1,     0,   -11,     8,     2,     7,    -4,    -7,    -7,    -7,   -10,    -8,    -8,     0,   -10,    -4,     1,    -4,    -6,    -4,    -8,    -2,    -4,    -8,    -4,     3,   -19,    -1,     1,    -1,   -10,     7,    -6,    -3,     2,     5,     5,     0,     2,    -4,    -2,     0,     0,     2,    -3,    -4,    -6,    -9,    -3,    -1,    -1,    -9,     1,    -3,   -12,    -2,     0,     0,    -8,     6,    -2,    -4,    -3,     1,     0,    -4,     0,    -5,    -4,     0,     0,    -6,    -5,    -3,    -3,    -2,    -1,     4,     4,    -2,     0,     0,    -2,     1,     0,     1,    -8,    -8,    -1,     4,    -5,     3,    -2,    -1,     2,     4,    -2,    -3,    -8,    -1,     1,    -5,     1,     2,    -4,     1,     6,     7,     0,    -3,    -4,     0,    -1,     1,     6,    -5,     7,     3,    -9,   -11,    -4,    -2,    -7,    -6,     2,    -1,     8,     0,     3,     6,     6,     4,     8,    10,     2,    -2,    -3,     0,    -5,     1,     0,     0,     0,     4,     5,     0,     2,     0,     2,     2,    -5,    -1,     6,     2,     8,     2,     3,     9,    11,     3,     8,     8,     4,     5,     5,     1,     1,    -1,    -1,     0,     0,     0,    -6,    -7,     3,     2,     4,     2,    -1,     2,     1,    -4,     5,     4,     3,   -10,    -3,     5,     1,    -6,     2,    -6,     1,    -1,     0,     0),
		    50 => (    0,    -1,     1,     1,     1,     0,     0,     0,     1,     1,     0,     1,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,    -1,     1,     1,     0,    -1,     0,    -1,     1,     1,     1,     1,     1,     1,     1,    -1,     0,     0,     1,     1,    -1,     1,    -1,    -1,     0,     1,    -1,    -1,     1,    -1,    -1,     0,     1,     0,     0,     0,     0,     2,     3,    -2,    -2,    -1,    -2,    -3,    -4,    -7,    -8,    -8,    -4,    -6,    -5,    -5,    -2,     1,     1,     0,    -5,    -1,     0,     0,    -1,     0,     1,    -1,     0,     1,     0,     2,    -3,    -2,    -8,    -8,    -3,     0,     0,     3,     0,    -7,    -8,    -4,    -2,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     1,    -1,    -1,     0,     1,    -2,    -7,     4,    -1,     5,     5,     3,     4,    -2,    -1,    -1,    -5,    -1,     2,     3,     1,    -6,    -8,    -2,     0,    -1,    -1,    -2,     0,     0,     1,     0,     2,     1,    -4,     0,    -2,    -7,    -1,     2,     3,     1,     3,     2,    -1,     3,     1,     2,    -1,    -2,    -2,     0,    -1,    -4,    -5,    -4,    -5,     0,     1,    -3,    -2,     3,    -2,     0,    -3,    -3,    -1,     1,     2,     0,     0,     1,     1,     5,     2,     3,    -2,    -1,    -5,    -2,     8,     5,    -6,    -7,    -1,     1,    -2,    -3,    -2,    -3,     4,     3,     2,    -1,     3,     5,     1,     1,     0,     2,     0,     0,     3,     0,    -2,    -6,    -5,    -3,     3,     4,    -5,    -5,     2,     2,     0,     1,    -3,    -3,     0,    -1,     0,     5,     5,    -1,    -1,     7,     3,     4,    -2,     1,    -3,     0,    -3,    -1,    -2,     2,     0,     1,    -5,    -7,    -3,    -1,     0,     0,    -2,    -6,     5,    -5,     0,    -1,     2,     0,     0,    -2,    -1,     1,     1,    -4,    -5,     6,     6,     6,     3,     4,     0,     7,    -8,    -7,    -1,     1,    -1,     0,    -2,    -8,     1,     0,    -1,     2,     1,     4,    -1,    -7,    -3,    -1,    -1,    -4,     3,     4,    -2,    -5,    -3,     7,     2,     6,    -5,    -4,    -1,     0,     3,    -4,    -4,    -6,    -1,     1,    -1,     1,     1,     3,    -7,    -7,    -7,    -6,    -7,    -2,    -1,     0,    -5,    -4,    -5,    -3,     1,     4,    -3,    -1,    -1,     1,     1,     0,    -3,     0,    -5,     2,    -2,     0,    -1,    -5,    -2,    -5,    -5,    -5,    -6,    -4,    -2,    -5,     1,    -1,    -3,    -1,    -7,     1,    -2,    -5,    -2,     0,     3,     1,     1,     6,    -1,     0,     0,     6,     2,    -4,   -11,   -10,   -15,   -12,    -8,    -6,    -5,    -1,    -4,     0,    -1,     1,    -5,     0,    -1,    -2,    -2,    -1,     0,    -1,    -3,    -3,     7,     3,     5,     2,     2,    -4,   -14,   -10,   -12,    -5,    -7,   -10,    -8,    -2,     1,    -3,     1,    -3,     3,     6,     0,    -5,     0,     1,     1,     0,    -8,     2,     6,     7,    -2,     1,     4,     3,    -9,   -16,   -10,    -3,    -4,    -6,    -6,    -4,    -1,    -1,     2,     1,    -2,     2,     0,    -1,    -4,     1,     0,    -1,   -10,     5,     6,     1,     8,    -4,    -1,     1,    -5,    -4,    -8,     0,    -5,   -12,   -10,    -8,    -7,     2,     6,     1,     0,    -1,    -3,    -3,    -1,    -1,     0,    -2,    -2,     3,     5,     3,     1,    -2,    -3,     3,     6,     3,     2,    -3,   -13,   -16,    -9,   -11,    -6,    -2,    -1,    -2,     1,    -4,    -4,    -7,     1,     0,     0,    -1,     3,    -4,     5,     7,     5,     1,     2,    -2,    -2,     0,    -5,    -7,   -10,   -13,    -6,    -2,    -1,     6,     3,     3,     2,     1,    -3,    -5,    -2,     0,     0,     1,     1,     0,     4,    -1,     1,     1,    -2,    -2,    -1,     3,    -2,    -2,    -5,     0,     4,    -5,     0,     3,     5,     5,     0,     1,    -3,    -1,    -2,     0,     1,    -1,     1,     7,     8,    -3,     0,    -3,    -6,    -5,     1,     2,    -1,    -1,     0,     2,     2,     1,    -1,     2,     3,    -3,    -1,     1,    -4,    -1,    -1,     1,    -2,     0,     6,     9,     2,     5,     1,    -5,    -2,    -4,    -1,    -4,    -2,     4,     4,    -3,     0,     0,    -1,     0,     4,     5,    -1,    -2,    -1,     0,     3,     0,     0,    -1,    -1,     1,     4,     4,     7,     5,    -1,     1,    -2,    -1,     0,     2,     2,     2,     2,     0,    -2,     1,    -1,     2,     1,    -4,     0,     0,     2,     0,    -1,    -1,    -6,    -6,     1,    -3,    -4,     0,     0,     2,     1,     4,     0,    -2,     3,     0,     5,     1,     0,    -5,    -5,    -2,    -2,    -9,     0,    -2,     0,     1,    -1,     0,    -2,    -3,     0,     3,     2,    -1,     5,     6,     1,     2,     4,    -4,     2,    -1,     5,     3,     5,    -5,    -6,    -6,    -3,     2,     2,     0,    -1,    -1,    -1,     0,    -1,     0,    -2,    -1,    -1,    -2,     0,    -2,    -6,    -4,    -4,    -6,   -10,   -11,   -11,   -14,    -9,    -7,    -9,    -5,    -1,    -3,    -1,     1,     1,     1,    -1,    -1,    -1,    -1,    -2,    -3,    -2,     1,    -3,    -2,    -3,    -1,    -7,    -6,   -10,    -7,    -6,    -8,    -9,    -7,    -8,    -5,    -5,     1,    -1,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,     1,    -1,     0,    -1,     0,    -2,     1,     0,    -1,     0,    -2,    -1,    -1,    -1,    -5,    -4,    -6,    -1,     1,     1,    -1),
		    51 => (   -1,    -1,     0,    -1,     0,     1,     1,     0,     0,     1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     1,    -1,     1,    -1,    -1,     0,    -1,     0,     1,    -1,    -1,     0,     1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     2,     1,    -1,    -1,    -2,     1,     0,     0,     1,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -4,    -7,    -7,    -5,     1,    -5,    -2,     7,     2,    -7,    -7,    -2,    -4,    -4,    -2,    -1,     1,     0,    -1,     0,     0,    11,     6,     0,    -5,    -3,    -1,    -3,    -4,    -7,   -10,    -5,    -1,    -4,    -6,    -2,    -3,    -1,     9,     7,    -7,    -1,    -4,    -1,    -1,     1,    -1,     0,     0,    10,    10,    -1,    -5,    -3,    -2,    -3,    -7,    -9,    -3,    -1,     5,     5,     0,    -6,    -9,     5,     2,     3,    -3,    -1,    -2,     0,    -1,    -4,    -4,    -1,     0,    10,     5,     2,    -1,     0,    -4,   -11,   -12,    -3,     1,    -3,     2,     1,     1,     3,    -7,    -4,    -2,    -6,    -4,    -2,    -1,    -1,    -1,    -4,    -4,     0,     0,    -4,     1,     0,    -2,    -4,    -1,   -10,   -13,    -7,     0,     2,     6,     2,    -4,     1,    -8,    -2,    -8,    -7,    -2,    -1,     1,     0,     0,    -3,    -3,     0,    -1,    -4,     1,    -1,    -6,    -7,    -2,   -15,    -9,     0,     2,     4,     7,     2,    -2,    -5,    -6,    -3,   -14,    -6,    -3,     0,    -1,     0,    -2,    -8,    -4,     1,    -2,    -4,     2,    -2,    -4,    -6,    -5,   -14,    -7,     1,     0,     1,     5,     8,     5,    -6,    -5,    -4,   -14,    -4,    -3,     3,     0,    -1,    -1,    -5,    -2,     1,    -2,    -5,    -2,    -2,     0,    -3,    -3,    -7,     0,     3,    -1,    -7,     0,     9,     7,    -5,   -10,     0,     1,    -5,    -1,     2,    -1,    -4,    -2,    -4,    -7,     0,    -2,    -2,    -2,    -4,    -1,    -7,    -3,    -3,    -7,     6,    -1,    -3,     3,     5,    -1,    -3,    -8,    -6,     0,    -2,   -10,     1,     4,    -6,    -3,     1,     6,     0,     1,    -1,    -2,    -2,    -4,    -9,    -5,    -8,    -5,    -1,     3,    -3,     1,     7,    -2,     0,    -5,    -7,    -3,     4,    -1,     3,     4,    -5,    -3,    -3,    10,     1,     0,    -9,     4,     0,     0,    -3,    -3,    -2,     6,     2,    -1,     2,     1,     4,    -3,    -1,    -8,    -9,    -5,     8,     1,     1,     5,    -5,     1,     1,     8,     1,    -1,    -9,     1,     1,    -1,    -1,     2,     6,     4,    -9,     2,     2,    -4,    -3,    -3,    -1,    -5,    -6,     2,     9,    -3,    -4,    -7,    -6,     5,     4,    -1,     0,     0,    -1,     1,    -1,    -5,     0,     3,    -2,    -3,    -8,    -6,     2,    -1,    -1,    -4,     1,     0,     0,     1,     2,    -4,    -7,    -1,    -1,    -2,     6,     1,    -1,     0,     1,     3,     0,    -6,    -5,     0,    -2,    -4,    -3,     8,     4,     6,     2,    -6,     0,    -1,     4,    -2,     5,    -2,    -6,    -2,    -6,    -4,     1,    -3,     0,    -1,     1,    -4,     0,    -3,    -2,     0,    -2,    -5,    -3,     4,     2,     0,     2,    -5,    -5,    -1,     2,    -5,     1,    -3,    -4,    -5,     0,    -5,     0,    -2,    -1,     1,     0,    -2,    -1,    -6,    -4,    -6,    -2,    -4,    -4,    -2,     1,     1,     1,    -3,    -4,    -5,     1,    -5,    -6,    -4,     3,     3,    -3,    -5,    -1,     1,    -1,     0,    -1,    -1,    -3,     0,    -4,    -2,    -6,    -4,   -13,    -3,    -4,     7,     4,    -1,     1,    -2,     3,    -8,     2,    -1,    -7,    -6,    -6,     0,     0,     5,    -1,    -1,     1,    -1,    -1,    -1,    -1,    -4,     2,    -7,    -7,    -2,    -1,     3,     6,     3,     0,    -5,    -3,   -11,    -3,    -3,    -9,    -6,    -2,     3,     4,     6,     1,     1,     0,    -3,    -3,    -2,    -4,    -8,    -2,    -3,    -2,    -1,     5,     2,     3,     2,     1,    -2,    -3,    -5,     0,    -8,   -12,    -4,     0,    -1,     6,    -1,     2,     2,     1,    -3,    -3,    -1,    -5,   -11,    -1,     0,    -3,     0,     0,     1,    -1,     0,    -2,    -7,     5,    -2,     2,    -3,    -9,    -8,    -3,     2,    -2,     0,     3,     1,     1,     1,    -2,    -1,    -2,    -9,     1,    -1,    -2,    -4,    -3,    -1,     1,    -2,    -2,    -3,     3,     1,     5,    -1,    -7,    -3,    -6,     5,     4,     0,     1,     0,    -1,    -3,    -1,     1,     5,    -3,     1,     7,     1,     4,    -1,     0,     0,     0,     2,     7,     6,     2,     4,    -3,    -1,    -4,    -4,    -1,     9,     1,    -1,    -1,    -1,    -2,    -1,    -1,     6,     1,    -1,     1,     5,     7,    -1,    -6,    -6,    -8,   -11,    -4,    -8,    -5,    -5,    -3,    -8,    -1,    -4,     6,     5,     1,     1,     0,    -1,     0,    -1,    -1,     0,    -1,    -2,    -4,   -16,   -13,    -9,    -8,    -2,   -10,    -9,   -11,    -9,    -9,   -15,    -6,    -4,    -4,     0,    -1,    -1,     1,     1,    -1,     0,     0,    -4,    -7,    -5,    -5,    -5,    -4,    -3,    -4,    -8,    -8,    -8,    -8,    -6,    -6,    -2,    -3,    -1,    -4,     0,     0,    -1,     1,     0,     0,    -1,     0,     1,     0,    -1,     1,     0,     0,    -1,     1,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1),
		    52 => (    0,     1,    -1,    -1,     1,     0,    -1,     1,    -1,     0,     1,     1,    -2,    -1,     1,     2,     0,     1,     1,     0,     0,    -1,     1,    -1,     0,     1,     0,     0,     0,     0,     1,    -1,     1,     1,    -1,    -1,    -1,     1,     1,    -1,     1,     1,    -2,    -2,     1,     2,    -1,    -5,    -3,     0,     0,     1,     1,     1,     0,     1,    -1,     0,    -2,    -2,    -2,     1,    -1,    -2,     5,     7,     9,     4,     4,    -3,     0,    -3,    -9,    -7,     0,     2,     0,     2,    -3,     2,     4,     2,    -1,     0,    -1,    -1,    -2,    -8,    -6,    -7,    -2,    -4,     2,     3,    -1,    -1,    -3,     2,     3,    -2,     0,    -1,    -2,     6,    -2,    -1,    -2,    -9,    -5,     2,    -2,     0,     0,    -1,    -1,    -2,     6,    -1,    -1,     1,     0,     1,    -2,     0,     4,     1,     0,     2,    -4,     2,    -5,    -2,     3,    -5,    -2,    -8,    -9,     4,    -7,    -3,    -1,    -1,     0,    -3,     1,    -7,    -8,   -11,    -5,    -1,     5,     1,    -4,     3,     2,     1,    -3,     2,    -1,     0,     0,     2,     0,     4,    -7,     7,    -5,    -1,    -1,     0,     0,     7,     6,    -6,    -5,    -3,     2,     5,     5,     0,     1,     6,     1,     0,    -2,     1,     0,    -1,    -2,    -5,    -2,    -1,     1,    -6,    -6,    -1,     0,     0,    -2,    10,     7,     5,    -2,     1,    -2,     0,    -1,     2,     2,     3,     1,     4,     5,     4,     1,     4,    -2,    -4,     6,     1,    -5,    -6,    -5,    -4,    -4,     7,    -1,     7,     5,     4,    -5,    -2,    -2,     4,     0,    -1,    -2,    -4,    -1,     1,     4,     5,    -1,     6,    -4,     0,     6,     5,   -14,    -9,    -6,    -4,     1,    -2,     2,     1,    -2,     1,    -3,    -4,    -2,     5,    -5,     1,     3,    -7,    -2,     1,     3,     2,    -1,     6,     0,    -3,    -4,     5,   -11,    -7,    -3,    -2,     0,     0,     1,     4,    -8,     9,     4,    -1,    -2,     0,    -5,    -6,     0,     3,    -2,    -2,    -2,    -3,    -1,     1,     3,    -1,    -3,     5,    -2,    -3,     1,    -1,     0,    -4,    -1,     5,     1,     2,     4,     0,    -2,    -5,   -11,     0,    -4,    -6,    -7,    -6,     0,    -2,    -6,    -1,    -3,     0,    -3,     3,    -1,     0,    -6,    -1,    -1,     0,    -7,    -1,     2,    -8,    -3,    -6,    -7,    -5,    -6,    -6,    -2,   -10,   -12,    -3,     0,    -1,    -7,    -1,    -4,    -2,    -1,    -4,    -2,     3,     0,    -3,     0,     1,     0,    -1,    -1,    -3,   -11,    -9,   -16,    -9,    -7,    -9,   -12,    -7,    -5,    -3,    -2,    -5,    -4,    -6,    -5,    -5,     2,    -4,    -1,     3,     5,    -3,     1,    -4,    -5,    -2,    -6,   -11,   -12,   -13,   -20,   -13,    -6,    -7,    -2,    -4,     0,    -3,    -7,    -3,    -2,    -2,    -6,    -9,    -1,   -10,    -1,     0,     7,     3,     1,    -3,    -1,    -3,   -12,    -6,    -6,    -8,     2,    -1,    -3,     3,     0,     4,     1,    -6,     1,    -1,    -7,    -9,    -8,    -5,    -9,    -5,     2,    -3,     7,    11,     0,     0,    -5,    -8,   -14,    -5,    -5,    -4,    -2,     2,     2,     3,    -4,     2,     2,    -3,    -4,    -2,    -4,    -8,    -5,    -2,     4,    -3,     3,     7,    10,     6,    -1,    -1,     0,    -5,    -5,    -6,    -1,    -2,     0,     1,     3,     1,    -4,     7,     5,     0,    -1,    -2,    -1,    -7,    -4,    -2,    -2,    -2,    -5,    12,     7,     6,    -1,    -1,    -2,   -10,    -4,    -3,     3,     5,    -2,    -3,     1,     0,     2,    -1,    -1,    -2,    -1,     3,    -4,    -5,    -6,     4,     5,     5,     9,    15,    -1,     8,    -1,    -2,     2,    -5,    -6,    -2,     5,     3,    -3,    -5,     2,     1,     0,     9,     8,     2,     4,    -1,    -2,    -4,     1,     5,     2,     5,    -1,     4,     4,     8,     0,    -1,     5,    -1,    -1,    -3,    11,     4,     3,     4,     8,     7,     5,    13,     4,     4,     7,    -1,    -1,    -1,     8,     7,     3,     2,     2,     6,     3,     0,     1,     2,     2,     6,     2,     2,     6,     4,    -1,     3,     3,     3,     0,    10,     8,     6,     4,     5,     2,     4,     4,     3,     6,    13,     6,     6,     6,    -2,     1,     0,     0,     0,    -1,     6,     9,     5,     1,     5,     1,     2,     1,     1,     3,     2,    -2,    -6,     0,    -5,     2,     5,     9,    11,     9,    -1,    -8,    -3,    -1,    -1,     1,    -6,    -3,     2,     6,     3,     3,     6,     2,     8,     6,     4,     2,    -2,    -5,    -3,    -4,     0,     5,     6,    12,     8,     7,     1,    -4,     0,     1,     0,    -6,    -4,    -1,    -4,     0,     3,     9,    -3,     1,     1,     6,    -3,     4,     2,    -6,    -2,     0,     0,    -7,    -4,    -1,     7,    13,     7,     4,     0,     1,     0,    -4,    -1,    -5,   -13,     6,    -2,    -7,   -13,   -17,    -5,    -3,    -1,     6,     4,    -4,     2,    -9,   -11,    -1,     2,    -9,    -4,     2,     7,     5,     0,     1,    -1,    -1,     0,    -4,    -8,    -9,    -6,    -5,    -8,   -14,   -12,    -7,    -7,    -7,    -5,   -11,   -10,    -8,    -1,    -4,    -5,    -3,     0,    -1,     0,    -1,     1,    -1,     1,    -1,     1,    -1,     0,    -2,     0,     1,     0,    -4,    -6,     0,    -3,    -1,     0,     0,    -1,    -1,     0,    -2,    -4,    -2,     0,    -1,     0,     0,     0),
		    53 => (    0,    -1,     0,    -1,     0,    -1,     1,    -1,     1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     1,    -1,    -1,     0,     1,     0,     0,     0,    -1,     0,     1,     0,    -1,     0,     1,    -1,     1,    -1,     0,     0,    -1,    -1,    -2,    -1,    -3,    -1,     0,    -1,     0,     0,     1,     0,     1,     1,     0,    -1,     1,     1,     0,    -1,     0,     1,     1,     0,    -5,    -6,     4,     5,     3,    -2,    -5,    -5,    -7,    -7,    -5,    -3,    -1,    -3,    -4,    -6,    -2,    -1,     0,     0,    -1,     0,     0,    -3,    -1,     0,    -2,     2,     1,    -1,     4,     4,     3,     3,     1,    -3,     2,     4,     5,    -2,    -2,    -3,    -1,    -9,    -4,    -1,     0,     0,    -1,     2,     1,     0,    -2,     1,     1,     3,     2,    -1,    -2,    -4,    -6,    -6,     0,    -3,    -3,    -8,    -3,     0,    -5,    -4,     5,   -10,    -8,    -4,    -1,     0,     0,     1,     1,    -2,    -1,     4,     5,     8,     1,    -6,    -8,    -4,    -3,    -3,     0,    -1,    -1,    -1,    -1,     1,    -1,    -3,    -5,    -4,    -4,    -1,    -4,    -1,     0,     2,     0,     2,     1,     0,     1,    -1,    -7,    -5,     4,    -1,     1,    -2,    -4,    -2,    -1,     0,     0,    -5,    -4,    -2,    -2,    -1,    -1,    -8,    -5,    -2,     1,     2,     3,    -5,   -11,    -5,     0,    -4,    -6,    -2,    -2,     1,    -2,     0,     1,     1,    -1,     3,     0,    -5,     1,    -3,    -1,    -4,    -3,    -6,    -5,    -2,     0,    -1,     3,    -7,    -9,     0,    -3,    -5,    -3,     2,     2,    -1,     0,    -4,     1,    -3,     1,     0,     4,     1,     2,     7,     4,    -9,   -15,    -5,    -6,     0,    -1,    -6,    -5,    -5,     1,     0,     3,    -1,    -2,    -2,     3,     5,     7,     4,     3,    -2,    -3,    -2,    -4,    -2,     4,     3,     3,    -7,   -18,    -7,    -7,    -1,     0,    -6,    -3,     4,     2,     2,     7,     1,    10,     5,     5,     4,     0,     0,    -1,    -3,    -9,    -1,     4,     4,     3,    -1,     3,    -2,   -16,    -2,    -5,     1,    -1,    -6,    -3,     9,     8,     8,     2,     5,     3,     7,     3,    -5,   -10,   -10,    -8,     3,     2,     3,     4,     5,     8,     2,     2,     0,   -10,    -9,    -2,    -1,    -1,    -6,    -6,     9,     5,     4,     0,     2,    -6,    -6,    -8,   -18,   -13,    -3,     4,     8,     3,     1,     4,     0,    -2,    -4,    -3,    -6,     0,     1,     0,     1,     1,    -4,   -12,     4,    -6,    -4,    -3,    -4,    -8,   -17,   -17,   -11,    -2,     3,     6,     1,     1,    -1,    -4,    -5,    -3,    -2,    -9,    -7,     5,    -3,    -3,    -1,    -2,     2,    -2,    -3,    -8,   -10,   -14,   -13,   -12,    -6,    -3,    -5,     3,     4,     2,     2,    -1,     1,    -6,    -4,    -5,    -4,    -9,    -2,     8,    -2,    -4,    -3,    -1,     4,     2,     1,    -3,    -5,   -11,   -14,   -10,     0,     3,    -2,     3,     7,    11,     0,     4,    -1,    -2,     0,    -2,     0,    -5,    -3,     6,    -2,     5,     1,     0,     1,     3,     6,     1,    -4,    -6,    -4,    -8,    -6,    -6,   -11,    -1,     1,    -2,    -5,     4,     3,    -3,     1,     1,     7,    -2,    -5,     3,    -6,     2,     0,     0,     1,     1,     1,     0,    -1,    -2,    -5,   -11,   -14,   -17,   -19,   -23,   -19,   -12,    -7,     5,    -1,    -6,     4,     4,     7,     2,    -5,    -2,    -9,    -1,     0,    -2,     1,     7,     2,     9,     1,    -4,     0,    -2,    -9,    -8,   -12,   -18,   -14,    -8,    -8,    -1,     6,     4,     4,     1,    -1,     3,    -2,   -11,    -3,     1,    -3,     0,    -4,    -4,    -4,     2,     4,     0,     0,    -3,     2,    -1,    -4,    -3,     0,     0,    -2,    -2,     0,    -3,     0,     1,     0,     5,     0,    -3,     2,    -2,    -3,     1,    -1,    -4,    -1,     2,     4,     5,     3,     1,     6,     5,     7,     3,     0,    -2,    -7,    -3,    -5,    -4,     1,     5,    -1,     2,    -4,    -5,    -4,    -1,    -1,    -1,     3,    -2,     0,    -2,     3,     1,     5,     6,     2,     0,     0,     1,    -2,     0,    -5,    -5,    -7,    -2,     2,     3,     0,    -3,    -4,    -6,    -3,    -2,     0,    -1,     1,    -3,     1,     1,    -2,    -3,    -4,    -1,    -1,     1,     1,     2,     2,     2,    -1,    -1,     0,    -1,     4,     0,     1,    -7,    -6,    -5,    -3,    -2,     1,     0,     1,     3,     5,     6,     4,    -1,    -2,    -2,    -1,    -6,    -3,    -5,    -2,    -2,     4,     1,     3,     4,     0,     2,     3,    -7,    -5,     5,     3,     0,     0,    -1,    -1,     0,     4,     5,     0,    -4,    -2,     1,     3,     0,     1,     3,     1,     1,    -2,     5,     4,    -3,    -7,    -2,    -2,    -5,    -8,    -5,    -3,    -1,     0,     0,     1,     0,    -5,    -4,     2,     3,     2,    -3,    -3,    -9,    -8,    -6,   -11,    -8,     0,     0,    -6,    -6,    -6,    -3,    -4,    -4,    -7,     0,     0,     1,     0,    -1,     0,     0,    -4,    -9,    -9,    -6,    -7,    -9,    -8,   -12,   -10,    -9,    -4,    -3,    -4,    -5,   -12,   -11,   -10,    -1,    -4,    -1,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -6,    -5,    -6,     0,    -4,    -4,    -5,    -4,    -4,    -4,    -6,    -2,    -1,    -1,     0,    -1,     0,     1,     0),
		    54 => (   -1,    -1,    -1,     1,     0,    -1,     1,     0,     0,    -1,     0,     0,    -2,    -2,    -2,    -1,     1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,     1,     1,     0,     1,     1,     1,     1,    -1,    -5,    -4,    -1,     0,    -2,     0,    -2,     2,     5,    -1,    -1,    -1,    -1,    -1,    -3,    -2,    -2,    -1,    -1,     1,     0,     0,    -1,     0,    -1,    -2,    -7,    -1,    -3,    -5,    -8,    -3,    -2,    -1,    -2,    -5,    -4,    -7,    -9,    -4,    -2,    -1,    -6,    -5,     0,    -2,    -1,    -4,     0,     0,     0,     0,    -2,    -3,    -6,    -2,    -4,    -6,    -2,    -1,    -3,    -2,     1,    -3,    -5,    -1,     1,     4,    -5,    -3,    -5,    -2,    -3,     0,    -1,    -2,     1,     0,     1,     0,    -2,    -1,    -2,    -4,    -6,     3,     7,     4,    -3,    -9,   -12,    -7,    -6,    -6,   -10,   -12,   -13,    -8,    -4,    -3,     1,    11,     8,     5,    -9,    -2,    -1,    -1,    -3,     1,    -3,     0,    -3,     3,    11,     3,    -7,   -12,    -8,    -5,    12,     7,     5,    -2,   -12,   -15,    -5,    -5,    -1,     3,     2,    -3,    -1,    -1,     0,     1,    -1,    -4,     4,     6,    -2,     4,     5,    -5,   -14,   -16,    -3,     2,     2,     6,     5,     2,   -11,   -22,   -20,    -2,     7,     7,     4,   -10,     2,    -7,     0,    -4,     0,    -4,     3,     5,     2,     3,    -1,    -2,    -8,    -5,    -7,    -1,     6,     6,     4,     3,   -17,   -23,   -10,     3,    10,    10,     1,   -12,     1,    -9,    -3,    -4,    -1,    -5,     0,     6,     4,     4,    -1,    -2,    -5,    -8,   -10,     1,     4,     9,    -3,   -11,   -20,   -11,    -2,     5,     3,    -1,    -1,    -4,     2,    -6,    -1,    -2,    -2,    -6,     2,     0,     3,     8,     0,    -4,    -5,   -10,    -3,     0,     7,     4,    -2,   -11,   -10,    -4,     4,     4,    -2,     2,    -2,    -3,     3,    -5,     1,    -2,    -6,    -7,    -2,     0,     1,     1,    -6,     2,    -2,    -8,     3,    -1,     6,     2,    -2,    -6,    -7,     0,     2,     0,     1,    -4,     1,     3,    -1,    -5,    -1,     1,    -5,    -3,    -5,     2,    -1,    -2,     1,     3,    -1,     2,     2,    -6,     1,     1,    -3,    -7,    -5,    -1,     0,     1,     2,     0,    -5,     0,    -4,    -9,     0,     0,    -4,   -13,    -4,     3,    -2,     0,     2,     1,     3,    -5,     2,     1,    -1,    -3,    -4,    -4,    -6,     1,     2,     1,     1,    -5,    -1,    -4,   -10,    -7,    -1,     1,    -4,    -9,    -6,    -1,     0,     2,     0,     3,     8,     0,    -6,     3,    -6,    -4,     3,     0,    -2,     3,     0,     1,     0,    -1,    -6,    -8,    -9,    -1,     1,     0,    -4,    -8,    -2,     0,     4,     0,     0,     3,     4,     1,     0,     4,     2,    -3,     0,     4,    -2,     0,     1,     3,     3,    -3,     0,    -5,    -2,     1,    -1,    -1,     0,    -8,    -1,     1,     2,     6,     5,     4,     4,     3,     3,     0,     2,    -1,    -4,     1,     1,     1,    -2,    -3,     1,     0,    -3,    -4,    -2,     2,     1,    -1,    -1,    -6,    -4,     2,     6,     7,     3,     0,    -3,    -1,     0,    -1,     0,     5,     2,     1,    -1,     0,     2,    -2,    -5,    -5,    -2,    -3,    -7,    -2,     0,     0,    -2,    -4,    -2,     0,     2,     0,     4,    -3,     0,    -3,     0,    -1,     5,     2,     1,    -2,    -3,    -3,    -3,    -2,    -1,    -3,    -7,    -6,    -4,    -3,    -4,    -1,     0,     5,     4,    -2,    -4,    -5,    -3,     2,    -8,    -8,    -4,     1,     4,    -1,    -2,    -3,    -2,    -5,    -9,    -4,    -4,    -5,    -3,    -5,    -2,    -3,    -1,    -3,    -3,     8,     2,   -11,    -8,    -4,    -2,    -1,   -11,    -7,    -4,    -6,     0,    -1,    -3,    -2,     3,    -4,    -7,    -8,    -6,    -7,     0,    -4,    -2,    -2,     0,     0,     0,    -3,     0,    -3,    -3,    -4,    -7,     2,    -5,    -1,     0,    -6,     5,     1,    -3,     0,     5,    -5,   -11,     0,    -3,    -2,     3,    -5,    -1,     1,     0,     0,    -3,   -10,    -5,     1,    -6,    -7,     2,     2,    -1,     1,    -2,    -9,     0,    -3,    -1,    -3,     1,    -2,    -8,    -1,    -3,     1,     1,    -6,    -3,     0,     0,    -1,     1,    -6,    -6,     1,    -1,     2,     4,    -4,    -2,     0,    -3,    -5,    -2,    -3,     1,    -4,     1,     5,    -2,     1,     3,    -1,     4,     1,     1,     1,    -1,     0,     0,    -3,    -4,    -9,    -2,     2,     2,     0,     7,     3,     2,    -6,    -4,    -6,    -6,    -4,     1,     2,     4,    -1,    -3,     0,     2,     3,     0,     1,     0,    -1,     0,     0,    -7,    -6,     3,     2,     2,     1,     1,     6,     5,    -4,    -1,    -1,    -9,     0,     2,     2,     5,     1,     5,     2,    -1,     7,     1,    -1,     1,     0,    -1,    -1,    -5,   -11,     2,     0,     0,    -1,     3,     4,    -9,   -13,    -4,     1,    -8,     2,    -5,    -8,     0,     1,     4,     0,    -1,    -2,     0,     1,     1,     0,     1,    -6,    -2,    -6,    -7,    -3,    -4,    -5,    -7,    -5,    -6,    -9,    -2,     1,    -2,     2,    -6,    -8,    -9,   -10,    -7,     0,    -1,     1,     0,     1,     0,     0,     0,     1,     0,    -1,    -2,    -3,    -3,    -2,    -6,    -5,    -4,    -5,    -8,    -1,    -4,    -6,    -6,    -5,    -7,    -4,    -5,    -1,     0,     0,     0,     0),
		    55 => (   -1,     0,     1,     0,     0,     1,     0,     1,    -1,    -1,     1,     0,     0,    -2,     1,     1,     1,    -1,     0,     0,     1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,     0,     0,    -1,    -4,    -2,    -2,    -5,    -6,    -6,    -6,    -5,    -5,    -7,    -7,    -2,    -1,     0,     1,    -1,     0,    -1,    -1,    -4,    -4,    -2,    -2,    -4,    -4,    -6,   -10,    -9,   -10,   -13,   -16,    -8,     3,     3,     5,     2,    -2,    -1,    -6,    -6,    -1,    -5,    -4,     1,    -1,     1,     1,    -2,     0,    -2,    -6,   -11,    -7,   -15,     3,     6,    -1,     2,     0,    -4,    -7,    -6,     0,     3,     7,    -1,     6,     0,    -5,    -3,     3,    10,     0,    -1,    -3,    -5,     0,    -7,    -1,     0,     1,     0,    -1,     2,    -1,     2,    -3,    -2,    -4,    -6,    -4,     4,    -6,    -5,    -1,    -3,    -3,    10,     7,     1,    -3,    -1,     1,    -5,     0,    -5,    -2,    -4,     1,    -4,     0,     0,     9,     7,    -2,     3,     5,    -1,    -5,   -11,    -2,    -1,     0,     1,     5,     0,     6,     2,    -1,     1,     0,     0,    -7,    -7,    -4,     0,     3,     3,    -1,     0,     6,     8,     1,     1,    -3,    -4,    -6,    -6,    -1,    -2,    -2,     2,     8,     8,    10,    -1,     1,     1,    -4,     1,   -12,   -11,    -5,     3,     8,     7,     6,     6,     2,    -1,     1,     3,     0,     5,     2,    -7,    -2,     2,     0,     1,     0,     2,     2,    -2,     4,    -1,    -3,    -9,   -15,    -8,     5,     0,    -6,    -1,     2,     2,    -1,    -1,     1,     4,     5,    -1,     3,    -5,   -10,    -3,    -3,     1,     0,    11,     4,    -8,     2,     0,    -1,    -7,   -11,    -4,     4,     2,    -7,     1,    -3,     1,     8,     5,     8,    11,     7,     1,    -3,   -11,   -12,   -12,    -6,     2,     0,     6,     7,    -4,    -3,     0,     0,    -9,   -19,     7,     7,     4,     2,    -3,    -2,     4,     7,    12,     8,     8,     9,     0,   -11,    -6,    -8,    -8,    -5,   -15,   -13,     5,     7,     7,    -4,     1,    -2,    -1,    -4,     2,     4,     3,    -1,    -2,    -3,     0,     3,     5,     6,     2,     6,     3,    -1,    -4,   -10,    -6,    -4,   -16,   -18,    -1,    -1,     3,     1,    -1,    -1,    -2,    -3,     5,     2,     0,     1,     0,    -1,     0,    -6,     1,     1,    -1,     1,    -4,    -4,     0,    -2,    -7,    -2,   -11,    -8,   -18,    -7,     7,    -7,     0,     0,    -3,    -1,     0,     4,    -3,     0,    -1,    -1,     0,     3,     1,     1,    -1,     2,    -2,    -6,     0,     3,     1,     1,    -3,    -9,   -14,   -11,     0,    -5,     1,    -1,    -1,     1,    -7,    -1,    -2,    -2,    -3,    -1,    -1,    -3,     0,    -4,     1,    -3,     3,    -1,    -3,     1,     3,    -1,     0,     8,     1,    -7,    -4,    -3,     0,     1,    -4,    -3,     1,     0,    -1,    -1,    -9,    -6,     1,    -1,     1,    -3,    -1,     0,    -2,    -1,     1,    -3,    -4,    -9,     0,     8,     4,    -7,    -7,    -8,     0,    -2,    -9,     8,     1,     3,   -10,   -15,    -7,    -8,    -4,     7,    -1,    -1,    -2,    -5,    -2,    -5,     0,     2,    -3,    -3,    -1,     4,    -2,   -15,    -9,    -9,     0,    -2,   -13,    13,     3,     0,    -3,   -14,    -9,    -7,    -3,    -1,    -5,    -3,    -4,    -3,     2,     5,     2,     5,     0,     0,     1,     3,    -8,   -15,   -12,   -12,    -2,     1,    -9,    13,    13,     7,    -1,    -8,   -11,   -15,    -2,    -6,    -4,    -6,     0,    -1,     3,     4,    -1,    -3,     3,     4,     4,     7,    -1,    -2,   -13,    -4,     0,    -3,     7,     1,    10,    10,     3,    -5,    -2,    -9,    -4,    -4,    -1,    -1,     0,     3,    -3,     2,     7,     0,     8,     0,     5,     7,     8,     5,    -8,    -9,    -1,    -4,     5,    -1,     5,     5,     1,     0,     1,    -1,    -5,     0,    -1,     4,    -1,    -3,     4,     6,     1,    -5,     4,    -1,    10,     4,     4,     8,    -7,     0,    -1,    -1,    -7,   -12,    -1,     5,    -3,    -4,     5,     4,     0,    -2,    -3,     0,     2,     6,     6,     3,     6,     5,     1,     6,    -1,     6,     3,    11,     4,    -2,    -1,    -1,   -10,    -4,    -8,    -7,    -4,     1,     1,     3,     3,    -1,     0,     2,    -2,     0,     2,     0,     1,     5,    -3,     0,     0,    11,    11,    14,     9,     0,     1,     1,     2,     2,    -3,    -2,     1,    -2,    -6,     0,    -2,    -1,    -3,     2,     2,    -1,     2,     2,     4,     5,    -2,     2,    -3,     8,     8,    10,     6,     0,     1,    -1,    -6,    -2,    -5,    -3,    -4,     3,     3,     9,     6,     5,    -1,    -4,    -7,     1,    -2,     6,     5,     6,     2,    -3,     2,     0,     9,    -6,    -3,     0,     1,     0,     0,     5,    -9,   -12,    -4,    -2,     2,    -4,    -6,    -6,     0,    -3,    -7,     0,     7,     9,     8,     6,     1,     7,    11,     9,     9,    -3,    -1,    -1,     1,     1,    -1,    -3,    -4,    -9,   -12,   -11,    -4,    -1,     3,     2,     0,    -2,   -10,     3,    -2,     3,     3,    10,     3,     0,    -2,    -5,    -3,     1,     1,     1,    -1,     1,     1,     0,    -2,    -2,    -1,    -2,    -2,    -3,     1,     1,     2,     1,   -12,    -9,    -3,    -4,    -3,    -6,    -7,    -8,    -4,    -1,     1,     1,     1,     0),
		    56 => (    0,     0,     0,    -1,     1,    -1,     1,     0,    -1,     0,     0,    -1,     2,     3,    -1,     1,    -1,     1,     1,     0,     1,     0,     1,     0,     0,     0,     1,    -1,     1,     0,     0,    -1,    -1,    -1,     3,     3,     6,     4,     3,     2,     1,     4,    -1,    -2,    -1,    -1,     0,     1,     7,     4,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     4,     0,     2,     6,     5,     5,     3,    -2,    -3,    -3,    -3,    -1,     0,    -1,    -1,     3,     4,     5,     4,     7,     3,     3,    -1,    -1,    -1,    -1,    -6,    -6,    -1,     4,     4,     3,     2,     3,    -1,    -4,    -6,   -11,    -5,    -3,    -1,    -5,     2,     7,     4,     3,     1,     6,     5,     1,    -1,     0,     1,     0,    -7,    -7,     5,     7,     4,     1,    -2,     2,     1,    -6,    -8,   -12,    -8,    -1,    -2,    -3,    -8,     0,     1,    -2,    -5,     0,     5,     4,     8,     8,    -1,     1,    -4,    -6,    10,     6,     2,     1,     2,     1,     0,    -3,    -5,    -9,    -3,     3,    -2,     1,    -3,    -4,    -4,    -2,    -3,     2,     3,     4,     9,     6,     0,     0,     2,    -1,     8,     2,     4,     1,     8,     4,    -4,    -8,    -8,    -9,    -2,    -3,    -7,    -3,     0,    -7,    -4,     0,    -1,     0,     1,    -5,     2,    10,     0,     0,     1,    -2,     8,     3,    -1,     5,     4,     5,    -3,    -7,   -10,    -5,     0,    -7,    -8,     0,     0,    -1,    -1,    -4,    -4,    -5,    -5,    -2,     4,     9,     0,     0,     1,    -3,     6,     2,    -2,     3,     1,    -1,    -6,   -10,   -11,     0,     1,    -8,    -1,     3,     2,     3,     3,     1,    -4,    -1,    -1,    -3,     4,    -5,    -1,    -1,    -1,    -5,     4,     1,    -2,     3,    -1,    -5,   -10,   -12,   -10,    -3,    -1,    -3,     2,     6,     1,     2,     4,     0,    -2,     1,    -1,    -5,    -2,    -2,    -1,    -1,    -2,    -5,     6,     4,     2,     7,     1,    -5,    -8,   -10,    -8,    -2,    -1,     1,     1,     5,    -4,    -2,    -3,     2,     0,     1,    -2,    -2,     0,    -1,     0,     1,     1,    -1,     5,     5,     3,     2,    -1,    -4,    -6,    -8,    -4,    -1,     1,    -1,    -2,    -9,    -6,    -2,    -4,     0,     2,     3,     1,     1,    -2,    -3,    -1,     0,    -1,    -3,     3,     7,     0,     2,    -1,    -4,    -6,    -8,    -2,     9,     2,     1,     1,    -3,    -3,    -5,    -2,     3,     5,     4,     3,    -1,    -1,    -5,     1,     1,    -1,    -2,     1,     1,    -1,     0,     2,    -3,    -4,    -9,     0,     5,    -2,    -5,    -1,     0,    -3,    -3,    -2,     2,     2,     4,     3,     0,    -1,    -1,    -1,     0,     1,    -3,     1,     2,    -2,     2,     0,    -1,    -5,    -3,     4,     6,    -8,    -6,     0,     1,    -1,    -1,    -5,    -2,     1,     3,     2,     0,    -2,    -2,    -1,     0,     0,    -2,     3,     1,    -2,    -1,     0,     0,    -4,     0,     0,     3,    -3,    -1,     1,    -2,    -1,    -5,    -5,     0,     2,     5,     2,    -1,     1,    -8,     1,     1,    -2,    -1,     4,     1,    -4,    -3,    -3,    -2,    -2,    -2,     3,     0,     2,     6,     1,     1,     3,    -5,    -3,    -1,     3,     2,    -1,     1,     0,    -4,     0,     1,     0,     3,     0,     1,    -2,    -3,    -2,     0,     2,     0,    -2,     3,     0,     1,     7,     0,     3,    -1,    -4,     0,    -1,     3,     0,     0,    -1,    -3,     1,     0,    -1,     1,    -2,     1,    -5,    -4,    -4,    -1,     0,     3,    -3,     1,    -3,     3,     2,     1,     5,     2,    -1,    -2,     2,     3,     0,    -1,     0,    -3,    -1,    -1,    -1,     4,     1,    -1,    -5,    -6,    -5,     0,     0,     0,    -2,     0,     1,     3,     0,     1,     5,     5,     3,     1,     0,    -4,    -2,     1,    -5,    -1,     0,    -2,    -1,    -3,    -3,    -4,    -1,    -7,    -6,    -2,     1,    -2,    -2,     2,     1,     4,     2,     5,     4,    -3,     0,    -3,    -7,    -4,    -3,     2,    -2,     0,    -1,     1,    -1,    -3,    -1,    -4,     0,    -4,    -3,     1,     0,     0,     0,     4,     2,     2,     2,    -3,    -4,    -2,     0,    -2,    -4,    -3,    -3,    -3,    -1,     1,     0,    -1,     0,    -3,     0,    -2,    -5,    -3,     1,     0,    -2,    -3,     0,     3,    -2,     1,    -1,    -2,    -7,     1,     0,    -4,    -5,    -6,    -6,    -2,     0,     1,     0,     1,     0,    -2,    -2,     0,    -2,    -3,    -2,    -3,    -1,    -4,     0,    -5,    -3,     2,    -3,    -7,    -3,    -3,    -2,    -1,    -4,    -4,    -5,     0,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -2,     1,     0,    -2,    -1,    -4,    -2,    -1,    -1,    -2,    -1,    -1,    -1,    -3,    -6,    -3,    -2,    -1,    -1,     0,     0,     1,    -1,    -1,     0,    -1,     1,    -1,    -2,    -3,    -2,    -1,    -2,     0,    -1,    -2,    -1,     0,     0,    -1,     0,     0,    -1,    -4,    -2,     0,     2,    -1,    -1,     0,     0,    -1,     1,     0,     1,    -1,     0,     0,     0,    -1,     1,    -1,     0,     0,     0,     1,     0,     1,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,     1,     1,    -1,     0,     1,     0,     1,    -1,     0),
		    57 => (    0,    -1,     1,    -1,    -1,     1,    -1,    -1,    -1,     0,     0,     0,     1,    -1,    -1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,     1,     0,     0,     0,    -1,     1,    -1,     1,     0,    -1,    -1,    -1,    -5,    -5,    -5,    -3,   -11,   -12,   -13,    -3,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,     1,     1,    -2,    -2,    -8,    -8,   -11,   -10,    -6,    -4,    -3,    -7,    -5,    -3,    -4,     0,    -6,    -6,    -5,    -4,    -4,    -2,     0,     0,     0,    -1,    -1,    -3,    -2,    -8,   -13,   -13,   -12,    -8,   -12,   -17,   -17,   -12,   -11,   -10,    -7,    -5,    -5,    -8,    -4,    -6,   -19,   -12,    -6,    -3,     0,    -1,     0,     1,    -1,    -5,    -6,    -9,   -13,   -18,   -19,   -23,   -25,    -4,    -1,    -2,    -3,    -6,   -13,   -18,   -15,   -10,    -7,    -7,   -11,   -15,   -16,    -9,    -2,     1,     1,     1,     0,    -7,   -10,    -4,    -8,    -5,    -1,     3,    -3,     3,     5,     4,     0,    -1,    -3,    -9,   -12,   -16,   -16,   -10,   -11,   -23,   -17,   -15,    -1,     0,     0,    -1,    -4,    -3,    -2,     3,     2,     2,     0,     2,     7,     6,     0,     1,    -6,    -2,     2,    -4,    -1,    -7,    -9,    -4,    -7,    -8,   -10,   -11,    -6,    -5,     1,     4,    -3,     1,    -1,     9,     5,     6,     5,     5,     7,     0,     3,     4,     4,     1,     3,     4,     6,     3,    -2,    -1,    -2,    -3,    -8,   -16,   -10,    -6,    -4,     3,    -1,     5,     0,     8,     1,     2,     1,    -3,     4,     4,    -5,    -7,    -5,     3,     4,     3,     5,     4,     3,     3,    -2,     0,    -7,    -9,   -10,    -4,    -1,     3,     4,     3,     5,     1,    -2,    -1,     0,    -2,     1,     3,    -1,    -2,    -6,     0,     1,     6,     5,     1,     0,     5,     2,     4,    -7,    -2,     9,    13,    -1,     6,    -1,    -3,     3,    -6,     1,    -3,     1,     2,     0,     3,    -4,    -6,    -1,     1,     5,     5,     6,     4,     3,    -1,     4,    -1,    -1,     5,     8,    11,    -1,     0,     0,    -3,     4,     3,    -4,    -3,    -1,     4,     2,    -4,    -2,     5,    -1,     0,     4,     2,     5,     3,    -3,     1,     6,     4,    -2,    -8,     0,     7,    -1,     3,     5,     1,     5,     7,     1,    -5,     5,    -2,    -5,    -2,    -2,    -2,    -2,     6,     4,     5,     2,     0,    -1,     1,     0,     3,     1,     4,     7,    11,     0,     2,     7,     0,     5,     6,    -2,    -3,     2,     0,     0,    -1,    -3,     0,    -3,     2,     1,     1,     0,     1,    -2,    -1,     6,     2,     6,     6,    -1,    -3,     0,     3,     2,     1,     0,     4,    -5,     3,     3,    -1,     0,    -1,     1,    -3,    -2,     0,    -3,     3,     0,     3,    -2,    -2,     1,    -2,    -2,   -12,   -11,    -2,     1,     0,    -1,    -1,    -3,    -4,     0,     1,     1,     3,     3,     2,    -2,     1,     3,     4,    -3,     0,     2,     3,    -1,     0,    -4,    -7,   -10,   -12,    -1,    -8,     0,     0,    -2,    -6,     1,     3,    -3,    -4,    -2,     2,     3,     0,     2,     7,     4,    10,     2,     1,     0,    -3,    -4,    -3,    -1,    -2,    -5,   -11,    -8,    -8,    -1,    -1,    -4,    -9,     2,     1,    -1,    -5,    -4,    -8,    -2,    -3,     5,     6,     4,     4,    -1,    -3,    -4,    -3,    -2,    -2,     0,    -1,     5,    -7,    -4,    -9,     2,     1,     2,   -14,     1,    -1,    -6,    -4,    -4,    -4,    -4,     0,     1,     2,     2,    -3,    -8,     1,     0,    -3,     6,     5,     2,     6,     2,   -10,     1,    -6,     1,     1,    -1,    -5,    -4,    -1,    -3,    -7,     0,    -4,    -5,    -1,     3,     4,    -1,    -8,    -1,     0,    -1,    -1,     2,     7,    -2,    -5,     4,   -11,    -9,    -3,    -1,    -1,    -3,    -3,   -11,    -8,    -7,    -5,    -8,    -3,    -8,    -8,    -3,     2,     1,    -4,    -1,     1,    -9,    -1,     1,     2,    -4,   -11,    -4,    -9,    -8,     1,    -1,     0,    -4,    -8,   -10,    -1,    -3,    -3,    -3,    -7,    -2,    -3,    -2,     2,    -3,    -2,     1,     0,    -7,    -3,    -4,     5,    -4,    -9,   -13,    -3,    -2,     0,    -2,    -2,    -6,    -7,     0,     1,     0,    -3,     3,     0,    -3,    -1,     1,    -3,     0,     1,     6,    -1,    -2,     2,     5,     0,    -6,   -24,   -13,    -1,    -4,     0,     0,    -1,    -5,    -8,     2,     2,     2,     1,     5,     3,     0,     2,     7,     4,     8,     1,     4,     4,     0,     0,     4,    -1,    -6,   -21,   -11,    -6,    -9,    -1,    -1,     1,     4,    -3,     8,     8,     8,     7,     7,     0,     4,     5,     6,    13,    11,     1,     7,     5,     1,     4,     4,     2,    -2,   -14,    -8,    -8,    -6,     1,     0,    -1,    -1,     3,     3,     5,     4,     5,     4,     5,     9,     9,     7,     6,     2,    -3,    11,     4,     3,     3,     0,     6,     7,    -2,    -2,    -6,    -4,     1,     0,     1,     1,    -4,    -3,    -6,     0,     4,     5,     7,     7,     8,     7,    -6,   -11,    -1,     4,     1,     2,     7,     4,     6,     7,     2,    -3,    -1,    -1,     0,    -1,     1,    -1,     0,     2,     3,    -2,    -3,     0,     3,     6,     1,    -1,    -8,    -2,     2,    -3,     4,     2,     3,     2,     6,     3,     8,     1,     0,    -1,     0),
		    58 => (    1,     0,     0,     0,     1,    -1,    -1,     1,     0,     1,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,     1,     0,     1,     0,     1,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,     1,     0,     0,     0,     0,     1,    -2,    -3,    -2,    -3,    -1,    -4,    -4,    -4,    -2,     1,     1,    -1,     1,     0,     1,     0,     1,    -1,    -1,    -1,     0,     0,    -1,    -2,    -3,    -8,    -7,   -11,    -5,    -1,    -1,    -4,    -4,    -6,     1,     1,    -3,    -3,    -3,    -3,    -1,    -1,    -1,     0,    -1,     0,     0,    -2,    -3,    -2,    -4,    -8,   -15,     1,     4,     4,    -1,    -4,    -5,    -3,     4,    -5,    -6,     1,    -4,    -3,    -3,     3,     7,     0,    -2,    -4,     1,     0,    -4,    -3,    -9,    -8,    -9,    -5,     5,    11,     9,     7,     4,    -1,    -1,     3,     4,     3,     8,    -1,    -5,    -7,    -8,    -4,    -7,    -9,     1,     5,    -2,     0,     1,    -6,    -8,    -6,    -9,    -1,    13,     5,     5,     3,     6,     7,     3,     1,     2,     3,     7,     0,     8,     0,     1,     3,    -2,    -3,    -2,    -7,    -3,     1,    -1,   -10,    -8,    -9,    -4,    -3,     6,    -3,     1,     5,     1,    -1,     2,    -1,     2,     0,    -2,     2,     2,     5,     0,    -1,     4,    -3,    -4,    -2,    -2,     0,    -7,    -8,   -10,    -8,    -6,     0,     1,    -1,     0,    -1,     5,     0,     2,    -5,     3,     2,    -1,    -2,     1,    -3,    -1,    -2,     9,     6,    -9,    -6,     3,     2,    -5,    -7,     1,    -1,    -1,    -1,     5,     2,     1,     1,     0,    -1,     1,    -1,    -1,    -1,     0,     3,     8,    -3,     7,     5,     9,    10,    -6,     8,     9,     1,    -2,    -9,     2,     5,    -3,     0,     4,     2,     0,    -3,     0,    -1,     0,     3,    -1,    -2,     2,     1,    -1,     6,     5,     6,     4,     2,    -3,     8,   -10,    -1,    -1,   -11,    -8,    10,     3,    -4,     3,     4,     2,     5,     2,     2,    -1,     5,    -8,    -6,     1,    -1,     0,     2,     6,     3,     6,     4,    -8,     3,    -4,     1,    -1,    -5,     0,     9,     8,     2,     6,     2,     1,     2,     0,    -3,    -2,     2,    -7,    -6,    -5,     1,     0,     3,     4,     4,     5,     6,     2,    10,    -2,    -1,     1,    -8,     2,     9,    16,     0,     1,     6,     2,     0,    -3,    -5,    -5,    -1,    -4,     0,     0,    -4,    -2,     3,     4,     8,     1,     4,    -4,     5,    -9,     1,    -1,    -5,    -1,     3,     9,     3,     2,     4,     1,    -1,    -1,    -1,    -2,    -1,     1,     0,    -7,    -3,    -3,     4,     2,     7,     0,    -5,    -5,     4,     1,     0,    -2,    -2,    -6,    -9,     1,     6,    -8,     4,   -10,    -7,    -2,    -4,    -5,     0,     1,    -3,    -7,     0,    -6,    -8,     3,     0,    -2,    -7,    -1,    -4,    -3,     1,     1,    -3,     3,   -15,    -4,    -5,    -6,     2,    -6,    -2,    -2,    -7,     1,     3,    -4,    -3,     1,    -5,    -2,    -4,    -7,    -2,    -8,   -11,    -2,   -11,    -7,     1,    -1,    -2,     4,   -14,    -6,    -7,   -12,    -6,    -1,    -7,    -5,    -1,     4,     0,    -2,    -5,   -10,    -5,    -1,    -5,    -8,    -4,    -3,    -4,    -4,   -13,    -7,     0,    -1,    -3,    -7,    -4,    -7,    -8,    -8,    -1,    -5,    -5,    -8,    -2,    -2,    -4,    -7,    -4,    -3,    -3,    -2,     1,    -2,    -2,    -1,    -1,   -12,    -6,    -9,    -1,    -2,    -5,   -13,     0,    -7,     0,     2,     1,    -1,    -2,    -3,     1,     0,    -5,   -13,     0,     1,     0,     2,    -1,    -2,     1,     0,     0,   -11,    -5,    -6,     1,     1,    -9,   -12,    -3,    -7,    -4,     2,     8,     2,     1,    -3,    -5,    -4,    -8,    -5,    -2,     6,     1,     3,     3,    -4,     2,     6,     8,   -15,   -11,    -7,     0,     0,    -4,   -10,    -8,     2,     4,     1,     7,    -3,     7,     0,     3,     0,    -5,    -2,     6,     4,     1,     0,     5,     5,     5,    12,     3,   -18,   -11,     1,    -3,    -5,    -4,    -5,    -6,     1,     8,     1,     5,     8,     4,     3,     2,     5,     4,    10,     0,     7,    -7,     3,     1,     1,     9,     8,    -3,   -14,    -9,     0,    -3,    -4,    -2,    -4,     4,     8,     5,     8,     7,     7,     9,     9,     4,     7,    11,    12,     2,     1,     3,    -3,     0,     0,     8,     5,    -4,    -1,    -9,    -1,    -1,     1,    -1,    -2,     8,    -1,     3,    -2,     4,     4,     1,     1,     8,     8,     7,     8,     7,     6,     7,    10,     2,    -3,    11,     5,    -3,    -1,    -9,     0,     1,     0,    -4,    -5,    -3,    -3,    -2,    -3,     3,     5,     2,     1,     7,     2,     3,     5,    11,    -1,    -1,    -1,     1,    -5,     1,     2,    -5,   -12,    -6,    -1,     1,     0,    -4,     0,   -15,   -12,    -1,    -1,    -5,    -9,    -5,    -5,    -3,    -2,     3,     4,    -1,    -3,     2,    -1,    -8,    -8,    -8,    -4,    -5,    -3,    -2,     0,     0,     1,     0,    -3,    -7,   -12,   -11,    -3,     2,     1,    -6,    -3,     3,     2,   -10,   -20,    -9,    -5,    -5,   -15,   -13,    -6,    -7,    -3,    -1,     0,     0,    -1,     0,     0,    -1,     1,    -3,    -2,    -3,    -2,    -4,    -4,    -1,    -1,    -5,    -8,   -10,    -8,    -4,    -6,    -3,    -4,     0,     0,    -3,     0,     0,    -1,     0,     0),
		    59 => (    1,    -1,     1,     0,    -1,     1,    -1,    -1,     1,     0,     1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,     1,     1,     1,     1,    -1,     0,     1,     0,    -1,    -1,     1,     0,     0,    -1,     0,     0,    -1,    -2,    -3,     1,    -2,    -1,    -2,     0,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     1,     0,    -1,     0,     1,    -1,     1,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -4,    -1,     1,    -1,     1,    -1,    -1,     1,    -1,     0,    -1,    -1,     0,     1,     0,    -1,     1,    -1,    -2,    -2,    -2,     0,    -3,    -5,    -2,    -4,    -1,    -5,    -4,    -4,    -1,     1,     2,     0,    -5,    -4,    -2,    -1,     0,    -1,     0,     1,     1,     0,     1,     0,     0,    -1,    -5,    -2,    -1,     0,    -3,     0,    -7,   -10,    -8,    -7,    -5,    -5,    -3,    -7,    -8,     0,    -1,     0,    -1,    -5,    -4,    -1,    -1,     0,     0,     0,    -1,     1,    -1,    -3,   -10,    -4,    -5,     0,     1,     0,     2,     0,    -2,    -8,   -10,    -5,    -1,    -2,     0,     0,     1,    -5,    -2,     1,    -1,     1,    -1,    -1,    -4,    -5,    -5,    -7,    -2,     3,     1,     6,     6,     5,    -1,    -3,     4,    -2,   -12,   -12,    -6,     0,     0,    -1,     0,     0,    -1,    -3,    -1,     0,    -1,     1,    -2,    -6,    -9,    -7,    -1,    -4,     2,     5,     1,     3,    -3,    -8,    -6,    -6,   -13,   -17,    -6,     1,     0,     0,    -2,     0,    -1,    -3,    -2,    -1,    -2,     3,     1,    -6,     5,    -1,     5,     0,     0,     1,    -2,     1,    -1,    -6,    -6,    -3,     2,    -4,    -9,    -2,    -2,    -2,    -3,    -1,    -1,     0,    -1,    -4,    -4,     2,     0,    -4,     4,     4,     2,     3,     5,    -3,    -3,     1,     1,    -5,    -8,     3,     3,    -3,    -6,    -5,    -6,    -2,    -4,    -6,    -3,    -3,     0,    -1,    -2,     2,    -1,    -6,     5,     3,     2,     1,     1,   -11,    -9,     2,     6,    -1,     4,     0,     0,    -3,    -5,    -6,    -7,    -4,    -4,    -5,    -1,    -5,    -1,    -7,    -3,     3,    -3,    -7,     2,     6,     4,     1,    -2,    -1,     4,    13,     0,    -1,    -1,     4,    -2,    -1,    -9,   -10,    -6,    -6,    -2,    -4,     0,    -4,     1,    -3,    -3,     4,    -2,     2,     2,    -1,     0,     5,     2,     1,     4,     9,    -3,    -7,    -1,     4,     0,     0,    -4,    -6,    -9,    -7,    -4,    -3,    -4,    -5,     1,    -3,    -2,    -3,    -4,     0,    11,     2,    -5,     1,     2,    -2,     0,    -2,    -2,    -2,     0,    -1,    -4,     2,    -4,    -5,    -5,    -5,    -2,    -3,    -3,     0,    -1,    -1,    -2,    -2,    -3,    -3,     7,     1,    -3,    -2,     5,     0,    -4,    -2,     2,     2,    -1,     0,     0,     0,    -4,    -7,    -7,    -7,    -3,    -5,     0,     0,    -1,     0,    -2,    -3,     4,    -5,    -5,     1,    -1,    -4,     3,     1,    -3,    -7,    -3,     2,     2,     0,    -2,    -2,   -11,   -10,    -7,    -6,    -2,    -1,     0,    -3,    -1,     0,    -4,    -1,     0,    -3,   -11,    -1,     2,    -4,     1,    12,     4,     2,     1,    -5,    -4,    -4,    -2,    -4,   -15,    -6,    -3,    -2,    -2,    -1,     0,    -5,    -1,    -1,    -4,     0,     0,    -4,    -8,   -10,    -1,    -8,    -3,     3,     6,     4,     1,     1,    -6,    -6,    -4,    -3,   -10,    -6,    -2,    -4,    -6,     4,    -4,    -2,    -1,     0,    -4,     0,     0,     0,    -3,    -6,    -8,    -8,    -8,    -3,     4,    -2,    -2,    -3,    -2,     0,    -6,    -2,    -4,    -7,     0,    -2,    -6,    -1,    -3,    -3,    -1,     0,    -3,    -1,     0,    -2,    -1,     0,    -2,    -1,    -7,   -10,   -10,    -9,    -7,     4,     2,     1,    -4,    -4,    -6,    -7,    -3,     0,    -4,     5,    -3,    -3,    -1,    -2,     0,    -2,     0,     0,     0,    -5,     0,    -5,    -5,    -9,   -12,    -7,     0,     1,    -1,    -2,    -3,    -4,    -3,    -2,    -3,    -3,     1,     3,    -4,     0,     1,    -1,     1,    -2,    -1,     4,    -1,    -2,    -1,     1,     1,    -1,    -3,    -1,     1,    -4,    -1,     0,     0,    -7,    -2,    -4,    -2,    -1,     2,     5,    -5,    -1,     0,    -1,    -2,     3,     0,     1,     2,     2,     2,     4,    -2,     1,     4,     2,     1,     2,    -1,     3,    -2,    -6,    -4,    -7,    -1,     0,     2,    -1,     0,    -1,     1,     1,    -3,     2,    -1,    -1,     3,     0,     2,    -2,     1,    -1,     0,     0,    -1,     4,     0,     2,     3,    -2,    -3,    -3,    -1,     2,     1,     1,    -3,     0,     0,     0,     0,     0,    -1,     1,     0,    -3,     0,    -3,     3,    -3,    -8,    -6,    -2,     2,     3,     2,     2,     3,     2,     0,    -1,     2,     1,     2,    -1,     0,     0,     0,     2,    -1,    -1,     0,     1,    -2,    -1,     2,    -4,    -5,    -3,     1,    -6,    -5,     1,     5,     1,    -5,    -6,    -5,    -5,    -2,    -2,     2,     0,     1,     1,    -1,     1,     2,     0,     0,     0,     1,     1,     3,    -3,    -6,     5,     0,     5,     3,     2,    11,     4,    -5,     1,     0,    -1,     2,     2,     1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     2,     3,     1,    -4,    -2,     1,     0,    -4,    -5,     9,     9,    -1,    -2,     4,     2,    -3,    -3,    -1,     0,     0,     1,     0),
		    60 => (    0,     0,     1,     1,     1,     0,     1,     1,     0,     0,     0,     1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,     1,     1,     0,    -1,     0,     0,     0,     1,     0,    -1,     1,     0,     0,     1,     0,    -3,    -2,    -3,    -5,    -2,     1,     1,    -7,     7,     9,     9,     0,    -1,    -2,    -1,     1,     0,     1,     1,     0,     0,     0,    -1,     1,     7,     9,    -3,    -4,     1,    -2,    -5,    -8,    -7,    -9,   -16,    -9,    -4,    -1,    -6,    -4,    -4,    -5,    -4,   -12,    -4,    -6,    -1,     0,     1,     1,    -1,     1,     8,     3,    -7,    -9,    -8,    -7,    -6,    -4,    -9,   -13,    -6,    -7,    -8,     3,     3,     0,    -6,    -6,    -9,   -13,    -6,    -5,    -5,    -9,     1,     0,     0,    -1,    -2,    -3,   -15,    -6,    -7,     1,     7,    -1,     1,    -7,     0,    -3,     3,     7,     3,    -1,     0,    -6,    -6,    -2,    -3,   -10,   -17,    -7,     1,     0,    -1,    -4,    -3,    -4,    -8,     3,    -1,     2,    10,     6,     5,     1,     1,     4,     4,     4,     4,     4,     0,     0,    -1,    -4,    -3,   -10,   -15,    -3,    -2,     1,     0,    -5,    -1,   -10,     3,     6,     6,     5,     4,     7,     3,     1,     0,     3,    -3,     1,    -1,    -5,     2,    -1,    -6,     0,   -12,    -7,   -18,    -5,    -2,     0,    -3,    -5,    -5,    -6,     0,     5,     5,    -3,     3,    -2,     1,     2,     2,    -6,    -6,    -3,    -1,    -2,    -5,    -2,    -5,    -1,     0,    -6,    -3,    -9,     2,    11,    -7,     0,    -8,    -7,     1,     1,    -6,     1,     2,    -3,    -5,     0,    -2,    -9,    -1,    -2,     5,    -1,    -3,    -3,     1,     0,     4,    -7,   -17,    -9,    -2,    -1,    -2,     4,     0,    -2,     2,    -6,    -3,    -1,     3,    -2,     2,     5,     2,     2,     4,     3,     4,     2,     3,     2,    -2,     0,     4,    -2,   -10,    -3,    -2,    -2,    -1,     5,     2,     1,    -4,    -1,    -4,     1,     4,    -1,    -2,     0,     4,    11,     8,     8,     9,    -2,     3,     2,    -3,     2,     4,     0,    -6,    -7,     0,    -1,    12,    -7,    -1,    -2,    -7,    -3,    -4,    -5,    -2,    -3,    -1,     3,    14,     5,     6,    15,    12,    10,     6,     5,     2,     2,     3,     7,    -7,    -8,    -1,    -1,     0,    -8,    -3,     4,    -7,    -7,    -8,    -6,    -1,    -3,     1,     7,    10,     7,     9,     6,     6,     6,     4,    -3,     0,     0,     2,     4,    -4,    -6,    -4,     0,     1,     0,    -3,     5,    -1,     1,    -4,    -1,    -5,    -4,     2,     3,     1,     0,     1,     0,    -2,    -1,    -2,    -3,     2,     1,     6,     2,     3,   -11,    -4,    -1,     0,    -1,   -10,    -4,    -2,    -5,    -1,     0,    -3,    -3,     0,    -3,    -2,   -10,   -11,   -11,    -5,     3,    -2,     4,     9,     9,     5,     8,     7,    -9,    -1,    -1,     1,    -6,    -9,    -2,    -4,    -6,     2,     0,    -7,    -6,    -5,    -7,    -7,   -15,    -8,    -6,    -2,    -3,    -1,     5,     4,     1,     4,     6,     8,   -10,    -8,    -1,     0,    -4,    -4,     3,    -2,    -6,     2,    -1,    -3,     0,    -3,    -6,    -8,    -8,    -1,    -7,    -6,    -2,     4,     3,    -2,    -3,    -6,    -1,    -3,   -14,    -3,     0,    -1,    -5,     0,     2,     1,    -4,     2,    -1,     2,     3,     5,     2,     5,    -3,    -3,    -5,    -1,    -1,     3,    -1,    -8,    -2,    -3,    -2,    -9,    -9,     2,    -1,     0,    -4,    -3,     5,     4,     3,    -2,     1,     5,     6,     2,     1,    -3,    -7,    -2,    -2,     2,     1,     1,    -6,    -5,    -3,     3,    -8,    -8,    -7,    -5,     1,     2,    -1,    -3,     0,     7,     4,     7,     6,     1,     0,     1,     6,    -3,    -4,     0,     0,     1,     1,     6,    -3,    -4,    -1,     3,     0,   -14,    -2,    -1,     0,     2,    -6,    -4,     7,     5,     4,     6,     3,     9,     0,     3,     8,     2,     1,     3,     0,     2,    -1,     1,    -5,    -7,    -3,    -2,    -5,   -16,     1,     0,     1,    -1,    -6,    -3,     1,    -1,     6,     9,     7,     5,     4,     1,     5,     0,    -1,     3,     2,     0,     2,     2,    -2,    -5,    -1,     1,    -8,    -8,    15,     0,    -1,    -1,    -3,    -4,   -10,    -6,    -1,     8,     7,     1,     9,     4,    -1,    -3,     2,     6,     3,     3,    -2,    -2,    -6,    -6,    -3,     0,    -5,    -3,     9,     2,     0,     1,    -3,    -7,    -2,    -7,    -5,    -1,     6,     5,     3,    -4,     5,    -1,     1,     3,     2,     6,    -1,    -7,   -11,    -7,    -9,    -3,    -6,    -8,    -8,    -1,     1,    -1,    -2,    -4,     2,     4,    -7,    -4,    -4,    -2,    -3,   -11,    -7,    -7,    -6,     4,    -1,     0,    -4,   -10,    -6,   -10,    -8,    -6,    -5,    -3,    -1,     0,     1,     1,    -1,    -2,   -10,    -6,   -11,   -16,    -9,    -9,   -10,    -6,    -9,    -6,    -6,    -8,   -18,   -16,   -16,   -18,   -12,   -14,   -10,    -4,    -1,     0,     1,     1,     0,     0,    -1,     0,    -3,   -10,   -14,    -7,    -5,    -9,    -7,    -8,    -5,    -6,    -8,   -12,   -10,    -9,    -9,   -11,   -10,   -11,    -7,    -5,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -6,     0,     0,     0,    -7,    -2,    -1,     0,     1,    -4,    -4,    -3,    -5,    -3,    -4,     0,     1,    -1,     1),
		    61 => (   -1,    -1,     1,     0,    -1,     1,    -1,     1,     0,     0,    -1,     0,     0,     1,    -1,     0,    -1,    -1,     0,     1,    -1,     0,     0,    -1,     0,     1,    -1,    -1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     1,     0,    -1,    -2,    -2,     2,     0,    -2,    -1,     0,     1,     1,    -1,     0,     0,     1,     0,     1,     1,     0,     1,     1,     0,    -1,    -1,    -1,     1,    -1,    -1,     0,     0,    -5,    -5,    -5,   -10,   -10,    -4,    -3,    -1,     3,    -3,    -2,    -1,    -3,    -3,     1,    -1,     0,     0,    10,     7,     1,    -2,     0,     4,     2,     1,    -2,    -1,    -8,   -20,   -15,   -12,    -8,    -7,    -5,     0,    -1,    -1,    11,     2,    -1,    -3,     0,     1,     1,    -1,     9,     7,     3,    -3,    -5,    -3,    -8,    -4,    -6,    -7,   -12,   -14,     6,     3,     5,     3,     3,     3,     1,     3,     3,    -4,    -6,    -8,    -7,    -5,     1,    -1,     6,    10,     6,     2,    -2,    -4,   -15,    -9,   -14,   -13,   -13,    -8,     0,     3,    -2,    -4,    -9,    -4,    -2,     2,     5,     0,    -5,    -8,    -7,    -7,    -1,     0,    -5,     4,     8,    -4,     6,     9,    -6,   -14,   -15,   -15,    -7,    -3,    -1,    -3,    -2,     1,    -3,    -2,     3,     0,     1,    -2,    -7,    -6,    -4,    -4,    -1,    -7,    -9,    -2,    -6,     6,     7,     9,   -10,   -10,   -22,   -13,    -7,    -3,     0,     0,     3,     3,     0,     5,     5,     1,    -4,    -3,    -8,    -5,    -4,    -3,     0,    -7,    -7,     3,    -6,     5,     6,     2,    -6,    -8,   -10,   -11,   -13,    -6,    -1,     4,     3,     3,     1,     3,     2,     1,    -3,    -6,   -10,    -4,    -9,    -1,     1,    -1,    -7,     1,    -3,    -4,     5,     8,     4,     2,    -2,   -13,    -4,    -9,    -1,     6,     9,     3,     3,     1,    -1,    -4,    -4,    -3,    -7,    -2,    -1,    -2,    -1,     3,    -7,    -3,    -3,    -7,     0,     6,    -2,    -1,     4,    -1,    -4,    -8,     0,     2,     4,     3,    -2,    -3,    -9,   -12,     0,    -1,    -6,     0,     0,     8,     1,     1,    -1,     4,     0,     6,     4,    -8,   -11,    -4,     3,    -3,   -11,     0,     1,     3,     2,     0,    -4,   -10,    -4,    -2,     0,    -2,    -1,     0,     0,     6,     0,     1,    -3,     6,    -2,     8,     7,    -3,    -4,     1,    -1,    -4,    -3,     3,     5,     1,     3,     3,    -6,    -8,    -3,     6,    -2,    -3,    -5,     4,    -1,     5,    -1,     0,    -2,     4,     2,     3,     6,     2,     4,     4,    -2,    -5,    -5,     0,     5,     0,     1,     5,   -10,   -17,    -9,     5,    -4,    -4,    -6,     0,     1,     1,    -1,     0,     4,     2,     8,    -4,    -4,   -12,     4,     0,     1,    -3,    -3,     2,     2,    -3,     3,    -2,     1,    -8,    -5,     8,     5,    -1,    -3,     7,     8,     0,     1,     0,     1,     9,     4,   -10,     0,    -1,     4,     1,    -2,     2,     0,     2,    -3,    -3,     6,     4,   -11,   -12,    -4,     1,    -1,    -4,    -6,     4,     4,    -2,     0,     1,     4,    -2,     0,     1,     0,    -7,     1,     0,    -9,     1,    -3,     3,    -1,    -1,     6,     1,    -7,   -12,    -7,     3,     0,     3,     4,     2,     0,    -2,    -1,     1,     0,    -7,     2,    -1,     1,    -2,    -3,    -4,    -6,     4,     1,     3,    -1,    -5,    -1,   -10,    -9,    -7,    -5,     2,    -3,     0,     2,     4,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -9,    -7,    -7,    -2,     0,    -1,     2,     1,     2,    -2,    -4,    -9,    -9,    -6,    -8,    -7,     1,     0,     4,     1,     4,     0,     5,    -1,    -1,     4,     2,     0,    -8,    -2,    -5,    -1,     4,     1,     2,    -1,     3,     0,     1,    -6,    -4,    -2,    -8,    -6,    -1,    -4,     4,     6,     7,     2,     5,     0,     0,     4,    -1,     4,    -2,    -1,    -4,     0,    -4,     1,     0,    -3,     2,     4,    -2,    -1,    -8,    -1,    -3,     4,    -3,    -1,     3,     9,     8,     1,    -1,     5,     6,     5,     4,     2,     5,    -3,    -1,     0,    -3,     2,    -4,     0,     0,     1,     1,    -5,   -10,     0,     4,     8,     3,    -1,     4,     7,     4,     0,    -1,     4,     6,     4,     3,    -1,     2,     1,    -6,    -5,    -2,    -4,    -4,     0,     0,     5,     8,     3,     1,     9,     4,     0,    -1,     2,     6,     1,    -1,     3,     0,     1,     1,     0,    -1,    -2,    -1,     5,     7,     9,     9,    -1,    -2,    -1,     2,     2,    10,     4,     6,     5,    -1,    -8,    -8,    -2,    -2,     3,     7,    10,    -1,     1,     0,     1,    -2,    -9,    -9,    -8,    -1,    -1,     9,    -3,    -2,    -3,     1,     1,     6,    -1,    -1,    -1,     2,    -1,     4,     1,    -4,    -3,     4,     3,     0,     1,     0,     1,    -2,    -5,    -4,    -3,   -13,     0,     6,   -16,   -13,     0,    -2,     5,    -2,    -7,   -13,    -7,    -4,    -7,    -5,    -4,    -3,    -1,     1,     0,    -1,    -1,     0,     0,     1,    -2,    -4,   -10,   -12,   -11,   -11,    -4,    -6,   -11,   -11,    -6,    -3,     3,    -7,    -1,    -2,    -1,    -2,     0,     0,     1,    -1,    -1,    -1,     0,     1,     1,     0,     1,     1,     0,    -1,    -1,    -2,    -5,    -4,     0,    -1,    -4,    -1,    -2,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     1),
		    62 => (   -1,     0,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     1,     2,     1,     1,    -1,     1,     1,     0,     1,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,    -1,     0,     0,    -1,     1,     1,     2,     1,    -1,     0,     0,    -1,    -3,     3,     1,     0,    -5,    -1,    -1,     0,     0,     0,     1,     0,     1,     1,     1,    -1,     0,    -2,    -1,     1,    -1,     1,    -1,     3,     9,     7,    11,     4,    -2,    -3,    -3,    -6,   -16,   -11,    -3,    -2,    -1,     0,     2,     0,     0,     0,    -1,    -1,    -4,    -4,     3,     6,    -1,    -1,     5,    -2,     1,    -2,     1,     0,     2,     5,     0,    -8,    -7,    -8,    -5,     4,     1,     0,    -1,     1,     0,     1,     1,    -3,     2,     3,     4,    11,    10,    -3,     1,     6,     6,     4,     9,     6,     6,     0,     1,     1,    -4,     2,     2,     1,    -7,    -7,    -3,    -4,    -1,     1,     1,     2,     0,    -1,    -4,    -3,     6,    -1,    -4,     2,     1,     3,     3,     0,     3,     4,     0,     1,    -1,    -5,     4,     8,     1,    -4,    -4,    -5,    -2,     1,     0,     3,     2,    -2,    -7,     2,     3,    -2,     0,    -1,    -3,     0,    -1,     3,     0,     0,    -4,     2,    -5,     1,     3,    10,     2,    -4,    -5,    -3,    -1,    -1,     0,    -1,     5,     0,    -2,    -7,     0,     3,    -1,     3,     0,     1,     2,     6,     4,    -1,    -3,    -3,    -7,     2,     0,     5,    -8,    -6,    -8,    -2,    -2,    -4,     3,     3,     1,     5,    -4,    -5,    -3,     2,     0,     5,     5,    -1,    -3,    -4,     1,     1,     1,    -1,     0,     0,     0,     1,     0,    -4,    -5,    -6,    -1,     0,    -3,    10,    -2,     4,     5,    -7,     1,    -1,     0,     0,    -4,     1,   -11,   -18,    -2,     3,     2,     0,    -1,     0,     0,     0,     3,    -9,    -5,     3,    -3,    -1,    -2,     5,     2,    -2,    -1,    -3,     6,     2,    -4,    -4,    -5,   -10,   -14,    -7,    -6,     1,     0,    -3,    -1,    -5,     2,    -8,     4,    -3,    -2,     3,    -1,     0,     0,    -2,     4,     5,    -2,     0,    -1,    -2,   -11,    -8,   -14,   -15,   -16,    -4,    -2,     0,    -5,    -6,    -5,    -2,    -3,    -4,     6,     0,     0,    -3,     0,     1,    -1,    -3,    -2,     0,    -1,    -5,   -13,   -10,   -12,   -12,    -9,   -12,    -4,    -1,    -4,     3,    -1,    -5,    -5,    -1,     0,    -4,     4,    -1,     2,     6,    -3,     0,     1,     4,     0,    -3,    -7,   -12,   -17,   -20,   -19,   -10,    -8,    -4,     5,    -3,    -4,     2,     0,    -3,    -7,    -6,    -2,    -5,     1,    -2,     0,     6,     1,     0,    -2,    -2,    -1,    -1,    -8,   -10,   -14,   -15,   -10,    -2,    -1,     1,     2,    -5,    -4,     0,    -2,    -6,    -4,    -6,    -1,     0,    -2,    -2,     0,     4,     4,    -1,    -3,     0,    -1,    -8,    -6,    -2,    -5,    -2,     4,     6,     4,    -3,     2,    -2,    -4,    -1,    -4,    -7,    -5,    -9,     1,    -1,    -3,    -1,     4,     4,     8,    -1,     0,    -1,    -3,    -7,    -5,     0,    -5,    -3,     2,     2,     3,     1,     1,     1,    -8,    -2,    -5,   -10,    -5,    -9,    -2,     0,     0,    -3,     9,     4,     3,     1,     0,     1,    -1,    -6,    -2,    -7,    -3,    -1,     0,     1,     3,     5,     3,    -1,    -3,    -5,    -8,   -12,    -7,     1,     0,    -6,    -6,    -5,     5,    -2,     3,     1,     1,    -3,     2,     6,    -1,    -1,    -2,     6,     4,     1,     2,     7,    -2,    -1,   -10,    -7,    -6,    -2,    -3,     1,     1,     0,    -4,    -3,    12,    -4,     8,     1,    -1,     2,     5,     5,     1,    -1,     4,     8,    -2,     4,     4,     7,     4,    -5,    -3,    -6,    -8,    -2,    -1,     0,     0,    -6,    -7,     4,     5,     7,     9,     0,    -1,     6,     7,     7,     6,    -6,     3,    -1,    -1,     2,     4,     5,     3,     0,     4,     1,     5,    -7,     1,     2,     2,     0,    -1,     4,     5,     6,     1,    -1,     3,     7,     6,     4,     4,    -4,    -3,    -3,     2,     2,     0,     3,    -1,     0,     2,     4,    -3,     1,     6,     1,     4,     4,     4,    12,    13,     4,    -1,     0,    -1,     6,     6,     2,     0,    -1,     1,     2,    -3,     3,     1,     2,    -1,     4,     4,     1,   -10,    -2,     3,     4,    -2,     3,    -4,     0,     2,    -5,    -3,    -1,    -1,    -1,     1,    -4,     3,     0,     2,     6,    -1,    -1,     3,     0,    -3,     2,     7,     2,    -6,     4,     2,     0,     5,     3,     5,     4,     3,    -4,     0,    -1,     0,    -4,    -2,    -5,    -7,   -12,   -18,   -11,    -5,     1,     1,     2,     2,     9,     1,    -4,     2,     6,     6,    -5,     3,    14,     8,     8,     3,     3,    -1,     0,    -1,    -2,    -1,    -2,    -4,    -3,    -6,   -11,   -12,    -2,    -1,    -2,     0,     6,     7,     4,    10,    -1,   -10,     1,     2,     2,     0,     4,     4,     3,     1,    -1,     0,    -1,     0,     0,    -1,    -3,    -3,    -3,    -2,    -1,    -5,     0,    -7,    -7,    -4,   -11,    -8,    -5,    -2,    -1,    -1,    -4,     1,    -1,    -1,     0,     1,     1,     1,     1,     1,     1,     1,    -1,     1,     1,     1,    -1,    -1,    -1,    -1,     0,     1,    -1,    -1,     1,    -1,    -3,    -2,     0,    -1,     0,    -1,     0,     1),
		    63 => (    1,     1,     1,     0,     0,     1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     1,    -1,     1,     0,     0,    -1,     1,    -1,     0,    -1,     0,     1,    -1,    -2,    -2,    -3,    -4,    -3,    -2,    -6,    -3,     0,     1,    -1,     1,     0,     0,     0,     0,     0,     1,     0,     1,    -1,     0,     0,     0,    -3,    -9,    -8,     4,     4,    -3,    -7,    -9,     0,    -3,    -2,    -1,    -2,    -6,    -5,    -4,    -5,    -2,     0,     0,     1,     1,     1,     0,    -2,     0,     3,     3,     7,     5,     0,    -3,     5,     4,     4,     8,     3,    -4,    -2,    -4,    -3,     2,     0,   -11,   -16,    -8,    -6,     1,     1,    -1,    -1,    -4,     5,    -8,     1,     8,     3,     1,    -3,    -3,    -2,     1,     4,     6,     0,     0,    -8,    -5,    -2,    -3,     2,     1,   -20,   -18,    -9,    -8,     1,    -1,     0,    -1,     0,    -3,    -2,     4,     0,    -4,    -6,    -1,     5,     6,     1,     2,    -1,     2,     1,    -1,     2,     2,     9,     4,     6,     5,   -17,    -3,     1,     1,    -1,     3,     1,     4,    -2,     2,     6,    -7,    -1,     2,     7,     3,     2,    -4,    -4,    -3,     2,     3,     0,     7,     9,     0,    -1,     4,   -12,    -9,    -2,     1,     2,     1,     4,    11,     3,     8,     3,     1,    -1,     2,     6,     3,     1,     4,     4,    -6,    -2,     1,     6,     0,     1,    -7,    -1,     2,   -11,   -14,    -4,    -3,     0,     0,     1,     4,     1,    -2,    -4,     1,     1,     1,     2,    -1,    -4,     5,     3,     2,    -4,     3,     8,     4,     6,    -4,    -3,    -2,   -14,   -14,    -2,     1,    -5,    -1,    -3,     3,     3,    -1,    -2,     0,    -2,    -4,     0,    -1,     2,     4,     2,     6,     4,     3,     2,    -2,    -3,    -3,    -4,   -16,   -17,   -16,    -6,     0,    -6,    -4,    -4,    -1,    -5,    -6,    -1,    -2,     1,    -2,     1,     4,     3,    -3,     0,     2,     8,     2,    -7,    -1,   -11,    -6,    -1,   -11,    -8,   -12,    -5,    -1,    -6,    -6,     1,    -2,    -2,    -2,     2,     0,    -4,     0,     2,     0,    -3,    -3,    -3,     0,    12,     5,     0,    -2,    -6,    -6,    -5,   -15,   -19,   -11,    -1,     0,    -4,    -8,     0,    -3,     1,    -1,    -4,    -3,    -1,     0,     2,     5,     0,    -3,    -1,     3,     7,     5,     6,     4,    -2,    -1,    -2,   -20,   -10,    -5,     0,    -1,    -2,    -6,     0,    -6,    -5,    -3,     0,     0,    -6,    -2,    -1,     5,    -1,    -2,    -4,     8,     6,     1,     5,     3,     1,    -4,    -2,    -1,   -12,   -10,    -3,    -2,     3,     0,    -3,    -6,    -1,     0,    -1,    -2,    -4,     1,     3,     1,    -1,    -4,    -2,     2,     7,     5,     9,     4,     6,    -1,    -1,     3,   -13,    -9,    -1,     0,     2,     0,     0,    -2,     8,     7,     0,     0,    -2,    -5,    -1,    -4,    -1,    -5,    -3,     2,     4,     3,     6,     3,     1,     3,     2,     6,    -9,    -5,    -3,     0,     1,     0,     3,    -1,     2,     8,     4,    -2,     0,    -1,     1,     1,    -3,    -4,    -5,     5,     7,     4,     2,     6,     5,    -1,    -4,     0,   -12,   -13,    -5,     0,     0,    -1,     6,    -1,    -1,     7,     8,    -4,    -3,    -1,     0,     3,    -2,    -7,     1,     5,     5,    -1,    -3,    -1,    -1,    -2,    -3,   -14,   -12,    -6,    -1,    -3,     1,     2,     7,     1,    -1,     6,     3,     1,     2,     4,     2,     0,    -8,    -2,     4,     4,     0,    -3,     0,     2,     1,    -3,    -5,   -12,   -13,    -3,    -3,     0,    -5,    -1,     0,     6,     6,     4,     7,     3,     3,     4,    -1,    -9,   -10,    -5,     0,    -8,    -8,    -3,    -1,    -1,    -3,     5,     1,    -8,   -11,   -11,    -6,     0,    -3,    -3,    -2,     2,     7,     4,     6,    -1,     2,     3,     3,    -9,    -8,    -5,    -5,    -9,    -9,    -5,    -3,    -3,    -7,     6,    -1,    -2,    -8,    -2,    -1,     0,    -1,     3,     1,    -2,     2,     5,     1,    -1,     0,     3,     8,     1,    -6,    -1,     1,     0,    -4,    -1,     2,    -2,     0,     2,     0,    -6,    -9,    -4,     1,    -2,    -2,     4,     0,    -2,     2,     4,    -3,     2,    -2,     8,     9,     6,    -5,    -2,     5,     1,     1,     3,    -2,     0,     0,     6,    -3,   -12,    -8,    -6,    -1,     0,     1,     1,     1,     0,     0,    -2,     1,     1,     5,     8,    10,     2,     6,     5,     6,     3,     2,     5,     0,    -1,     2,    -2,    -5,    -5,    -7,   -10,     0,     0,     0,    -3,     6,     0,    -2,     0,     6,     8,     8,     9,     1,     2,     2,     4,     5,     8,     3,    -3,    -5,     0,     1,    -1,     0,   -11,    -8,    -4,    -1,    -1,     0,     1,    -4,    -3,     6,     5,     5,     6,     7,     4,    -1,     2,     0,     4,     5,     6,     5,     4,     5,     5,     0,    -6,   -15,    -9,    -3,    -2,     0,    -1,     1,     0,    -4,    -8,     6,     4,     5,    -6,    -6,     2,     1,    -2,    -7,    -6,    -3,     3,     1,    -1,    -2,    -2,    -6,    -5,    -4,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,    -2,    -1,     0,    -2,    -4,    -5,    -6,    -3,    -5,    -6,    -4,     0,    -1,    -4,    -5,    -4,    -3,    -1,     0,     0,    -1,    -1,    -1),
		    64 => (    0,     0,    -1,     0,     1,    -1,     1,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     1,    -1,     1,     0,    -1,    -4,    -4,    -3,    -2,    -5,    -4,    -1,    -5,    -2,    -3,    -2,     0,     1,     0,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,     1,     0,     0,     1,    -1,     0,    -6,    -5,    -6,    -9,    -8,   -10,    -6,    -4,    -2,    -2,    -2,    -1,    -2,    -1,    -4,    -1,    -2,    -2,    -1,     0,    -1,     1,     0,    -1,     1,     0,    -3,    -3,    -1,    -3,    -9,   -13,    -7,     0,    -3,    -7,    -5,     0,     0,    -1,     6,     2,    -3,    -1,    -4,     0,     3,    -1,     1,     0,    -1,     0,    -1,    -2,    -4,     0,     1,    -1,    -3,    -5,     0,    -2,    -3,    -5,    -4,    -5,    -3,    -4,     0,     3,    -3,    -2,     2,     8,     3,     3,    -4,    -2,     0,     1,     0,    -2,    -2,    -5,    -1,    -5,     3,     0,     4,    -8,   -14,   -17,   -15,    -4,     6,     4,    -7,    -8,    -4,    -5,    -1,     6,     1,     3,    -4,    -1,     1,     1,    -1,    -6,    -5,    -1,     4,     2,     3,     5,    -6,   -13,   -16,   -23,   -17,    -3,     2,     5,    -2,   -11,    -4,     1,     5,     7,    -3,    -7,     2,    -3,    -1,    -6,     0,    -5,    -4,     0,    -1,     0,     5,     8,     3,    -8,   -20,   -27,    -9,     5,     3,     4,    -9,    -1,     3,     6,    13,     4,    -9,    -8,    -2,    -8,    -3,    -5,    -2,    -6,    -5,    -2,     3,     0,     2,     8,     3,    -5,   -23,   -17,    -5,     2,     6,    -1,    -8,    -6,     1,     5,     1,     4,   -10,    -1,    -6,    -6,     0,    -2,    -1,    -7,    -4,    -1,    -4,     4,     6,     6,     4,    -3,    -9,    -7,    -3,     0,     2,    -2,    -2,     0,     0,     1,     0,     5,    -4,    -3,    -4,    -2,    -1,     1,     0,    -7,    -1,     0,    -1,     3,     4,     9,     6,     1,    -8,   -11,    -2,     4,     1,     0,     1,    -1,    -4,    -4,    -3,    -1,     3,     2,    -2,    -4,     1,    -2,    -1,    -4,     1,     2,     2,     1,     6,     8,     3,    -4,    -7,    -7,    -5,    -2,    -1,     0,    -4,    -2,     1,    -1,     1,    -3,    -1,     3,    -3,    -7,     1,    -2,     1,    -9,    -3,    -1,     3,    -2,     1,     5,     3,    -1,    -1,     1,    -1,     2,     0,     1,    -1,     2,     5,    -1,     1,    -7,    -6,    -1,    -3,    -7,    -1,     0,    -2,    -6,    -7,    -5,     4,     2,    -2,     6,     2,     0,     0,     3,     1,     3,     0,     1,     4,     7,    -1,     1,     1,    -9,    -9,     0,    -4,     1,    -1,     2,    -7,    -2,     0,    -3,    -3,     2,    -5,    -3,     0,    -1,     0,    -2,     2,     6,     2,     5,     4,     1,     2,     4,    -4,   -10,    -8,     1,     8,     1,     1,    -1,     5,     1,     6,    -1,     5,    -1,     5,    -4,    -3,    -4,    -5,     0,    -3,     4,     1,     0,    -2,     1,    -7,    -1,     2,     4,    -6,     3,    10,     1,     1,     0,    -4,     4,    -1,    -6,    -5,     3,    -1,     2,    -1,    -3,    -2,    -2,    -5,     2,    -1,    -1,     0,    -4,   -11,     0,     1,    -1,     7,     9,     3,    -1,     1,     0,    -2,     1,     0,    -4,    -4,     2,     2,     1,    -2,    -3,    -4,    -3,    -6,     2,     0,    -2,     0,    -6,    -5,     4,    -1,     2,     3,    10,     8,    -3,     0,     0,    -2,    -1,    -1,    -5,    -4,     1,    -1,     0,    -5,    -8,    -8,    -2,    -4,     3,    -4,    -3,     2,    -2,    -3,    -1,    -2,     1,    -4,    -2,     0,    -2,     1,    -1,    -3,     2,    -2,    -5,    -1,     2,    -3,    -3,    -4,    -7,    -7,     0,    -1,     4,    -1,    -3,     5,    -2,    -7,    -2,     0,    -3,    -4,    -5,     0,    -2,     1,     0,     0,    -3,    -4,    -5,    -4,     3,    -2,    -2,    -5,    -3,    -8,    -3,    -2,     1,     2,    -1,     1,     2,    -1,     1,     3,     1,    -1,    -8,     0,     0,     1,     1,    -4,    -5,     0,     0,    -2,     3,     1,    -3,    -5,   -12,    -7,    -1,     5,     1,    -1,    -2,     0,     2,     0,     0,    -2,     5,     0,    -9,    -4,    -1,     1,     0,     0,    -3,    -5,     1,     1,    -1,     2,    -4,    -7,    -8,    -5,    -1,     1,     1,    -3,    -6,    -1,     6,     1,     2,     3,     7,    -3,    -4,     2,     0,    -1,     1,    -1,    -1,    -3,    -3,     0,    -1,    -2,    -1,    -3,    -9,    -2,     2,     2,    -1,    -3,    -6,     3,     4,    -3,     6,     0,    -3,    -7,     3,     1,     0,     0,    -1,    -1,     0,    -4,    -3,    -3,    -4,     1,    -1,    -3,    -4,    -3,    -1,     3,     3,     0,     0,     2,     1,     2,     2,     5,    -3,    -9,     1,    -2,     1,     0,     1,     0,     0,    -1,    -1,    -3,    -2,     2,    -2,    -4,    -4,     0,     3,    -7,    -4,    -3,     2,     2,     1,     5,     3,    -3,    -3,    -4,    -2,    -2,     1,     1,    -1,    -1,    -2,    -1,    -2,    -1,     0,     1,     1,    -4,    -2,    -2,   -14,   -15,   -15,    -8,    -1,    -3,    -8,   -11,   -10,   -13,    -1,    -4,     0,    -1,     0,     1,     1,     0,     0,     1,     0,    -2,    -5,    -5,    -3,    -2,    -5,    -5,    -4,    -5,    -2,    -5,    -8,    -6,    -5,    -6,    -6,    -7,     0,     1,     0,     0,     1),
		    65 => (   -1,     1,     0,     0,    -1,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,     1,    -1,    -1,     1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     1,     1,     0,    -2,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -2,     0,    -1,    -1,     1,     1,     0,    -1,     0,    -1,     0,     1,    -1,     1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -6,    -5,    -6,    -8,    -4,    -5,     5,     0,     2,     6,    -2,     0,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -3,    -2,    -3,    -5,     1,    -2,    -4,    -2,    -1,     2,    -4,     4,     3,     3,     8,     8,     5,    -6,    -5,     2,     8,     1,     0,     1,    -3,    -2,    -2,    -3,    -7,    -3,    -6,     5,     5,     0,     1,    -7,    -4,    -2,    -8,    -2,     4,    -3,    -3,     2,     0,    -3,    -1,     6,     5,    -5,    -1,     1,    -4,    -3,    -2,    -4,   -13,   -14,    -3,     5,     1,    -1,     3,     6,    -1,   -13,    -5,    -4,    -5,    -3,     6,     3,     3,    -3,    -3,     4,     6,    -2,    -1,    -1,     5,    -3,    -5,   -10,   -13,   -13,    -7,    -1,     4,    -2,     7,     7,    -1,    -4,    -4,     0,    -1,     2,     6,     3,     5,     0,     0,    11,    11,     4,     1,    -1,     5,    -6,    -3,    -3,   -11,   -11,    -6,     4,     1,    -1,     5,     4,    -4,     3,     6,     6,     7,     7,     8,     2,     5,    -1,    -3,     5,    11,     0,     0,    -3,    -5,    -5,    -3,   -12,   -10,    -5,    -1,    -1,    -4,    -3,     0,    -3,     0,     3,     5,     7,    11,     9,     7,    -1,     2,     4,     0,    -1,     6,     3,     1,     0,    -8,    -9,    -8,    -8,    -5,    -4,    -6,     0,    -2,    -2,    -4,    -3,    -6,    -6,    -3,     7,     3,    -1,    -5,    -4,    -1,    -2,    -3,     5,     1,     6,     1,    -1,    -1,    -1,     1,    -4,    -2,    -9,    -4,     3,    -4,     0,     1,    -4,    -8,   -19,   -20,   -15,   -12,   -17,   -14,    -5,    -7,   -15,    -7,     1,     7,     7,    -1,     0,     0,    -2,     9,     0,    -9,    -5,    -3,     0,     0,    -3,     0,    -3,    -5,   -12,   -15,   -22,   -20,   -18,   -20,   -12,   -10,   -12,    -8,    -4,     1,     6,     0,    -1,     0,     2,     4,    -4,    -7,    -3,    -2,    -1,     3,     1,     0,     6,     1,    -1,    -3,    -8,    -5,    -8,   -10,   -13,   -13,   -10,    -8,    -3,    -1,    -3,     0,    -1,     0,     4,     2,    -3,    -1,     1,    -3,    -4,    -2,    -2,    -1,     3,     4,     3,    -3,    -3,    -4,    -5,    -1,   -11,   -17,   -10,    -8,    -3,     0,    -3,     0,    -2,    -2,     5,     2,    -5,    -2,     3,     1,     2,     0,     1,     2,    -1,    -2,     1,    -3,    -2,    -3,     0,     5,    -1,    -4,    -3,    -3,    -2,    -1,    -1,     2,    -2,    -6,    -4,     2,     0,     4,    -4,    -2,     4,    -1,     0,     1,    -3,    -1,    -2,     2,    -2,     0,    -3,     2,     6,    -3,    -2,     2,     1,    -2,    -4,     1,    -1,    -4,    -3,    -2,    -1,    -4,    -7,     0,     1,     2,     3,     1,     3,     0,    -4,     0,     1,    -6,     1,    -1,    -3,    -6,    -8,     0,    -4,    -6,    -4,     0,    -1,    -5,     0,     1,    -5,    -6,    -2,    -5,    -2,     5,     4,     2,     5,    -3,    -2,    -2,    -2,    -2,     1,     3,    -3,    -5,   -10,    -1,    -4,    -1,    -6,     0,    -1,    -4,     2,     2,    -1,    -8,   -11,    -8,   -10,    -5,     3,    -1,    -1,    -7,    -6,     4,     2,     1,     0,     5,    -4,    -3,     0,     1,    -1,    -5,    -3,     1,     0,    -3,    -5,     8,     0,     0,    -5,    -6,   -14,   -13,   -14,    -5,     1,    -4,    -8,     0,     4,     1,    -2,     5,    -5,    -4,     3,     4,    -3,    -1,    -2,     0,    -2,    -2,    -3,     1,     4,     1,     1,    -2,    -7,    -1,    -6,   -10,    -1,    -2,     2,    -3,     1,     1,     4,     3,    -2,    -1,     2,    -1,    -1,    -2,     1,     0,    -1,    -6,     0,     6,     4,     1,     1,     0,     2,     3,    -1,    -1,     3,     1,     1,    -3,    -3,     1,     5,     1,    -3,     4,     3,    -2,    -1,    -4,     0,     1,     1,    -7,     6,     3,    -4,    -2,    -3,     2,     8,     6,     5,     1,    -4,     2,    -3,    -1,     2,    -1,     0,     1,     0,    -1,     7,    -1,    -2,    -1,    -1,     0,     1,     3,     8,     7,     4,     5,     1,     1,    -5,     2,     4,     2,     0,    -1,     1,    -4,    -2,    -1,     1,     1,     0,     2,     8,    -2,    -5,     1,    -1,     1,     1,    -4,     2,    -2,    -2,     0,     0,    -2,     1,     1,    -2,    -2,    -1,     0,     0,    -4,    -2,     3,    -2,    -4,     2,    10,     2,     4,    -6,    -3,    -1,    -1,    -1,    -1,     9,    -7,    -7,    -3,    -4,    -7,     1,    -4,    -3,     1,     5,    -2,    -1,   -11,     2,     2,     1,     3,     8,    13,     6,     4,     0,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -6,    -2,     5,     5,     3,   -11,   -12,   -10,   -11,    -5,     3,    -4,     3,     3,    -1,    -1,     0,    -1,    -1,     1,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     0,     1,     2,    -3,     0,     0,     0,    -2,    -1,     1,    -1,    -3,    -1,    -1,     0,     1,     0),
		    66 => (    0,     1,     0,    -1,     1,     1,     0,     0,     1,    -1,     0,     0,     4,     5,     1,    -1,     0,     0,    -1,    -1,     0,     1,     0,     1,     1,    -1,     0,     0,     0,     1,    -1,    -1,     0,     0,     2,     2,     1,     0,     6,     1,     2,     6,    -3,    -2,    -1,     1,     3,     5,     6,     5,     4,     4,     0,     1,     0,     0,     0,    -1,     0,    -1,     2,     4,     3,    -1,     1,     5,     4,     4,     3,     4,     4,    -2,     4,     4,     5,     8,     7,     4,    12,     8,     6,     5,     0,     0,     1,     1,    -7,     4,    -1,     7,     8,     7,    10,    10,    12,    12,    15,    10,    13,     9,     2,     1,     1,     1,    -4,    -5,    -3,     0,     5,   -10,    -8,     0,     1,    -1,    -5,     0,     4,     6,     7,    10,     5,    10,     9,     5,     9,     1,    10,     8,     2,     4,     2,     5,     6,     3,    -2,    -3,    -3,    -7,    -3,     7,    -1,    -1,    -3,    -6,     9,     4,     5,     6,     4,     4,     8,     2,    -5,     4,     9,     4,     1,     6,     1,    -2,     2,    -5,    -1,     1,     7,     3,     7,     2,     1,     0,     0,     1,     7,     2,     7,     4,    -1,     3,    -2,    -4,     2,     2,     2,     1,     1,     0,    -8,     2,    -1,    -5,    -5,    -4,    -1,     3,     6,     9,     0,    -1,     0,    -2,     7,     5,     3,     2,     1,    -2,    -4,    -2,    -6,    -8,     3,    -3,    -1,    -3,    -2,     1,    -2,    -1,    -2,    -2,     3,     1,     5,     6,    -1,    -3,    -4,   -13,     8,     3,     1,    -3,     0,     4,    -3,    -4,    -2,    -5,     0,    -6,   -11,    -5,    -3,    -1,     3,     3,    -2,    -5,    -5,   -11,    -1,    -8,     0,    -1,    -5,    -7,     6,    -1,    -4,    -3,     1,    -2,    -4,    -5,    -7,    -8,     0,     0,    -4,   -10,    -2,    -2,    -1,     5,    -1,    -1,    -7,   -13,    -8,    -7,    -1,    -1,    -5,    -4,     2,     1,    -4,    -5,    -1,    -3,    -2,    -7,    -8,    -4,     1,    -3,    -9,    -5,    -8,    -6,     1,     1,    -6,    -5,    -9,   -10,    -8,    -8,     0,    -1,    -1,    -8,     2,     1,     0,    -1,    -4,    -1,    -3,    -6,     1,    -1,    -1,    -5,    -5,    -4,    -5,    -3,    -2,     1,    -5,    -1,    -4,    -8,    -9,    -6,     1,    -1,    -4,    -8,    -1,     2,     6,     2,    -2,     2,     0,     1,    -2,     3,    -4,    -3,    -7,    -4,    -6,    -4,     3,     2,    -4,     4,     5,    -1,   -12,    -6,     0,     1,    -3,    -7,    -3,     3,    -1,    -3,    -3,     5,     6,     4,     4,     2,     3,     1,    -2,    -8,    -2,     3,     4,     4,    -3,     4,     3,    -4,   -12,     0,     0,    -1,    -1,    -6,    -9,     3,    -4,    -6,     2,     2,     6,     6,     7,     4,     1,    -5,    -1,    -4,     2,     2,     1,     3,     3,    -3,    -2,     6,   -10,    -2,     0,     0,    -4,    -4,   -10,    -4,    -3,    -1,    -3,    -1,     2,     3,     0,     8,     5,    -3,    -3,    -8,     1,     4,    -1,     1,    -6,     1,     0,     6,    -4,   -12,     1,     0,    -6,    -5,    -2,     2,     2,     3,    -3,     3,     3,     1,    -2,    -4,    -3,    -3,    -3,    -4,     5,     6,    -2,    -2,     2,     0,    -2,     4,    -6,   -10,    -1,     0,    -7,    -7,    -4,     6,     0,     2,    -1,    -4,    -3,    -1,    -2,    -4,     1,     2,     2,     4,     3,     4,     3,    -2,    -1,    -3,    -1,     4,    -6,   -14,     1,    -1,    -6,   -10,    -2,    -1,    -4,     1,    -1,     1,     4,    -7,     0,    -1,     0,    -5,     0,     4,    10,     8,     1,    -3,     0,     2,     1,     6,     0,    -6,     1,     0,    -8,    -8,     1,     3,     3,    -1,     1,     0,     8,     8,     4,     2,     1,     2,     0,     6,     0,     8,    -1,    -1,    -1,    -3,    -7,     2,    -4,     0,     0,     0,    -7,   -11,     0,     0,     0,     3,     1,     2,     7,     7,     6,    -4,     2,     2,     1,     4,     4,     4,     4,     0,    -1,    -8,    -9,    -3,    -3,     0,    -1,    -1,    -9,   -10,    -7,    -8,    -2,     6,     7,     0,     4,     0,    10,     5,     2,     1,     8,     5,     5,     3,     2,    -3,    -2,    -8,    -4,     0,    -1,    -1,     0,     1,    -7,    -7,   -13,   -17,   -22,     0,     0,     4,     2,     1,     0,     0,     1,     6,     7,    10,     6,     1,     2,     2,    -7,    -6,   -15,    -4,    -2,    -1,     0,     1,     1,    -8,   -10,   -12,   -11,    -1,    -3,     0,    -4,     1,     5,    -1,     2,     5,     0,    -4,     1,     0,     1,     3,    -8,   -10,   -10,    -7,    -8,     1,    -1,     0,    -1,    -1,    -3,    -4,    -6,   -11,   -15,   -19,   -13,   -17,    -8,    -8,    -5,     1,     3,     4,     9,   -13,    -2,    -7,    -6,    -5,    -4,    -3,    -1,     0,     1,     1,     0,    -1,    -1,    -2,    -4,    -4,    -3,    -4,    -5,     2,     4,    -2,    -2,    -4,    -6,    -6,    -3,   -10,    -9,    -2,    -5,    -5,    -4,     1,    -1,     1,     0,     1,     0,     0,    -1,    -2,     1,    -1,     0,    -1,    -1,    -2,    -1,     0,    -1,    -2,     0,    -1,     0,    -1,    -1,     1,    -1,    -1,     1,     1,     1,     1,     0,     1,    -1,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,     1,     1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     1,    -1,     0,     0,     0),
		    67 => (   -1,    -1,     1,    -1,     0,     0,     0,     1,    -1,    -1,     1,     1,     1,     0,     0,     0,     1,     1,     1,     1,     0,    -1,     1,     1,     0,     1,    -1,    -1,     1,    -1,     0,     0,     1,     0,     1,    -1,     1,     0,     0,    -1,    -1,    -2,    -2,    -5,    -5,    -3,     0,     0,     0,    -1,     0,    -1,     1,     1,     0,     1,    -1,    -1,     1,    -1,     0,     0,    -1,    -1,    -2,     1,    -1,    -4,    -7,    -3,    -3,    -3,     1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -1,     1,    -1,     0,    -2,    -4,    -4,    -7,    -3,    -1,    -3,    -5,    -8,    -9,    -6,    -6,    -4,    -3,    -1,     0,    -1,     1,    -3,    -1,    -2,    -2,     1,     0,     1,     0,     0,    -1,    -3,    -1,    -5,    -5,    -8,    -9,   -13,     1,     1,     0,    -2,    -6,   -15,   -11,    -8,    -9,    -6,     1,    -4,    -5,    -6,    -4,    -1,    -1,    -1,    -1,     0,    -3,    -5,    -2,   -10,     0,    10,     2,    -2,     0,     3,    -1,     3,     1,     1,     0,     7,     0,    -5,    -3,    -2,    -4,    -8,    -1,    -2,    -1,     0,     0,     3,    -2,    -2,    -2,    -6,     3,     4,     7,     3,    -1,    -2,    -2,    -2,     3,     1,     0,     5,     2,    -9,    -4,     0,    -5,    -5,    -4,    -4,    -2,     1,     3,     4,     0,     2,     0,     3,     2,     4,     3,    -1,    -3,    -5,    -5,    -6,     0,     5,     5,     4,     6,     9,     2,    -4,    -4,    -7,    -4,    -3,    -2,    -5,     2,    10,     1,     4,     3,     2,     6,     6,     1,    -1,    -2,    -2,    -4,     1,     6,     1,     1,     2,     3,     6,     3,    -1,    -9,    -6,    -1,    -3,    -2,     2,     2,     2,     5,     4,    -7,    -2,     0,     2,     0,     2,    -4,    -2,     2,     0,    -1,     2,     5,    -2,    -1,     3,    -4,    -3,    -5,    -3,    -1,    -5,     2,     1,     1,    -1,     1,     7,    -2,    -2,     1,    -3,     2,     2,    -4,    -8,     2,    -1,     1,     1,    -1,     0,     1,    -2,    -6,    -2,    -5,    -5,    -1,    -3,     0,     2,     2,    -1,    -5,     0,     1,    -2,     4,     2,    -3,     1,     0,    -8,    -5,     0,     7,    -1,     0,     0,    -1,    -5,    -3,    -5,   -10,    -5,    -6,    -5,     2,     1,     1,    -4,    -1,    -4,    -1,    -4,     4,    -1,    -5,    -3,    -9,   -10,    -7,    -4,     5,    -2,    -6,    -2,    -9,    -5,    -5,    -9,    -9,   -10,    -3,    -3,     1,    -1,     3,     4,    -2,    -1,    -1,    -3,     0,     1,    -4,    -5,    -9,   -17,   -11,    -6,    -1,    -3,     0,    -3,    -8,    -7,    -7,    -8,   -11,   -10,    -1,    -6,    -3,     0,     4,     1,     4,     0,     3,    -7,    -3,    -7,   -10,   -18,   -14,    -9,    -7,    -5,     0,    -5,     2,     4,     1,    -3,     2,    -6,    -7,    -3,    -1,    -5,    -2,     1,     0,     0,     3,     3,    -2,    -5,   -13,    -8,    -7,   -10,     1,    -2,    -1,    -6,     0,    -1,     5,     5,     1,     3,     3,    -1,     1,     1,     2,    -2,    -2,     0,     0,     0,    -3,    -2,     0,    -8,    -4,     7,    -2,    -2,     6,     2,     0,    -1,     5,     2,     1,     5,    -3,    -1,    -5,    -3,    -1,    -1,    -8,    -4,    -1,     1,     0,    -4,    -3,    -5,    -9,    -4,    -3,    -2,     0,    -5,     1,    -1,     0,    -2,     2,     2,     5,     3,     0,    -9,    -9,    -8,    -6,    -2,   -12,    -7,    -8,     2,     0,     2,    -4,    -4,    -1,    -3,     0,    -3,     2,     0,     1,    -5,     4,     2,     6,    -1,     7,    -4,     2,     4,     1,    -6,    -8,    -5,    -9,     1,    -6,     0,     1,     0,    -1,    -1,    -8,    -3,    -3,     3,    -2,    -2,    -6,    -3,    -3,     6,     9,    -4,    -3,    -3,     3,     4,     5,    -3,    -1,     2,    -4,    -5,    -4,     0,     3,    -2,     0,    -1,    -7,    -5,     0,     2,     3,    -1,   -13,    -4,    -2,     3,     2,    -4,    -7,    -3,    -1,     4,     0,    -3,   -10,    -5,    -3,    -5,     1,    -1,     1,    -2,    -3,    -2,    -7,   -10,    -9,     2,    -3,    -4,    -7,    -1,     0,     4,     1,     5,    -7,    -3,    -5,    -3,     1,    -4,   -12,    -7,    -7,     0,     0,    -2,     1,    -1,    -1,    -2,    -6,    -8,    -8,    -4,    -6,    -3,    -7,    -4,     4,     1,     4,     1,     2,    -5,    -2,    -3,   -10,   -16,   -11,    -7,    -4,    -6,     0,     0,     1,    -2,    -4,    -9,    -9,    -8,   -12,   -10,   -14,   -10,    -8,    -5,    -2,    -2,     0,    -2,    -7,   -11,    -8,    -7,    -7,    -7,    -6,     2,    -4,    -6,    -1,    -1,    -1,     1,     0,    -3,    -9,   -10,   -10,   -15,   -14,   -11,    -7,    -2,     0,     2,     5,    -1,    -2,   -10,    -6,    -1,    -3,    -1,    -5,    -3,    -3,    -1,     0,    -1,     0,    -6,     0,     1,    -4,    -6,    -8,    -8,   -13,    -8,     2,    -4,    -3,    -1,     7,     1,     2,     0,     3,     5,     3,    -2,    -4,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -3,    -3,    -1,     4,     2,     2,    -3,    -2,     3,     5,     3,     1,     0,     2,    14,    12,     7,     2,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     0,     1,     2,     0,    -1,    -2,     0,     5,     7,     4,     3,     3,     1,     6,     5,     8,    12,     8,     4,    -1,    -2,     1,     0,    -1,    -1,    -1),
		    68 => (    1,     1,     1,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     1,    -1,    -1,    -1,     1,     1,     1,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -5,    -5,     0,     0,    -1,    -1,    -1,     1,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     1,    -1,    -3,    -1,     0,    -1,     1,    -1,    -3,     0,     0,     0,    -1,    -3,    -1,    -2,     0,    -1,     1,     1,    -1,    -1,     0,     0,    -1,    -2,    -1,    -3,    -2,    -2,     0,     0,    -1,     0,    -4,    -3,    -1,     0,     2,    -1,    -3,     0,     1,     1,    -1,     0,    -2,     1,     1,    -1,     0,    -2,    -1,    -1,    -4,    -4,     1,     0,    -1,     4,     4,    -3,     0,    -6,    -5,    -1,     2,     0,     2,    -2,    -3,     0,    -2,     1,     0,     0,    -1,    -1,     0,    -2,    -6,    -7,     0,    -1,     0,     0,    -3,    -2,    -3,    -3,     1,    -2,    -4,    -2,    -2,    -3,    -1,    -2,    -3,    -2,    -1,     3,     0,    -2,    -1,     0,    -3,    -5,    -1,     1,    -1,     3,    -1,    -2,    -4,    -6,    -2,    -6,    -3,     0,     0,     0,    -1,    -2,    -2,    -4,    -1,    -1,    -1,    -2,    -1,     0,     1,    -1,    -2,     0,     1,     6,     1,     2,     1,    -1,    -1,    -4,     1,     0,     1,     2,     2,     1,     0,     1,    -4,    -1,     1,     0,     2,     0,     0,    -1,     0,    -3,    -1,     5,     7,     8,     3,    -1,    -5,    -3,    -1,     2,     1,     1,     0,    -3,    -4,    -2,    -2,    -2,     0,     1,     1,    -1,    -1,     1,    -2,     0,     0,    -3,    -4,     4,     6,     7,     3,    -3,    -6,    -4,     2,    -4,    -4,    -2,    -3,    -6,    -5,    -1,    -2,     3,     3,     3,     1,     0,     0,     3,    -2,    -1,    -1,    -2,    -4,     2,     2,     6,     5,     3,    -3,     1,     3,    -1,     0,    -2,    -2,    -3,    -3,     0,    -2,     0,     1,     0,    -2,    -3,     0,    -3,    -2,    -2,     0,    -1,    -5,    -3,    -2,     0,     5,     6,     4,     6,     4,     1,    -1,    -2,    -3,    -2,    -2,    -2,    -5,     0,    -1,    -1,     1,    -1,    -3,    -2,     0,    -5,     0,     0,    -3,    -7,    -5,    -1,     1,    -2,     2,     1,     4,     0,     0,    -5,    -5,     0,     0,    -1,    -1,    -3,    -3,     3,     1,    -1,    -2,    -3,    -3,    -6,     0,    -2,    -5,    -8,    -3,    -5,    -5,    -5,    -5,    -4,    -2,     1,     1,    -3,     1,     2,     0,    -3,    -3,    -6,    -4,    -1,    -1,    -1,    -3,    -5,    -3,     2,    -2,    -1,     1,    -8,    -3,    -3,    -4,    -6,    -6,    -9,    -4,    -6,    -3,     0,    -1,    -5,    -5,    -1,     0,    -2,    -5,    -2,    -1,    -1,    -4,    -2,    -9,    -1,     0,     1,    -2,     2,     0,    -2,    -3,    -6,    -3,    -5,    -4,    -2,    -3,     0,     0,    -2,     0,    -2,     0,    -3,     0,    -3,    -3,    -3,    -3,     2,    -3,    -4,     1,    -2,     0,     2,     0,    -2,    -4,    -2,    -1,    -4,     0,     1,     0,    -2,    -5,    -5,     2,     2,    -3,    -2,    -1,     0,     0,    -2,    -2,     1,    -4,    -3,     1,     0,     0,     3,    -1,    -3,    -3,    -2,    -3,    -3,     3,     4,     0,    -4,    -4,    -6,    -3,     2,     0,    -3,    -2,     1,     2,    -3,    -2,    -2,    -1,    -2,     0,    -1,    -1,     0,    -2,    -2,    -3,    -2,    -4,    -3,     1,     0,     2,     0,    -5,    -4,    -4,     3,     1,    -1,    -5,    -2,     4,    -1,    -2,     1,     0,    -4,     1,     1,    -1,    -1,    -3,    -1,    -1,    -2,    -7,     0,     3,     3,    -1,     0,    -3,    -4,    -4,    -1,     4,     1,    -1,     1,     2,     3,     0,     1,    -3,    -3,    -1,     0,    -2,    -2,    -2,    -2,    -1,    -2,    -5,    -1,     1,     4,     2,    -4,    -6,    -4,    -5,    -1,     2,     0,     0,     0,     4,     1,    -1,     0,    -3,     0,    -2,    -2,    -1,    -3,    -1,    -1,    -4,    -3,    -3,    -2,    -2,     1,     2,    -1,    -3,    -3,    -5,     1,     2,     1,     1,     1,     4,     0,    -1,    -2,    -2,     0,    -4,    -2,    -2,    -2,    -2,    -3,    -2,    -2,    -3,    -3,    -1,    -1,    -2,    -1,    -2,    -2,    -3,     2,    -1,    -1,     0,     3,     1,    -1,    -4,    -2,    -1,     0,     1,     1,     0,    -2,    -2,    -4,    -4,    -3,    -1,    -3,     0,    -4,    -2,     2,    -2,     0,     2,     0,    -1,     0,     2,     4,     1,    -2,     0,     0,    -5,     0,    -1,     1,    -1,     0,    -1,    -3,    -2,     1,    -2,    -1,     0,    -4,    -3,    -4,     1,     3,     3,    -3,    -5,    -3,     0,    -3,    -4,    -1,    -1,    -2,    -1,     1,     1,    -1,    -2,    -2,    -2,    -2,    -3,    -3,    -2,     0,     3,    -2,    -3,    -2,     0,     1,     0,    -1,    -2,    -2,    -4,    -3,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,    -1,     0,    -2,    -2,    -3,    -2,    -4,    -3,    -3,    -3,    -3,    -5,    -4,    -1,     0,     0,    -5,    -6,     0,    -4,     0,     1,     1,     0,     0,     0,     1,     1,     0,     0,     1,     0,    -1,    -1,    -2,    -2,    -1,     0,    -2,    -1,    -1,    -2,    -2,    -3,    -1,     0,    -1,    -1,    -1,     0,     1,    -1,     0),
		    69 => (   -1,    -1,     1,     1,     1,     1,     0,     1,    -1,     1,     1,     1,     0,     0,     0,     1,    -1,    -1,     1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,     0,    -1,    -2,    -3,    -2,    -2,    -3,    -4,    -6,    -3,    -7,    -6,    -6,    -3,     0,     1,    -1,    -3,     0,     1,    -1,    -1,    -1,    -1,     0,    -1,    -5,    -5,    -1,    -1,    -5,    -7,    -3,    -3,    -5,     0,     0,   -14,    -8,    -7,    -5,    -8,    -6,   -11,   -12,    -9,    -7,    -4,    -2,     1,     0,     0,     0,    -1,    -6,    -8,    -7,    -4,    -7,   -16,   -20,   -27,   -24,   -16,   -21,   -19,   -21,   -27,   -24,    -7,   -10,   -17,   -15,   -12,    -7,    -6,    -4,     1,     1,     1,    -1,    -3,    -5,    -9,   -11,   -16,   -11,   -12,   -13,    -8,    -2,     1,    -1,    -4,    -4,    -4,    -8,   -14,   -28,   -18,   -15,   -15,    -8,    -7,   -11,    -8,     1,    -1,     0,    -3,    -5,    -4,    -6,    -7,    -4,   -10,     2,     2,     1,     4,     8,     3,     3,     7,     7,    -1,    -4,    -8,    -3,   -16,    -7,   -10,   -11,    -7,    -2,    -1,     1,    -3,   -11,    -8,   -10,    -5,    -3,     0,     5,     5,    -3,    -2,     7,     3,     8,    12,     8,     2,     3,    -2,    -1,    -2,     2,     0,    -3,    -8,    -9,     0,    -4,    -7,    -9,    -6,   -10,    -1,    -1,    -2,     2,     2,    -1,     4,     9,     8,     7,    15,     9,     0,     3,     4,     0,     2,     2,     0,     1,    -9,    -7,    -6,    -8,    -6,    -7,    -8,    -1,     3,    -1,     0,     2,     1,     1,     6,     5,     8,    12,    10,     7,     6,     7,     1,     3,     2,     5,     5,     0,    -8,    -5,    -1,    -6,    -8,    -9,     5,     2,     5,     2,     3,     5,     1,    -2,     2,     7,     7,     4,     3,     2,     2,     2,     6,     0,     0,    -2,    -3,    -9,   -11,    -7,    -1,    -4,   -12,    -6,     5,     5,     0,     1,    -1,    -1,     0,     0,     4,     3,     2,    -5,     0,    -3,     0,     0,     2,    -5,    -3,    -3,    -7,     5,   -11,    -5,    -1,   -18,     0,    -4,     2,     6,     3,    -2,    -5,    -1,    -2,    -4,     0,    -7,    -6,    -6,     0,     2,    -5,    -2,     4,    -3,    -8,    -5,    -7,    -1,    -9,    -4,     0,    -2,    -1,    -4,     4,     3,     2,    -3,    -6,    -6,    -2,     0,    -5,    -7,    -3,    -5,    -3,     1,    -4,    -6,     1,    -4,    -4,    -1,    -8,   -13,    -8,    -6,    -1,    -4,    -6,    -4,     2,    -2,     2,     1,     0,    -4,    -1,    -4,     0,    -2,    -3,    -6,     1,     0,    -2,    -3,    -4,     0,    -5,    -5,    -3,   -10,    -6,    -2,    -2,    -3,    -4,    -1,     3,    -1,    -1,     2,     0,    -1,     0,    -2,     3,    -6,    -4,     2,     1,     0,     3,     2,    -1,    -4,    -5,   -11,    -5,   -12,    -7,     0,     0,    -1,    -8,    -3,     1,     1,     3,     1,     4,     3,    -4,    -6,    -5,    -2,     3,     2,     5,     2,     4,     6,     8,     3,     1,    -8,    -5,   -11,    -2,    -7,     1,    -2,    -6,    -4,     0,     5,     4,    -1,     2,     1,    -1,    -7,    -7,    -2,     5,     4,     1,     5,    -2,     4,     6,     1,     0,    -6,    -2,   -14,    -8,    -8,     0,     0,    -8,     1,    -5,     1,    -4,    -2,     0,     2,    -2,    -4,    -1,    -3,     4,     1,     1,     2,    -3,     0,     2,    -3,   -11,   -13,    -4,   -17,   -10,    -6,     3,     0,   -10,     7,    -5,    -4,    -1,     0,    -7,    -3,    -4,    -6,    -9,    -1,    -4,    -2,     3,     2,    -7,     1,     1,    -6,    -4,    -4,    -6,   -13,    -9,    -4,     1,    -2,    -8,     3,    -1,    -4,    -6,    -2,    -8,    -3,     0,    -2,    -1,    -4,     0,    -4,     2,    -2,    -2,     1,    -1,    -5,     0,     5,    -3,    -9,    -6,    -3,     1,    -3,   -16,     1,    -6,     2,    -1,   -10,    -3,    -5,    -3,    -3,    -6,    -5,    -3,    -5,     1,     1,    -3,     1,    -4,    -6,     0,     9,     8,     4,    -5,     0,     1,    -1,   -13,     2,    -2,     3,     2,    -2,    -3,    -7,     2,    -1,    -5,    -3,    -1,    -3,     5,     4,    -1,    -5,    -7,    -1,     2,     6,     6,    -1,   -13,     1,     0,     0,   -10,     4,    -4,     0,    -3,    -4,     0,    -3,     0,    -6,     2,    -3,     5,     1,     6,     5,     1,    -5,    -2,     1,     8,     8,     6,    -9,    -9,     0,     0,     1,    -1,     2,    -3,     1,     1,     7,     3,     0,    -3,    -1,     1,     3,     6,     5,     4,     3,     2,     0,    -2,    -1,     3,     6,    10,    -4,    -6,     1,    -1,     0,    -5,    -7,    -2,     3,     9,    11,     7,     5,     2,     4,     1,     3,    -6,    -4,    -4,     3,    11,     5,     6,     1,    -4,     1,     2,    -4,     0,     0,     0,     0,     5,    -6,    -1,     4,     7,    10,     7,     6,     0,     3,    -2,    -4,     3,    -2,    -1,     7,     6,     3,     5,    -2,    -1,    -4,     0,     0,    -2,     1,     0,    -1,     0,     4,     0,     3,     5,     9,    -2,     2,     0,    -3,     3,    -2,     7,     6,     3,     0,     3,    -1,     9,     2,    -3,     6,     2,     0,     1,     0,     1,     1,    -1,     1,     0,    -4,     2,     1,     2,     0,     2,     4,     4,     3,     3,     1,     3,    -5,     0,     2,    -3,    -7,    -5,    -5,     1,    -1,     1,    -1),
		    70 => (    0,    -1,    -1,     0,     1,    -1,    -1,     0,     0,     1,     0,    -1,     0,     0,    -1,    -1,     1,    -1,     0,     0,    -1,     1,     0,    -1,     1,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     1,     2,    -1,     0,    -1,     1,     1,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,    -2,    -2,     0,    -2,    -3,    -5,    -2,     1,    -2,    -4,    -2,    -1,     0,    -1,     0,    -1,    -1,     1,    -1,     0,    -1,     1,    -1,    -1,    -1,     2,    -2,    -3,    -3,   -10,    -5,    -3,     1,     4,     2,    -5,    -1,    -1,     0,     1,    -2,    -5,    -5,    -2,     1,     0,     0,    -1,     1,     1,     1,     1,    -2,    -9,    -3,    -1,    -3,    -1,    -2,     5,     7,     8,     4,     2,    -7,    -8,    -2,     1,    -6,    -7,    -4,    -2,    -2,    -4,    -2,     0,    -1,    -1,    -3,    -1,    -2,    -6,    -2,     0,     1,     0,     1,     2,     8,     2,     2,     4,    -2,    -7,    -6,     4,    -4,    -7,     1,     2,     0,    -6,    -5,    -3,     1,    -1,    -1,    -2,     2,     2,     3,     3,     3,     1,     0,     7,     1,    -1,     1,     0,     5,     3,    -4,     0,    -3,    -2,    -1,    -2,    -1,    -9,    -4,    -2,     0,    -1,    -2,    -5,     1,     3,     5,     4,     1,     3,     1,     4,    -1,     1,     6,     3,     7,     2,     2,     3,     4,     2,    -5,    -2,    -2,    -2,    -5,    -4,     1,    -1,     5,    -4,     3,     0,     3,    -3,    -1,     5,     4,    -1,    -3,     5,     4,    -1,    -3,    -4,     5,     0,     2,     4,    -1,     0,    -4,    -3,    -7,    -3,     1,     0,     6,    -1,    -1,    -3,    -5,    -5,     4,     4,     5,    -1,    -2,     5,    -1,     1,    -2,    -1,    -2,     6,    -1,    -3,    -2,    -3,    -5,    -5,    -6,     1,     0,     1,     6,     1,    -4,    -1,    -4,    -5,     3,     3,    -1,     0,     0,    -5,    -1,     3,     0,    -3,    -5,    -4,    -6,    -3,    -3,     3,    -1,    -2,    -5,     0,     1,     6,     0,    -3,    -4,    -1,    -2,    -3,    -1,    -1,     3,    -3,    -9,   -14,   -11,    -2,    -3,    -5,    -5,    -5,    -2,    -3,    -2,    -2,     2,    -3,    -2,    -3,     0,     0,    -1,    -2,    -4,    -6,    -2,    -5,    -3,    -1,    -4,     0,   -12,   -14,   -16,    -7,     4,    -3,    -4,    -2,     1,     1,    -1,    -3,    -6,    -4,    -4,    -3,     0,     1,     2,     4,    -2,     0,     1,    -3,    -2,     1,     2,     0,    -8,   -14,    -6,    -3,     0,     2,    -2,    -3,     2,     4,    -1,    -2,    -5,    -4,    -6,    -1,     0,     1,    -1,     4,     2,     0,    -3,    -3,    -5,     3,     7,     0,    -8,    -6,    -5,    -6,    -7,    -1,     2,     0,     1,     4,     1,    -2,    -3,     0,    -5,    -1,     0,     0,    -2,     2,     4,     1,    -8,    -3,     1,     6,     9,     0,    -4,    -7,    -2,    -6,   -12,    -1,    -1,    -1,     4,     3,     4,    -3,    -4,     4,    -4,    -5,    -1,     0,    -1,     2,     2,    -4,    -6,    -3,    -1,     2,     4,     4,    -6,    -3,    -4,    -3,   -15,    -1,    -2,    -2,     4,    -2,     3,    -3,    -6,    -3,   -10,    -3,     0,    -1,    -3,     2,     1,    -3,    -5,    -2,     0,     2,     4,     1,    -1,    -8,   -11,   -19,    -8,     0,    -5,    -2,     2,    -3,     0,     0,    -2,    -4,    -8,     0,     0,     0,    -2,    -1,    -1,    -5,    -6,    -4,    -3,     2,     5,     1,    -3,    -7,   -14,   -15,   -10,    -6,     6,     0,     4,    -2,    -1,     0,    -3,    -4,    -5,    -2,    -1,     1,    -2,    -1,    -1,    -2,    -6,    -4,    -2,     7,     2,    -2,     1,    -3,    -6,    -5,    -2,    -2,     0,    -1,     2,    -1,    -4,     1,     1,   -10,    -2,     0,     1,     1,    -1,    -3,     2,     5,    -7,    -4,    -4,     0,     3,     6,    -4,    -2,     5,     0,    -2,    -1,     1,    -3,     0,     2,    -4,     3,     1,    -7,     3,     1,    -1,     1,     0,    -1,    -1,     0,    -9,    -2,    -5,    -3,     1,     4,     5,     5,     3,     4,    -4,    -3,    -2,     1,     4,     1,     1,     2,     2,    -1,     2,     3,     0,     0,     0,    -2,    -3,    -1,    -4,    -2,    -2,     0,    -3,     4,    -1,     3,     4,    -1,     2,    -2,     0,     3,     4,     2,     1,     2,    -1,     0,     2,     2,     0,     1,    -1,    -3,     0,    -1,    -6,    -8,    -3,     3,    -1,    -2,    -1,     5,     3,     6,     8,     8,     2,    -5,    -4,    -2,    -1,    -3,     1,    -5,    -2,     0,     0,    -1,    -2,     1,     3,    -2,    -4,    -3,    -6,    -3,    -2,    -3,    -2,    -2,    -3,     0,    -1,     1,    -1,    -4,    -2,     0,     0,    -2,    -2,    -1,     1,     0,     1,     1,     1,    -1,    -1,     0,    -3,     0,    -1,    -1,    -1,    -2,    -1,    -2,     0,    -9,    -7,    -7,    -4,    -5,    -6,    -4,    -4,    -1,    -1,     1,     0,     0,     0,    -1,     1,     0,     0,    -3,    -5,    -1,    -1,     0,    -2,    -2,    -1,    -5,    -6,    -5,    -4,    -7,    -8,    -1,    -7,    -5,    -1,    -1,    -1,    -1,     0,     1,     0,     1,    -1,     0,     1,     1,    -1,     1,    -1,    -1,    -1,    -1,     0,    -3,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,     0),
		    71 => (   -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     1,     0,    -1,     1,     1,     1,     0,     1,     0,    -1,     0,    -1,    -1,    -1,     1,    -1,     1,    -1,    -1,     0,     1,     1,     1,     1,     1,    -1,     0,    -1,     1,    -1,    -1,     3,     1,     2,     0,    -2,    -1,    -1,     1,    -1,    -1,     0,     1,    -1,     0,    -1,     1,    -1,    -1,    -1,     1,     1,     1,    -4,    -4,    -2,    -2,    -6,    -3,    -4,     0,     6,    -1,    -2,    -1,    -4,    -9,    -6,    -4,    -2,    -2,     0,    -1,     1,    -1,     7,     1,     0,    -2,    -2,    -1,    -4,    -6,    -7,    -8,    -1,     1,    -8,    -2,     4,     4,     5,     4,     5,     5,    -2,     0,    -1,     0,     0,     1,     1,    -1,     5,     6,     1,     2,     1,    -1,     2,     0,     2,    -1,     0,     2,    -5,    -6,    -1,     2,     3,     5,    -3,     4,    -2,     1,    -1,    -4,    -5,    -2,     1,     1,     3,     1,     2,     3,     0,    -1,    -4,    -3,    -3,     0,     5,     0,     4,     4,     2,    -6,    -1,     3,     2,     2,     2,     1,    -1,    -4,    -1,    -2,     0,     0,    -4,    -4,    -1,     2,     1,    -1,   -11,   -16,    -7,     1,    -2,    -3,    -2,    -1,     1,    -6,     4,    -1,     1,     4,     2,     1,    -1,     0,    -3,    -1,     1,    -1,    -5,    -4,    -5,     2,     2,    -5,   -10,    -5,     0,    -4,    -1,    -4,    -1,    -5,    -3,    -3,     2,     1,     3,     6,     2,    -1,    -2,     0,    -5,    -1,     0,    -2,    -6,    -5,    -7,    -2,     7,     1,    -8,    -4,     1,    -2,     5,     5,     0,    -2,    -3,    -4,    -6,    -7,     0,     3,     4,    -3,    -4,    -1,    -5,     0,     0,     0,    -3,    -5,    -4,    -1,     1,     4,     3,     1,    -5,    -3,    -2,     3,     1,     0,    -4,    -4,    -7,   -10,    -4,    -1,     2,     5,    -2,     6,     5,    -2,    -1,    -2,    -4,    -2,    -3,    -3,    -5,    -3,     4,    -2,    -6,    -2,     1,     5,     1,    -5,    -2,     1,    -5,    -3,    -7,    -8,     4,     4,    -3,     5,     4,     4,     0,     0,    -2,    -1,    -3,    -3,    -5,    -5,    -7,    -8,    -7,     0,     1,     0,    -2,    -5,    -4,     0,    -6,    -5,    -3,    -4,     3,     4,    -2,     5,     3,     7,     1,     1,    -2,    -3,     0,    -1,     0,     0,    -5,    -3,    -1,     1,     4,     4,    -1,    -2,     1,     6,    -7,    -7,    -2,    -2,    -3,    -1,     0,     6,     8,     9,    -1,     1,     0,     0,    -1,     3,     2,     1,     4,     5,    -2,    -2,    -1,    -7,     0,    -1,     1,     1,    -9,    -9,    -6,    -5,    -6,    -9,    -5,     8,     6,    -1,     1,    -1,     0,     2,    -2,     3,     3,    -2,     9,     8,     3,    -5,    -8,    -6,     1,    -1,     5,     0,    -4,    -7,    -3,    -4,    -4,    -2,    -1,    -1,     1,     0,     0,    -1,     0,    -2,    -3,    -2,    -5,     3,     4,     9,     0,    -3,    -2,    -1,    -1,    -1,     3,    -1,    -2,    -6,    -5,    -7,    -5,    -5,    -6,    -1,     0,    -2,     0,     0,     0,    -3,     0,     2,    -5,     0,     4,     2,     1,    -5,    -1,    -1,     1,    -6,     0,    -3,    -5,   -10,    -7,   -10,    -6,    -5,     0,    -6,    -3,    -1,     1,     0,     0,    -3,     0,     2,    -3,    -6,    -2,    -5,    -6,   -11,     2,     4,     1,    -1,     0,    -5,    -9,    -8,    -4,    -6,    -5,    -2,    -2,    -4,    -4,    -7,     2,     0,    -2,    -1,    -5,    -5,    -7,    -8,    -9,   -14,   -11,   -12,    -5,    -1,     5,     1,     1,    -3,    -8,    -4,    -4,    -3,    -3,    -4,    -5,    -3,    -4,    -2,     0,    -1,     1,    -4,    -4,   -10,    -4,    -7,    -3,    -8,    -9,   -12,    -8,    -6,     6,     4,     0,    -1,    -5,    -2,    -5,    -3,     0,     1,    -2,    -2,    -3,     0,    -1,     0,    -2,     2,     3,    -2,     2,    -2,    -3,     3,     3,     0,     1,    -7,     6,     4,     4,     3,     8,     1,     4,    -4,    -5,    -1,     2,    -3,    -2,     0,     2,     0,    -3,     4,     6,     3,     5,     5,    -1,    -3,     1,    -2,    -5,    -4,     2,     3,     6,     0,     6,     2,     6,     2,    -8,    -5,    -2,    -1,    -4,     0,     2,     2,    -8,    -4,     8,    10,     6,     3,     1,    -4,    -6,    -3,     0,    -3,    -2,    10,     4,    -3,     2,     1,     3,     1,    -4,    -5,    -3,    -1,     0,     0,     1,     1,    -2,    -4,     1,     0,     4,    -5,    -7,    -3,    -8,    -6,     1,    -1,     0,     2,     1,     0,     1,    -2,     1,    -3,     0,    -2,    -2,    -5,     7,    -1,     1,     0,     0,    -2,     0,     0,    -2,    -2,    -5,     5,     4,     1,    -2,    -8,    -8,     2,    -2,     3,    -5,   -13,    -6,    -4,    -7,    -5,    -6,     8,     9,     1,    -1,     0,    -1,    -1,     0,    -1,    -3,    -1,    -1,    -3,    -4,    -7,    -5,   -11,    -5,    -8,    -6,   -12,    -8,    -6,    -9,    -3,    -2,    -2,     0,    -1,    -2,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,    -1,    -3,     0,     0,    -9,    -6,     3,     2,     5,    -8,    -3,    -2,     0,    -2,     0,     0,     1,     0,     1,     1,    -1,     0,     0,     0,     1,     1,    -1,     0,    -1,     1,    -3,    -2,    -1,    -2,    -3,    -3,    -2,     0,     1,     1,    -1,     1,     0,     0,     0,     0,    -1,     1),
		    72 => (   -1,     0,     0,    -1,     0,     1,    -1,     1,     1,     0,     1,     1,    -3,    -3,     2,     1,     1,     1,    -1,     1,     0,     1,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,     0,    -5,    -3,    -5,    -7,    -5,    -7,    -3,    -5,    -2,    -3,    -5,   -10,    -7,    -2,    -2,    -2,     1,     0,     0,     1,    -1,     0,    -2,    -1,    -4,    -1,    -1,    -6,    -2,     6,     5,    -1,    -2,   -10,    -8,   -13,    -9,    -2,     0,    -2,   -11,    -3,    -4,    -2,     3,     1,    -1,     1,     0,     1,    -2,    -5,    -2,     1,     0,     0,     2,     2,     4,     0,    -6,   -12,    -9,   -11,   -10,    -9,    -9,    -8,    -9,    -7,    -4,    -2,     0,     0,     1,     0,     1,    -1,    -3,    -1,     1,    -3,     3,     3,     1,    -2,     4,     1,    -4,   -11,   -10,    -8,    -9,    -5,    -9,    -9,    -6,    -7,    -4,    -4,     0,    -1,    -4,    -2,    -1,     1,    -2,     0,     3,    -4,     6,     5,     6,     0,     3,    -3,     2,     0,    -4,    -1,   -11,   -11,    -8,    -5,    -3,    -6,    -7,    -2,    -4,    -1,    -1,    -2,    -1,     0,    -1,     1,     2,     6,     4,     1,     4,     4,     0,    -1,    -1,     3,    -1,    -5,    -6,    -6,    -6,    -3,    -2,    -6,    -5,    -4,    -7,    -2,    -2,    -2,     0,    -1,     0,    -2,    -1,    -1,    -4,    -2,     0,     1,    -5,    -1,    -1,    -1,    -4,    -4,    -5,    -1,    -6,    -7,    -6,    -8,    -9,   -10,    -7,    -4,    -4,    -2,    -4,     7,    -2,     0,    -7,    -2,     2,    -2,     1,    -3,     3,    -2,    -3,     4,     4,     1,    -2,    -2,    -4,    -5,   -10,   -11,    -9,    -9,   -10,    -4,    -6,    -3,    -1,    -4,    -2,     2,    -8,    -1,     0,    -3,     0,    -1,     2,     1,     2,     1,    10,     3,    -2,    -5,    -6,    -5,    -7,    -6,   -13,    -3,     8,    -7,    -2,    -3,     0,    -3,    -2,    -1,   -10,     3,     0,     0,     0,    -4,    -4,    -2,     1,    -2,     2,     6,     5,    -4,    -6,    -4,    -4,    -7,    -7,     1,     5,    -4,    -5,    -5,     0,    -1,    -7,    -3,    -4,    -3,    -3,    -2,    -3,     0,     2,     7,    -4,    -6,    -1,     2,     1,    -2,    -1,    -5,    -6,    -9,    -5,     1,    -1,    -5,   -10,    -1,    -1,    -1,    -8,    -1,    -1,     2,    -5,    -9,    -1,    -3,    -5,    -3,    -1,     0,    -3,    -1,     3,    -1,    -1,    -7,    -5,    -2,     1,    -8,    -2,    -3,    -4,     1,    -1,    -1,    -6,     0,    -1,    -2,    -7,   -10,    -2,    -4,    -7,    -4,    -3,     0,    -3,     2,     1,     1,    -3,    -4,     2,     6,     8,     1,    -2,    -1,     5,     5,     1,    -1,    -1,    -2,    -6,    -1,    -9,    -6,    -3,    -6,    -2,    -3,     0,     2,     1,     2,     3,     0,    -3,     0,     2,     6,     4,    -1,    -2,     0,    10,     5,     0,    -2,     5,    -4,    -1,    -1,    -1,    -5,    -3,    -1,     1,     0,     4,     7,     2,     3,     0,    -2,    -1,     0,     3,     1,    -3,    -5,     0,     2,     3,     6,     1,     0,     6,    -1,     3,    -4,     1,    -1,    -8,    -2,     2,     5,     1,     3,     3,     3,     6,     3,     1,     3,     0,     3,     2,     3,     2,     3,    -1,     6,    -1,     0,     9,     1,     5,    -2,     4,     1,    -2,     1,     3,     4,    -1,     1,     4,     4,     5,     3,     5,     7,     4,     5,    -2,     1,     0,    -3,    -7,     5,    -1,     1,     4,     3,     3,     2,     7,    -1,    -4,     1,     4,     4,    -3,     1,    -2,     3,     2,     1,     4,     2,     1,     4,     3,     5,     8,     4,    -5,     4,     0,    -4,     1,     7,    -1,     4,     3,     2,    -1,     5,     1,    -1,    -4,    -3,    -1,     4,     0,     0,    -2,    -3,    -3,     0,     4,     8,     5,     2,     4,     9,     0,    -2,     1,     5,     1,    -1,     1,    -2,     3,    -1,     0,    -1,    -1,     0,     1,     0,    -6,    -9,    -8,    -7,    -7,    -2,    -3,    -2,    -2,    -6,     4,    -1,     1,     0,    -1,     3,     2,     2,     8,     0,     0,    -1,     4,    -4,     1,    -3,    -4,    -4,   -12,   -18,    -2,    -3,    -6,    -7,    -8,   -10,   -10,    -5,    -5,     0,     1,     1,     0,    -1,     0,     3,     1,    -3,    -4,    -4,    -5,    -2,    -2,    -5,    -4,   -11,   -17,   -16,    -5,    -3,    -6,    -9,   -11,    -8,    -8,    -7,   -11,     0,     1,    -1,     1,    -1,    -2,    -2,    -3,    -5,     0,     0,    -7,    -8,   -14,   -12,   -16,   -13,   -15,   -15,   -10,   -11,   -10,   -11,   -10,   -13,   -10,    -6,   -11,     1,     0,     1,    -3,    -1,   -12,    -3,    -7,    -2,     1,    -5,     1,    -3,   -22,   -16,   -14,   -12,   -13,   -15,   -12,   -12,   -11,   -12,    -9,    -9,     2,     4,     4,     0,     0,     0,     0,     1,    -3,    -2,    -1,    -2,    -9,   -12,   -13,    -8,   -13,   -12,    -8,   -10,   -10,    -8,    -6,   -10,   -10,    -9,    -2,    -3,     0,     2,     3,     0,     0,    -1,    -1,     1,     0,    -4,    -6,    -6,    -9,   -11,    -8,    -3,    -3,    -4,    -6,    -2,    -5,    -4,    -2,    -7,    -4,    -2,    -5,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     1,    -2,    -3,    -1,    -2,    -4,    -2,     0,    -2,    -2,    -4,    -2,    -3,    -3,    -3,    -1,     1,     1,     0,     0),
		    73 => (    1,     0,    -1,     1,    -1,     1,     0,    -1,    -1,     0,     1,     1,    -2,    -1,    -2,     0,     0,     1,    -1,    -1,     1,     1,     0,     0,     1,    -1,     0,     0,    -1,     1,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -3,    -2,    -1,     0,     1,     0,     0,     1,     0,    -1,     0,     1,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,    -2,    -4,   -10,   -10,   -10,    -2,    -2,     0,    -1,    -1,     1,     0,    -3,    -1,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,    -1,     0,     1,     0,    -2,    -6,    -3,    -5,    -7,    -8,    -7,    -3,    -2,    -1,    -2,    -3,    -4,    -5,     0,     0,    -1,     0,    -1,     0,     1,     1,     0,    -1,    -2,    -7,    -5,   -13,     2,     4,    -1,    -1,     4,     1,     0,    -1,    -1,     0,    -1,     4,     8,    -5,    -6,    -5,    -1,     0,     0,     0,     1,    -1,     0,    -4,    -3,    -4,   -10,   -10,    -4,     4,     4,    -5,    -2,    -2,     0,    -3,    -3,    -4,     0,    -5,    -2,    -4,    -3,   -12,    -4,    -1,     0,     0,     3,     2,     0,    -4,     1,    -2,    -1,     3,     7,     2,    -1,     2,    -1,     2,     2,    -5,    -2,    -6,     1,     0,    -4,    -1,    -3,    -6,    -8,    -3,     1,     1,     1,     0,     1,   -11,    -9,    -4,     1,     1,     0,    -5,     1,     8,     1,    -3,    -4,    -1,     0,    -2,    -2,    -4,    -2,    -6,    -8,    -5,    -6,    -1,     0,    -1,    -1,    -2,     0,    -8,    -6,     1,     1,     1,    -2,    -2,     4,     3,    -1,    -2,     1,    -2,    -2,    -1,    -1,    -1,     0,    -3,   -15,    -5,   -10,     1,    -1,    -2,     1,    -2,    -5,    -4,    -2,     3,    -1,     1,     3,     6,     4,    -1,    -1,    -3,     2,     3,    -2,     1,     1,    -1,     2,     1,   -12,    -4,    -6,    -5,     0,    -3,    -1,    -1,    -3,    -5,    -2,    -5,     2,     1,     2,     6,     4,    -6,    -7,    -3,    -3,    -2,    -4,     2,     5,    -4,     1,    -1,   -11,   -10,    -9,    -4,    -1,    -4,     0,     3,     6,     4,     2,     0,     6,     1,    -6,    -7,   -22,    -8,    -3,    -4,    -3,    -1,    -3,     1,     3,     6,    -1,     3,    -9,    -6,    -4,     1,     0,    -2,    10,     2,     7,     4,     0,    -8,    -7,   -11,   -11,   -15,   -11,    -1,     0,    -2,    -2,    -4,    -3,    -1,     2,     5,     4,     3,    -6,     2,    -3,     0,    -1,    -4,    -5,    -6,    -7,    -6,    -5,   -17,   -15,   -11,    -6,    -4,     1,     6,     6,    -4,     1,    -1,    -2,     0,    -1,    -2,    -2,    -1,    -7,    -4,    -6,    -2,     0,     1,     3,    -3,    -5,   -13,   -13,   -15,    -2,     4,     2,    -2,     0,     3,     0,     1,    -1,     3,     0,    -5,    -6,    -3,    -3,     1,    -4,    -9,    -6,    -2,    -1,     0,     0,    -1,    -7,   -14,   -18,     6,     6,     1,     1,     3,     5,     5,     5,     1,    -1,    -1,     1,    -1,    -7,    -4,    -8,    -4,    -4,    -5,     5,    -1,    -1,     1,     3,    -2,    -3,    -5,    -2,    -2,     3,     5,     5,     5,     4,     3,     4,    -1,     0,    -3,    -1,    -3,    -8,    -6,    -5,     1,    -2,    -3,    -2,    -2,     1,     1,     2,     2,    -6,    -6,    -3,    -4,    -2,     2,     7,     3,     7,     6,     1,    -7,    -5,     0,    -2,     0,    -8,    -6,    -4,    -3,    -9,    -3,    -1,    -1,    -2,    -2,     1,     2,    -6,   -11,   -12,    -4,    -6,     0,     3,     5,     7,     1,     0,    -3,    -3,    -5,     2,    -1,     1,    -3,    -3,    -8,    -9,    -2,    -1,    -1,    -1,    -3,     0,    -1,    -9,    -8,   -10,    -9,   -12,    -9,   -11,    -4,    -8,    -3,    -6,    -3,     4,     2,     5,     1,    -4,     2,    -4,    -8,    -9,     0,    -5,    -1,     1,    -3,     2,     6,    -2,    -1,    -9,   -15,   -16,   -24,   -32,   -24,   -19,    -7,    -1,    -3,    -1,     4,     6,     4,     1,    -2,    -4,   -11,    -9,    -6,    -1,     1,    -2,    -1,     5,    10,     6,     0,    -1,    -6,    -1,    -5,    -5,    -8,    -5,    -4,     0,     2,     0,     0,     3,     0,     3,    -1,    -3,    -8,    -6,    -2,    -3,     1,    -1,     0,     1,     6,    11,    10,     7,     4,     4,     2,     5,     2,    -2,     1,     1,     1,     3,    -1,    -2,     0,    -3,    -2,    -5,    -4,    -6,    -3,     0,     0,     1,     1,     1,    -2,     7,     7,     6,     5,     1,    -2,     3,     0,     4,     7,     0,     4,    -7,     1,    -1,    -5,     3,     1,    -2,    -2,    -6,    -4,    -1,     1,    -1,    -1,     1,     5,     9,    -2,     5,     4,     0,     1,     4,     4,     3,     3,    -1,    -1,    -3,     2,   -13,    -4,     3,     3,     5,     5,    -8,    -2,    -3,     0,     1,    -1,     1,    -5,     0,    13,     9,     7,     3,     4,     1,    -2,     1,    -2,    -5,    -2,    -2,    -5,   -13,    -3,    -4,    -8,    -3,   -10,    -6,    -3,    -4,     1,     0,     1,     0,    -4,    -8,     0,     1,    -2,    -2,    -6,     0,     1,    -2,     1,     0,    -7,    -1,     3,     2,    -3,    -2,    -3,     1,    -1,    -1,     0,     1,     0,     1,    -1,    -1,     0,    -1,    -3,    -1,    -1,    -1,    -7,    -7,    -5,    -4,    -4,    -5,    -5,     0,    -1,    -2,    -5,    -5,    -1,    -4,     0,    -1,     0,     0,     0),
		    74 => (    0,     0,    -1,     0,     0,     1,     0,     1,     1,     1,     1,     1,    -1,    -4,    -1,     0,    -1,     0,    -1,     1,    -1,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,     1,    -1,     1,     1,    -5,    -5,    -2,    -4,    -8,    -4,    -9,    -5,     2,   -14,   -12,    -9,    -3,     0,    -6,    -1,     0,    -2,    -1,     1,     1,    -1,     0,    -1,    -2,    -5,    -8,    -5,    -3,    -7,    -4,    -4,   -12,   -16,   -12,    -3,     2,    -4,    -7,    -6,    -8,   -10,   -11,    -7,    -7,    -8,    -2,    -5,     1,    -1,    -1,     0,    -3,   -10,   -16,    -5,    -6,    -1,   -11,   -12,    -8,   -10,   -18,    -6,     2,    -1,    -5,    -7,   -10,    -3,    -2,    -5,    -3,    -9,   -10,    -4,     0,     0,     0,     0,    -2,   -14,    -1,     0,     1,     2,    -1,    -7,    -5,    -5,    -1,     4,     4,     2,     1,     3,     5,     0,    -3,     1,    10,     0,    -1,    -2,    -9,    -3,    -1,     1,    -3,    -6,     1,     3,     2,     8,     5,     3,     3,    -1,     3,     5,     8,     2,     0,     6,     2,     7,    -1,     5,     5,     8,     8,     4,    -9,     0,    -1,     0,    -3,    -2,     5,     4,     1,     9,     7,     8,     5,     3,     2,     8,    10,    13,     8,     2,    -4,     0,     3,     0,    -1,     8,    10,     3,     2,    -5,     0,    -5,    -4,     3,     6,     3,     5,     9,     4,    19,    12,    16,     9,    10,     9,     8,     5,     6,     2,     7,     3,    -3,    -2,     1,     4,    -4,    11,    -7,    -5,    -6,     6,     3,     3,     0,     7,     4,    -1,    16,     9,    10,     2,    -2,    -1,     3,    -3,    -3,    -3,    -1,     1,     1,    -7,    -2,     0,     3,     5,    -8,     1,    -2,     5,    -4,     1,    -4,    -5,    -3,    -2,     0,     3,    -7,    -3,     1,    -2,     1,    -5,     2,    -1,    -2,    -2,    -2,    -8,     0,    -2,    -5,    -5,    -4,     1,    -3,     3,    -3,    -3,    -6,   -10,    -4,    -5,     1,    -3,    -8,     0,    -6,    -5,    -3,    -3,     0,    -7,     0,    -8,    -4,    -2,    -5,   -11,    -3,    -1,    -6,     1,    -5,     3,    -4,    -5,    -4,     4,    -8,     1,    -3,    -7,    -2,    -1,    -2,    -4,    -1,     1,     4,    -6,    -5,   -13,    -5,    -4,    -8,   -13,    -3,    -5,   -10,    -1,     1,     1,    -4,    -7,    -2,    -1,    -5,    -1,     1,    -4,     2,     8,     4,    -7,     0,     1,     3,    -2,    -3,     0,     4,    -2,    -5,     1,     6,    -5,    -9,     0,    -2,    -7,    -7,    -7,    -1,     1,     7,     4,    -3,     2,     7,     9,    -1,     2,     1,     0,     4,     4,    -1,     0,    -4,    -5,    -2,     1,     4,    -2,    -1,    -1,     4,   -13,    -9,     0,     0,     0,    12,     7,     4,     7,     5,     3,    -2,    -3,    -1,     2,     1,    -2,    -1,    -5,    -7,    -2,    -1,     0,     5,    -7,    -1,    -1,     1,     5,     1,     6,     0,     4,     6,     7,     3,     1,     1,     6,     4,     1,    -1,     3,     6,    -2,    -3,     0,     1,     6,     3,    -2,    -1,    -4,    -7,     1,     0,    -8,     2,    -3,    -3,    -3,    -2,     0,     0,     4,     3,     0,     0,     1,    -1,     2,     3,     1,     3,     6,     4,     4,    -1,     3,     1,    -4,    -3,     0,    -1,    -5,    -6,     0,     0,    -4,     6,     1,    -1,    -7,    -3,     1,    -5,    -1,    -5,     5,    -1,    -2,     2,     0,     4,     2,     8,     2,   -10,    -2,    -3,    -5,    -1,    -2,     0,     1,     5,     3,     1,    -5,    -2,    -7,    -5,     2,    -3,     1,    -3,    -4,    -8,    -2,     6,    10,     6,     4,     7,     5,    -3,    -4,    -6,     0,    -5,    -7,    14,    -4,    -2,    -4,    -7,    -3,    -6,    -7,    -8,    -1,     1,     2,     3,     1,    -8,     0,     3,     4,     3,     5,     1,     2,    -1,    -2,    -5,     1,    -2,    -4,     3,    -4,    -7,    -7,    -8,    -4,     3,     1,     1,     0,    -1,     0,     3,     4,    -1,     5,     5,     7,     5,     2,    -2,    -7,    -8,    -4,    -1,    -2,    -1,    -5,     4,     3,    -3,    -5,    -4,     1,     2,     0,     2,    -5,    -3,    -2,     3,     4,     3,    -1,     6,    14,    11,    11,     3,    -3,   -12,    -8,     0,    -2,    -2,    -2,    -7,   -14,    -8,     0,     3,     6,    -2,     7,     1,    -1,     0,    -5,    -3,     6,     5,     0,    11,    12,    13,     8,     7,     1,     0,    -2,    -2,     1,     1,     0,   -10,   -12,   -23,     4,     6,    10,     6,    11,     8,     3,     0,    -2,    -3,     2,    -1,     5,    11,    11,     5,    -5,     5,     0,     7,    -2,     0,     0,     1,     1,    -4,   -12,    -2,    10,    10,     3,     8,     1,     9,    -3,     0,     0,    -8,    -4,    -4,     6,    10,     0,    -3,    -2,    -1,    -6,     6,    -6,    -1,     0,     0,    -4,     0,    10,    14,     5,    -4,    -3,     1,     5,     5,    -5,     3,    -7,     2,     1,    -1,    -2,    -1,    -2,    -2,    -2,     1,    -3,    -7,    -5,     1,     0,    -1,     0,    -9,    16,    13,     8,    -3,    -6,    -9,   -15,    -3,    -5,    -5,    -3,   -11,   -12,    -8,    -2,    -1,    -9,   -18,   -16,    -4,     1,    -1,     1,     1,     0,    -1,     1,    -1,    -2,     0,    -5,    -6,    -4,    -5,    -6,    -8,    -6,    -2,    -5,    -2,   -10,   -15,   -12,    -7,    -7,    -3,    -5,     1,     1,     0,     0,     0),
		    75 => (   -1,     1,    -1,     0,     0,     0,    -1,     1,    -1,    -1,     0,     0,     1,     0,     0,    -1,     1,     0,     1,     0,     1,     1,     0,     0,     1,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,     1,     1,    -1,    -1,    -2,    -4,    -3,    -2,    -2,    -4,    -3,     0,    -1,    -2,     0,     1,    -1,     1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -3,    -2,    -6,    -6,    -7,    -7,    -4,    -5,   -12,    -2,     1,     1,    -1,     4,     6,     0,     0,     2,    -3,    -1,     1,     0,     0,     0,    -1,     2,     3,    -5,    -6,    -6,    -4,    -2,    -2,    -3,     1,     2,     4,     4,     3,    -1,    -4,    -3,     1,     4,     1,     3,     2,     1,     2,     1,     1,    -1,     0,     3,     0,    -1,     3,     5,     1,     5,     0,    -6,    -4,     0,     2,     5,     6,     1,     0,    -4,    -1,     0,     3,     4,     3,     4,    -2,    -4,    -1,     0,     1,     1,    -3,     0,     5,     3,     3,     1,    -1,    -5,    -6,    -1,     0,    -1,     0,     0,    -1,     6,     5,     0,     4,     4,     4,     3,    -3,    -3,     0,    -1,    -5,    -4,     2,     3,     7,     2,     1,    -1,     0,    -3,    -4,    -2,    -1,     0,    -1,    -3,     1,     6,     7,     5,     4,     2,     4,     4,     3,     1,    -1,     1,     0,    -4,     1,     8,     1,     2,    -3,    -1,    -2,    -1,    -2,    -3,    -1,    -3,     0,    -1,    -2,     0,     3,    -1,     4,     3,     7,     4,     3,     4,    -1,    -4,    -4,    -7,     1,     0,     0,     1,    -2,     1,     0,     3,     2,     2,     0,    -4,    -4,    -6,     1,     2,    -2,     0,     6,     7,     4,     5,     3,     2,     0,    -2,    -9,    -6,     1,     1,     0,     0,    -3,    -2,     3,     4,     6,     5,    -2,    -3,    -5,    -5,    -2,     0,     2,     6,     7,     7,     6,     1,     5,     1,     1,     0,    -1,    -9,     0,     0,    -1,     2,    -3,     1,     0,     6,     8,     1,     4,     0,    -6,    -2,     0,     3,     7,    10,    10,     7,     7,     3,     0,    -3,     1,    -1,    -1,    -6,     2,     0,     1,     2,     3,    -1,    -2,     6,     4,     0,     4,    -3,    -5,    -8,     6,     5,     9,     4,     4,     5,     6,     5,     1,    -4,     0,     1,     0,    -7,     2,     3,     4,     4,     6,     4,    -4,     0,     2,     1,     1,    -2,    -5,    -1,     3,     6,     4,     0,    -1,     4,     2,     3,     6,    -4,    -1,     0,    -1,    -8,     0,     2,     3,     5,     4,     5,     7,     3,     3,    -2,     0,    -5,    -3,    -2,     0,     5,     5,     5,     0,    -3,    -3,     0,     5,    -4,     1,     0,    -2,   -10,    -1,     1,     4,     5,     4,     3,     7,     1,     1,     0,     0,    -4,    -2,     2,     7,     6,     5,     4,     3,    -3,    -5,    -5,    -3,     0,     1,    -1,    -3,    -1,     2,     4,     0,     2,     4,     6,     7,    -1,    -1,     0,     4,     1,     0,     3,     4,     6,     3,     3,     2,     0,     1,    -5,    -3,    -7,     0,    -2,    -5,    -1,     2,     9,     2,     1,     4,     4,     4,    -4,     1,     1,     1,     3,    -3,     1,     0,     1,     5,     9,     4,     0,    -2,    -5,    -4,    -8,    -1,     0,    -4,     2,     3,     8,     6,     5,     6,     6,    -2,    -2,    -4,     0,     4,    -3,     1,    -1,    -1,     0,     4,     2,     4,     1,    -1,    -5,    -9,    -9,     0,     0,    -5,     1,     1,     7,     6,     4,     7,     5,    -1,    -5,    -8,     2,     3,     0,    -1,    -2,    -3,    -4,    -1,     0,    -1,     2,     2,    -4,   -10,    -6,     1,    -1,     4,     0,     2,     4,     4,     8,     5,     0,    -3,    -3,    -4,     3,     0,     1,    -3,     1,    -1,     1,     1,    -1,     0,     4,     1,    -4,   -11,    -5,     1,    -1,     3,     2,     2,     2,     4,     5,     7,     0,    -3,    -4,     1,     0,    -3,    -2,    -1,     1,     4,     4,    -2,     2,     2,     4,    -5,    -1,    -8,     0,     0,     0,     1,     1,     1,     4,     4,     6,     6,     5,     0,     3,     2,     1,     0,    -1,     0,     0,     2,     4,     5,     1,     2,     1,    -5,     0,    -5,    -1,    -1,     0,    -5,    -1,     2,     1,     4,     3,     6,     4,     2,     6,     3,     1,     1,     1,    -2,    -3,    -2,     1,     2,    -3,    -2,    -3,    -7,     1,     4,    -1,     0,     0,     1,     0,    -3,    -1,     3,     5,     3,     2,     0,     3,     3,     3,     2,    -2,    -7,    -5,    -3,    -3,    -1,    -5,    -3,    -5,    -2,     2,     3,     1,    -1,    -1,    -1,     0,    -4,    -2,     3,     2,     1,     3,     4,     3,     1,    -2,     1,     0,    -4,    -4,    -2,    -4,    -4,    -3,    -3,    -2,     1,    -8,    -3,     0,     1,     0,     1,     4,    -7,    -6,    -1,     2,    -3,    -4,     4,     2,     2,     1,     0,     2,     3,     5,     4,    -1,     3,     2,     6,     2,     0,     0,    -1,     0,    -1,    -1,     0,    -4,    -6,    -8,    -9,    -1,     0,    -2,    -2,     4,    -1,     1,     4,     2,     3,     1,    -2,    -1,    -4,    -3,     1,    -5,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -1,     0,     1,     0,    -2,    -1,    -2,    -1,     0,     1,    -1,    -3,    -2,    -6,    -5,    -2,    -1,     1,     1,    -1),
		    76 => (    1,     0,     1,     0,     0,    -1,    -1,     0,     1,     1,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,     1,    -1,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     1,     2,     2,     4,     2,     1,     2,     2,     1,    -1,    -2,    -3,     1,     0,     0,     7,     3,     1,     2,     1,     0,     0,     0,     0,     0,     1,     1,     6,     2,     0,     4,     5,     1,    -2,     0,     0,     1,    -3,    -2,    -2,     2,     0,     2,     2,     8,    10,     8,     8,     4,    -1,     0,     1,     0,    -3,    -3,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -8,    -7,    -7,    -4,    -5,    -6,     2,     8,     8,     5,     2,     7,     7,     1,    -6,    -1,     1,     1,    -2,     0,     3,     1,    -2,    -3,    -4,    -1,    -2,    -4,    -7,    -9,   -10,    -8,    -3,    -4,    -3,     1,     1,     6,     1,     7,     2,    -2,     4,     5,    -1,    -1,    -3,    -4,     3,     1,    -1,    -2,    -2,    -1,    -4,    -6,    -6,    -6,    -5,    -2,    -3,    -1,     0,     0,    -2,     2,     4,     6,     7,     6,     8,     5,    -1,    -1,     0,    -1,     1,     2,    -2,    -1,    -4,    -1,    -4,    -4,    -3,    -4,    -8,    -8,    -7,    -2,    -2,     2,     0,    -2,     1,     5,     7,     4,     3,     7,     1,    -1,     0,     0,     3,     2,    -4,    -1,     0,     3,    -6,    -6,    -5,    -9,    -6,    -9,    -3,     0,     2,    -3,    -3,     1,    -3,    -3,     2,     4,     3,     8,     0,     0,     0,    -2,     4,     0,    -7,    -3,    -2,    -1,    -8,    -8,    -9,    -9,    -8,    -5,     1,     1,     2,     0,     0,    -2,    -2,    -1,    -7,    -4,     6,    -4,     1,    -1,     0,    -3,     6,    -1,    -6,    -1,     2,    -1,    -7,    -8,    -9,    -9,    -5,     2,     3,     1,    -1,     1,    -1,    -3,    -2,    -5,    -6,    -4,    -3,    -2,    -1,    -1,     0,    -2,     4,    -1,    -4,    -1,    -1,    -6,   -13,   -10,    -7,    -1,     0,     3,    -2,    -3,    -7,    -8,    -2,    -2,    -5,    -5,    -4,    -4,    -3,    -4,     0,    -1,     1,    -3,     2,     1,    -7,    -6,    -5,   -13,    -8,    -7,    -3,     0,     3,     0,    -3,   -10,   -13,    -8,    -8,    -5,    -3,    -4,    -7,    -1,    -1,    -2,    -1,    -1,    -1,    -5,     1,    -2,    -5,    -6,    -8,    -8,    -8,     1,    -3,     2,    -1,    -2,    -3,    -7,   -11,    -8,    -6,    -4,    -2,    -3,     0,    -2,    -4,    -2,     1,     1,    -1,    -3,    -1,    -1,    -4,    -5,     0,    -2,    -3,    -2,     2,     3,    -2,     1,     0,     0,    -2,    -2,    -1,    -8,    -4,    -1,    -1,     0,    -4,    -1,     0,     0,     0,    -3,    -3,    -3,    -3,     1,     4,    -3,     1,    -2,     3,     1,     1,    -4,     2,     0,    -1,     0,     1,    -5,    -9,    -8,    -1,     0,    -2,    -2,     0,     0,    -3,    -1,    -3,    -4,     3,     2,    -2,     1,    -2,     2,     4,     0,    -1,    -2,    -1,     2,     1,    -3,    -6,    -6,    -8,    -3,    -2,    -1,    -1,    -4,     1,     1,    -2,    -3,     1,    -4,    -2,    -1,     1,     1,     0,     1,     3,     2,     0,     1,    -1,    -3,     1,     1,    -5,    -7,    -4,    -2,    -3,     1,    -2,    -2,    -1,    -1,    -3,    -5,    -1,    -5,    -4,     1,     2,    -1,     6,    -3,    -2,    -5,    -4,    -3,    -4,    -5,     5,     3,     1,    -4,    -1,    -2,    -3,    -2,    -3,    -6,     1,    -1,    -1,    -1,     4,    -2,    -5,    -2,     0,     1,     0,    -2,    -5,    -4,     0,     2,     0,     0,     6,     8,     5,     0,    -2,    -3,    -2,     0,    -6,    -1,     0,    -1,     1,    -3,     3,    -3,    -3,     1,    -4,     2,    -1,    -5,    -2,    -6,     0,     4,     1,     3,     7,     5,     4,     1,    -5,    -3,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -3,     3,     0,     5,     2,    -2,    -1,     0,    -2,    -2,     0,     7,     1,    -2,    -3,     0,     1,     0,    -3,    -4,    -4,     0,    -1,    -1,     0,     1,    -1,    -4,    -3,     1,     0,     0,     0,     4,    -4,     2,     5,     5,     3,     2,     0,    -1,    -3,    -3,    -4,    -6,    -5,    -4,    -1,     0,    -1,     0,    -1,     0,     0,    -2,     1,    -1,    -2,    -9,    -3,     4,    -2,     0,     4,     7,     3,    -5,    -5,    -2,    -6,    -4,    -5,    -5,    -1,    -1,    -4,    -2,    -4,     1,     1,    -1,    -1,     0,    -3,    -4,    -2,    -5,     3,     2,     1,     3,     4,     4,     1,    -1,    -3,    -1,    -7,    -6,    -4,     0,    -1,     0,     1,    -3,    -3,    -1,     1,     1,     1,    -1,     0,    -2,    -2,    -1,    -1,    -3,    -3,    -1,    -3,    -1,    -3,    -1,    -1,     2,     0,     0,    -3,    -1,    -2,    -1,     1,     0,    -1,     0,     0,    -1,     1,    -1,    -1,     0,    -4,    -5,    -6,    -3,    -2,    -1,     0,     0,    -1,    -1,     1,    -2,     0,    -1,    -1,    -4,    -1,    -1,    -2,     0,    -1,     0,    -1,     1,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -1,     0,    -3,    -2,    -1,     0,     0,     0,    -1,     0,     0,     1,    -3,    -1,    -2,     0,     0,     1,    -1,     1,    -1,     1,     1,     1,     1,     1,    -1,     1,     1,     1,     1,     0,     0,     0,    -1,     0,    -1,    -1,     1,     0,    -1,    -2,     1,     0,     0,    -1,     0,    -1),
		    77 => (    0,     0,    -1,     1,     1,     0,    -1,     1,     0,     0,    -1,     1,    -1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -1,     1,     1,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -2,     0,    -1,    -1,    -1,    -4,    -5,    -3,     1,     1,     1,     0,     0,     0,     1,     0,     0,     1,     1,     1,     0,    -1,     0,     1,     0,    -1,     0,     0,    -3,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,    -3,    -3,    -3,    -4,    -2,    -3,     1,    -4,    -4,    -9,    -3,    -4,    -3,    -2,    -5,    -1,    -2,    -1,    -1,     1,     0,     0,     1,    -1,    -3,    -2,    -3,    -8,    -7,    -6,    -8,   -12,   -14,   -11,    -7,   -14,   -10,   -12,   -11,    -6,    -7,    -3,    -9,    -5,    -3,    -3,    -1,    -1,    -1,     1,    -1,    -5,    -1,     7,     5,     4,     9,     8,     0,     3,     1,     3,    -2,     0,    -1,    -5,     0,    -3,    -5,   -10,   -11,    -8,   -10,    -8,    -3,    -1,     1,     0,    -1,    -3,    -2,     4,     5,     7,     7,     0,     1,     4,     6,     6,     8,     2,     7,     5,     3,     4,     5,     1,     3,    -1,    -1,    -3,     0,    -2,     0,     1,    -2,    -1,    -3,    -2,    -3,     5,    -1,     1,    -1,     5,     8,     7,     3,     4,     3,     7,     1,     2,     4,     0,     0,    -1,     1,    -1,    -2,    -1,    -3,     2,     0,    -2,    -2,    -5,    -5,    -4,    -7,    -6,    -7,     0,     1,    -2,     1,     2,    -1,     3,    -2,     0,    -4,    -3,    -6,    -5,    -5,    -2,    -4,    -4,     0,    -1,    -2,     1,     0,    -4,    -7,    -6,   -12,    -4,    -7,    -5,    -4,    -6,    -3,    -5,     1,    -6,     0,    -1,    -4,    -3,    -3,    -5,    -4,    -1,    -4,     2,    -1,    -2,    -5,    -4,     0,    -5,     0,    -3,    -5,    -3,    -6,    -4,   -10,   -12,   -12,    -3,    -2,     1,    -2,    -3,    -1,    -9,    -2,    -7,    -5,    -2,    -5,     2,    -1,    -1,    -4,    -1,    -4,    -4,    -4,    -8,   -10,    -8,   -13,    -9,   -14,    -9,    -6,    -2,     0,    -2,    -3,    -3,    -3,    -3,     4,     4,    -3,    -8,    -4,     3,     0,     0,    -2,     1,     0,    -3,    -5,   -10,    -8,   -12,    -8,   -10,    -8,    -5,    -4,    -2,     0,    -6,    -7,    -3,    -4,     1,     1,    -2,     0,     0,    -2,     3,     1,     0,     2,     0,    -2,    -4,    -3,     1,    -4,    -1,    -3,    -2,    -2,     0,    -1,     1,     3,    -3,     0,    -1,     4,     4,    -2,    -5,    -4,     0,    -5,    -4,    -1,     0,     0,    -2,     3,     0,     2,     4,     0,     1,     1,     3,     4,     3,     3,     2,     3,     0,     2,     8,     0,     1,     2,    -9,    -5,    -3,    -3,     1,     0,     0,    -2,     1,     4,     3,     3,     5,     5,    -1,     2,     0,    -2,     1,     0,     2,     6,     3,    -1,    -2,    -4,     1,    -3,   -10,   -10,    -6,    -1,    -2,     1,    -1,    -2,    -3,     1,     0,    -1,    -6,     0,     0,    -1,    -4,     0,     1,     1,     5,     2,     0,     0,    -2,     1,    -2,    -6,    -8,    -9,    -6,    -4,    -3,    -1,    -1,    -3,    -3,    -4,    -2,     4,    -5,    -2,    -1,    -2,     3,     0,    -2,     2,    -2,    -4,    -4,     0,     0,     3,    -1,     1,    -2,     2,     3,     5,    -6,     0,     0,    -1,    -3,     0,    -3,    -3,    -2,     0,    -6,    -3,     3,     2,    -2,    -1,    -1,   -10,    -7,    -1,     1,    -3,    -4,    -6,    -5,    -2,     3,     7,    -6,    -1,     1,     1,    -2,     3,    -4,    -1,    -7,    -8,    -2,    -4,     0,    -4,    -3,    -1,    -5,   -13,    -6,    -1,    -2,   -11,   -13,    -7,    -8,    -3,     4,    -3,    -2,     1,     2,     1,    -1,    -4,    -1,    -3,    -5,    -4,    -2,     0,     3,    -3,    -3,    -3,    -6,    -8,    -4,   -11,   -10,    -4,    -5,    -6,    -3,    -7,    -8,    -2,    -1,     0,     0,    -1,     0,    -3,     3,     0,     1,    -2,     1,     1,     0,     4,     2,    -3,    -2,    -4,    -2,    -6,    -4,    -9,    -6,    -3,    -2,    -4,    -4,    -1,     0,     1,     0,    -2,    -2,     5,     0,    -2,     2,     3,     0,     0,     1,     0,     2,    -6,     0,     3,     0,    -3,    -8,   -10,    -6,    -2,     0,    -6,    -2,    -3,     1,     1,    -1,    -2,    -8,    -1,    -6,     1,    -1,     0,    -3,    -2,    -1,     0,     4,    -3,    -2,    -7,    -8,    -5,    -4,    -9,    -4,    -4,     0,    -1,     0,    -3,    -1,     0,     0,    -2,    -5,    -2,    -4,     0,     4,     2,     1,    -5,     1,     2,     3,    -1,     4,    -7,    -8,    -2,    -2,    -8,    -8,    -6,     1,    -1,    -4,    -2,     1,     1,    -1,     1,     2,     2,     1,    -6,     2,     3,    -7,    -1,     3,     4,    -3,    -2,    -5,    -9,    -5,    -3,    -3,    -5,    -4,    -2,     0,     0,    -1,     0,     0,     0,     1,     0,    -4,    -1,    -4,    -1,     5,     5,     4,     0,     0,     4,     4,     5,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,    -1,     1,    -1,     0,     0,    -1,     1,     2,     0,     0,    -1,     2,    -1,    -2,     0,     1,     2,     1,     0,     0,     0,     2,     1,    -1,     0,     1,     2,     1,     1,     0,     0),
		    78 => (   -1,    -1,     0,     1,     1,     1,     0,     0,     0,     0,    -1,     1,     0,    -1,     1,     0,     0,     1,     0,     0,    -1,     0,     1,    -1,    -1,     1,     1,     1,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     0,    -1,     1,     0,    -1,    -3,    -6,    -4,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,     0,     1,    -1,     0,     1,     1,     0,     0,     0,    -2,    -3,    -7,    -5,    -2,    -1,    -1,     0,     0,    -2,    -2,    -1,    -2,    -3,    -5,    -2,    -2,    -2,     0,     1,     0,     0,    -2,     0,     0,    -4,    -3,    -6,     4,     2,    -1,    -2,     0,    -2,    -4,    -2,    -1,    -3,    -1,    -2,    -2,    -2,     0,     1,     0,    -2,    -3,     1,     0,     1,     0,     0,    -4,    -6,    -1,     0,    -2,    -6,    -6,    -7,    -2,    -2,    -1,    -5,    -2,     4,     5,    -2,    -2,    -3,    -4,    -3,    -1,    -2,     1,    -2,     1,    -1,    -1,    -1,    -4,    -5,     1,     1,    -3,    -7,    -5,    -4,    -4,    -1,    -2,     0,     0,     1,     3,     2,     0,     0,    -2,    -1,    -1,    -1,    -1,    -4,     0,     1,    -3,    -6,    -1,    -5,     0,     1,     0,    -1,    -4,    -3,     1,     1,     0,     2,    -1,    -1,     0,     0,     1,     0,     1,     0,     0,     0,    -1,     1,     0,    -5,    -2,     0,    -3,    -2,     2,     0,     1,     1,     3,     0,     1,    -3,    -1,     4,     1,    -1,     4,    -3,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,    -2,    -3,    -2,     0,    -3,    -2,     3,     0,    -1,     0,     1,     0,    -2,    -2,     0,     4,     2,    -5,     1,    -1,    -5,    -2,    -1,     0,    -1,     2,     0,     0,     0,    -2,    -5,     0,    -1,    -6,     1,    -1,     1,    -1,     0,    -4,    -3,    -2,    -1,     4,     1,    -5,     2,     0,    -1,     0,     0,    -2,    -4,    -1,    -3,    -6,     0,    -1,    -5,     1,    -1,    -6,    -5,     1,    -1,    -4,     1,     0,    -1,    -4,    -5,     2,    -3,     1,     0,     0,    -1,    -3,    -3,    -5,    -4,    -1,     4,    -4,     0,     1,    -2,     0,    -3,    -5,    -5,     2,    -2,    -5,    -2,    -3,    -5,    -6,    -2,     3,     0,     0,     3,     1,    -2,    -6,    -3,     2,     0,     0,     5,    -5,    -1,     1,    -3,    -3,    -4,    -3,    -4,     0,     0,    -3,    -3,    -3,    -2,    -5,    -5,     3,     3,     1,     2,     1,     0,     1,     2,    -3,    -2,    -3,    -2,    -7,    -1,     0,    -4,    -3,    -5,    -4,    -4,    -1,    -2,     0,    -6,    -4,    -7,    -7,    -3,     0,    -2,     1,     4,     1,     0,     2,    -2,    -3,    -3,    -4,    -4,     0,     0,     0,     0,    -3,    -1,    -3,    -6,    -2,    -1,     0,     0,    -2,    -1,    -9,    -2,    -3,    -6,    -4,    -2,     0,     0,    -1,    -4,    -4,    -4,    -1,   -12,    -1,     0,     1,     0,    -2,     0,     0,    -3,    -3,    -3,     1,     0,    -4,    -1,    -6,     0,     0,    -2,     0,    -2,    -2,    -2,    -1,    -2,    -3,    -2,    -1,   -10,    -4,     0,    -1,    -1,    -2,     1,    -2,    -2,     0,    -1,    -3,    -2,    -2,    -4,    -2,     2,     0,    -2,     1,    -2,    -2,    -3,    -1,    -3,    -2,    -1,     0,    -6,    -4,     1,     0,    -1,    -1,     0,    -2,    -3,    -1,    -2,    -6,    -5,    -4,    -6,     1,     3,     2,    -2,    -4,    -1,    -1,     0,    -2,    -3,    -1,     0,    -1,     0,    -4,     0,     1,     0,    -3,     0,    -2,    -2,     0,    -3,    -4,    -1,    -5,     0,     2,     1,    -1,     1,    -4,     0,    -1,    -2,    -4,    -1,    -2,     1,    -1,     0,    -2,     0,    -1,    -4,    -4,     1,    -2,    -1,    -4,    -6,     0,    -1,    -2,     2,     2,     0,     3,     4,    -2,    -1,    -2,    -3,    -2,    -2,    -1,    -1,     0,    -6,    -5,     0,     1,    -1,    -1,     0,    -4,    -3,    -2,    -3,     2,    -1,    -2,    -1,    -2,    -4,     0,    -1,     2,     1,    -1,    -5,    -3,    -3,    -1,     0,    -1,    -5,     1,    -4,    -2,    -2,     0,    -2,    -5,    -3,    -6,     0,     4,     0,    -5,     1,    -2,    -4,    -5,     0,     5,     1,     1,    -3,    -1,    -2,    -2,    -2,     0,    -5,     0,    -2,    -2,    -1,    -2,    -1,    -4,    -2,    -3,    -2,     3,     2,     1,     1,    -2,    -4,    -4,     3,     3,     0,    -1,    -2,    -5,    -4,    -2,    -2,    -1,    -4,     1,     0,     1,    -2,     0,    -2,    -3,    -3,    -2,    -3,     0,     2,     2,     7,     2,     1,     0,     6,     0,    -2,    -6,    -3,    -2,    -3,    -1,    -2,     0,    -6,     1,     0,    -1,    -1,    -2,     0,    -2,    -4,    -3,    -3,    -2,    -3,    -3,     1,     0,     1,     1,     3,    -6,    -6,    -5,    -4,    -2,    -1,    -1,    -4,    -1,    -1,     0,     0,     1,    -3,    -3,    -1,     0,    -2,    -4,    -4,    -4,    -3,    -9,    -1,     1,     1,     4,    -6,    -8,    -6,    -4,    -1,    -2,     0,     1,     0,    -2,    -2,     1,     0,     1,     1,    -1,     1,    -3,    -3,    -2,     0,    -3,    -5,    -6,    -5,    -7,    -9,    -4,    -2,     0,    -1,    -2,    -7,    -4,    -4,    -1,     0,     1,     0,     0,     1,    -1,     0,     0,    -1,     0,    -2,     0,    -2,    -1,    -2,     0,     1,    -3,     0,    -1,    -3,    -4,     0,     1,    -1,    -1,    -1,    -1,     0,    -1,     1,     1),
		    79 => (    0,     0,     1,     0,     0,     1,    -1,     0,     0,    -1,    -1,     0,     1,     1,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,    -1,     1,     1,     0,     0,     1,     1,     1,     1,     1,     1,     0,    -2,    -2,    -2,     1,     0,     1,     0,    -1,     0,    -1,     0,     1,     1,    -1,     0,     1,    -1,     0,    -1,     1,    -1,     1,     0,    -1,     0,     0,    -2,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     0,     0,     0,     1,     0,     0,    -1,     0,     1,    -1,    -1,    -1,    -2,    -1,    -3,    -5,    -1,    -3,    -5,    -4,    -4,    -1,     2,     4,    -2,    -1,    -3,    -1,     0,     0,     1,     0,     0,     1,     1,     0,     0,    -1,    -5,    -1,    -1,    -4,    -4,     4,     3,     3,     0,    -4,    -4,    -6,    -8,    -7,    -9,    -4,    -3,     1,     0,    -4,    -3,    -1,    -1,     1,     0,    -1,     0,     0,    -1,    -2,    -8,   -10,    -6,     7,     0,     1,    -2,     3,     9,    -3,    -1,    -1,     3,    -4,    -5,    -2,    -3,    -4,    -5,    -1,     0,    -4,    -1,     0,    -1,    -5,    -1,    -8,    -3,    -4,    -3,    -4,     3,     3,     5,     3,     1,     2,    -3,    -6,    -7,    -1,    -3,    -2,    -1,    -2,    -3,    -2,     1,    -1,    -2,     1,    -1,    -8,    -8,   -15,     6,    -9,     2,     6,     3,     2,     2,    -3,    -3,    -8,   -14,    -7,    -4,    -3,    -3,    -3,    -2,    -2,    -3,    -3,    -2,    -6,    -2,    -2,    -2,    -5,   -10,   -11,     7,    -2,     5,     6,     5,    -3,    -9,    -2,    -6,    -2,    -5,     3,    -2,    -4,    -2,    -4,    -5,    -3,    -8,     0,     0,    -4,    -2,    -1,    -6,    -6,   -14,    -2,     6,     0,     3,     1,    -7,    -7,    -5,     0,    -1,     3,    -5,     2,    -1,    -5,     1,    -3,    -2,    -6,    -3,    -2,     0,    -1,     0,     1,    -3,    -3,    -6,     4,     7,     4,    -3,     1,    -5,     3,     9,     6,     0,     4,     6,     4,    -4,   -10,    -4,    -6,    -3,    -4,     0,    -4,    -1,    -3,     0,    -1,    -3,    -3,    -2,     0,     4,     1,     1,     0,     5,     6,     9,     3,     5,     7,     2,     0,    -4,    -5,    -6,    -5,    -1,    -5,     0,    -4,     1,    -1,    -2,     0,    -1,    -3,    -6,    -3,    -2,    -2,    -2,     1,     0,     5,     0,     1,     2,     2,     0,     1,    -2,    -3,     0,    -9,    -9,    -4,    -5,    -1,     1,    -2,    -2,    -5,    -3,    -3,    -6,    -1,    -2,     1,    -5,    -2,    -1,     3,     0,     6,     5,     0,   -10,    -4,    -5,    -7,    -2,    -4,    -5,    -3,    -5,     0,     0,    -1,    -3,    -4,    -3,    -3,    -6,    -2,    -8,    -1,    -5,    -3,    -1,     3,    -3,    -2,     2,     1,    -4,    -7,    -5,    -1,     4,    -1,     0,    -4,    -2,    -1,     1,     1,    -1,    -3,    -1,    -2,    -2,   -12,   -11,     0,     3,     5,     4,    -1,    -1,    -5,     2,     2,    -9,    -7,    -9,     1,     3,    -2,     1,    -2,    -2,    -3,    -1,    -1,    -2,    -2,     0,    -3,    -3,    -6,   -15,   -13,    -7,     0,    -2,    -8,    -5,    -5,    -1,    -5,    -4,   -11,    -7,    -2,     2,     0,     1,    -3,     1,    -1,     0,    -1,    -3,     0,     0,     3,     2,    -3,    -5,   -10,   -12,   -19,   -10,    -6,    -2,    -4,    -3,    -3,    -5,   -10,    -6,    -2,    -5,    -5,     3,    -1,    -2,    -1,     4,     1,    -3,    -2,    -2,    -4,    -3,    -4,    -5,    -6,    -8,   -16,    -7,    -3,    -2,    -6,    -2,    -1,    -5,    -9,   -12,    -5,    -6,    -8,    -4,    -1,    -1,    -2,     1,    -2,    -1,     0,    -1,    -7,    -8,     5,    -5,    -6,    -7,   -10,    -3,    -3,    -2,    -3,    -4,    -7,    -3,     0,    -9,     2,     0,    -1,    -2,    -2,    -3,     1,     0,    -2,    -2,    -1,    -2,     2,    -5,     2,     2,    -3,     0,    -3,    -2,    -2,    -4,    -6,    -4,    -5,     0,    -3,    -8,     0,     3,    -1,     5,     1,    -1,     0,     0,     1,    -3,    -2,     3,     4,    -7,     0,     4,     8,     2,    -1,    -2,    -2,    -7,    -5,    -6,    -1,     0,     0,    -2,    -4,    -1,     5,     3,     3,    -4,     0,     1,    -1,    -7,    -4,     0,    -2,    -8,    -5,     4,     5,     0,     4,     1,     0,    -1,    -3,    -1,    -1,     3,     1,    -1,    -3,    -3,     2,     7,    -5,    -1,    -1,     1,     1,     0,    -3,    -1,    -4,    -4,    -6,     0,     4,     4,     6,     3,     3,     3,     2,     0,    -1,     3,    -1,     2,    -6,     2,     1,     5,    -2,    -1,     1,    -1,     0,     0,    -6,     0,     0,    -2,     0,     2,    -1,     2,    -1,    -5,    -3,     0,    -2,     1,     0,    -5,    -6,     3,     0,     0,     1,    -1,    -1,    -1,    -1,     0,     0,     2,    -3,     0,     0,     3,     6,     0,     2,    -4,    -4,    -4,    -5,    -2,     0,     1,     5,    -6,    -7,     4,     1,     3,     3,     0,    -1,     0,     0,     0,     1,     0,     3,     1,    -1,    -2,     1,   -10,    -1,     5,     2,    -1,    -1,     7,    -2,    -8,    -6,    -3,    -5,    -1,     0,    -2,     2,     2,    -1,    -1,    -1,     0,     1,     1,    -1,    -2,    -2,     1,     1,    -2,    -3,    -1,     3,     0,    -2,     0,     4,     7,    -4,     1,     0,     1,    -2,    -1,     0,    -1,     1,     1,    -1),
		    80 => (    0,     1,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,     0,     1,    -1,     1,     1,     1,    -1,    -1,     1,     1,     0,     1,    -1,     0,     0,    -1,    -1,     1,    -1,     1,     1,     0,     1,     1,     0,     1,     0,    -1,    -1,     1,     1,     1,    -2,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     8,     7,     0,     1,     2,    -1,    -2,    -1,    -5,    -5,    -8,    -8,    -8,    -5,    -6,    -4,    -6,    -4,    -4,    -5,    -3,    -4,    -2,     0,    -1,    -1,     0,     1,     9,     6,     3,    -1,    -2,    -4,    -3,    -4,    -2,    -3,     3,     1,    -3,     1,    -1,    -2,    -1,     1,    -8,    -6,    -5,     0,    -1,    -4,    -1,     0,     0,    -1,     0,    -2,    -3,    -4,    -4,    -4,    -2,    -3,    -3,    -6,    -3,    -2,     1,    -3,     1,     4,     2,     5,     3,     9,    -3,     0,    -3,    -5,    -1,     0,     1,    -2,     2,     1,     0,     2,    -7,    -9,    -7,    -8,   -11,    -6,     0,    -1,    -1,    -2,     3,     3,     2,     6,     4,     9,    -2,    -1,    -3,    -5,    -2,    -1,     1,    -2,    -1,     1,     6,     1,     1,    -6,   -11,   -10,   -10,    -2,     5,     0,     1,    -7,    -3,     0,     1,    -1,     7,     5,    -5,    -8,   -10,    -6,     0,    -1,    -1,    -1,    -2,     3,     7,     1,    -2,    -4,    -3,    -4,     1,     0,     1,    -4,    -1,    -2,    -2,     0,     4,     2,    -4,     3,     2,    -2,    -2,    -7,     2,     3,    -2,     3,    -2,     1,     4,     3,    -3,    -4,    -5,    -8,    -7,    -3,    -3,     5,    -4,     2,    -1,     2,     1,     1,     4,     4,     3,    -5,    -7,    -7,    -1,     0,    -1,     4,    -1,    -3,     4,    -3,    -4,    -2,   -10,    -3,    -6,    -2,    -1,     4,     2,    -5,    -1,     2,     0,     2,    -1,     2,     5,     4,     1,    -5,     1,     0,     0,     2,     0,    -5,    -2,    -8,    -3,    -4,     1,    -4,    -1,     4,    -1,     1,     3,     0,    -4,    -8,    -3,     6,     4,     5,     5,     4,     2,    -9,    -1,    -1,     4,    -3,    -2,    -6,    -6,    -4,     4,     1,    -1,    -2,     1,     1,    -3,    -1,    -4,    -9,   -11,   -11,     0,     2,     2,     0,     0,    -1,     0,    -5,    -1,     1,     3,    -1,    -2,    -3,    -4,    -4,    -1,    -1,    -1,     3,     4,     4,     4,     2,    -2,   -16,   -15,    -4,     3,    -5,    -1,     2,     8,    -1,    -2,    -4,     0,     1,     3,     2,    -4,    -3,    -3,     0,     1,     1,     3,     1,     4,     2,     3,     0,    -4,   -20,    -7,     4,    -1,    -4,    -5,     1,    16,     5,     3,    -4,    -1,     0,     0,     0,   -10,    -3,    -1,     2,     5,     0,     2,    -5,     0,    -1,    -2,   -17,   -14,   -15,    -6,    -3,    -3,    -3,     2,     1,     7,     2,    -2,    -7,     0,     0,     1,    -2,   -11,     2,    -4,     1,     6,     2,     2,    -7,    -3,     4,    -1,   -12,    -8,    -2,     0,    -4,    -3,    -8,     1,     2,     4,     7,    -5,    -8,    -2,     1,     1,     0,    -8,     2,     0,     0,     5,     4,    -3,    -3,     1,    -5,    -8,    -3,    -1,     0,    -2,     2,    -4,    -2,    -4,    -2,     0,     4,    -6,    -4,     1,     0,    -1,    -4,    -4,     1,     5,     2,     6,    -3,     2,     0,    -4,   -11,    -8,    -5,    -1,    -4,     0,    -1,     2,     2,    -6,    -4,     1,     4,    -7,    -4,     1,    -1,     1,    -3,    -1,     2,     1,     2,     5,     7,     3,    -6,   -11,    -8,    -4,     0,     1,    -1,     0,     2,    -4,    -1,    -2,     2,     1,     1,    -3,    -2,    -2,     1,     2,    -7,    -2,     8,     0,     1,     4,     2,     3,    -5,   -10,    -4,    -5,     0,     2,    -4,     1,    -3,    -2,    -6,    -2,     2,     0,     3,    -5,    -1,     1,     0,     2,    -9,     2,     7,     1,     3,    -1,     3,     2,    -1,     2,    -2,    -3,    -1,    -7,    -1,    -2,    -2,    -7,    -7,    -3,     1,    -1,     1,    -4,     1,     1,     1,     1,    -9,     2,     1,     1,     4,     6,     1,     3,     0,     0,    -3,    -2,     0,     3,     0,    -1,    -5,    -6,    -9,    -9,    -5,    -2,     5,    -3,     1,     2,     1,    -1,   -10,     0,     0,     5,     6,     2,     2,     2,     2,    -3,    -4,     1,     4,     0,    -9,    -7,    -3,    -4,   -10,    -6,    -1,    -1,     4,     0,     0,     1,     1,     0,    -2,    -7,    -8,     1,     1,     0,     1,     4,     4,     4,     0,     3,     3,    -5,    -8,    -5,    -8,    -7,   -10,    -5,     2,     0,    -6,     0,    -1,    -1,     0,     0,    -2,    -2,     7,     9,     0,    -2,     1,     5,     8,     5,     7,    -8,    -7,    -7,   -14,   -12,    -7,    -7,    -4,     1,    -1,     0,     3,     1,     0,    -1,     1,    -1,     0,     0,    -5,    -9,    -9,    -9,    -8,    -5,    -6,    -8,   -10,    -7,    -3,    -8,    -9,    -8,   -10,    -7,     0,    -2,    -2,    -1,     0,     0,    -1,     0,     1,     1,    -1,    -1,    -1,    -7,   -10,    -2,     0,    -2,    -4,    -5,    -2,    -3,    -3,    -5,    -5,    -9,   -10,    -2,    -6,    -2,    -2,    -1,     0,     1,    -1,     1,    -1,    -1,     1,     1,     0,     1,     1,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     0,     1,     0,    -2,    -1,    -2,    -2,    -1,     0,     0,     1,    -1),
		    81 => (   -1,     1,     1,     1,    -1,    -1,     0,    -1,    -1,     1,    -1,     1,     0,     0,     1,     0,     0,     0,     1,     0,     1,     0,     1,     0,    -1,     1,    -1,     1,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,    -2,     1,     2,    -1,    -2,     0,    -1,     0,     0,    -1,     1,     1,     0,     1,    -1,    -1,     1,    -1,     1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     6,     8,    16,    12,     6,    -4,     1,    -5,    -4,    -3,     0,     1,     1,    -1,     0,     0,     3,     2,    -1,    -4,    -9,    -3,     6,     2,    -4,    -6,    -5,    -1,     3,     9,    10,     2,     0,    -4,     0,     6,    -1,     0,    -4,     0,     1,     0,     1,     1,     3,     3,     6,     3,    -2,    -2,     9,     7,     4,    -1,    -1,    -4,    -1,     2,     3,     2,    -2,    -2,     4,     6,     3,     4,    -1,    -3,    -3,    -4,     0,    -1,    -1,    -1,     7,    13,     6,     5,     3,     1,     1,    -7,    -7,     1,     4,     1,    -2,     1,     0,     2,     4,     4,     4,     1,     1,    -1,    -4,    -4,     1,     1,    -8,     1,     1,     3,     6,     2,    -4,    -5,     3,    -1,     0,    -1,    -1,    -1,    -5,     4,     2,     6,     3,    -1,     2,    -1,    -1,    -1,    -2,    -1,    -1,     1,    -9,    -8,    -8,     0,     3,     4,    -6,     1,     4,    -4,    -1,    -5,    -1,     4,    -1,     1,     3,     7,     1,    -1,     2,    -2,    -2,     0,    -4,    -2,     0,    -1,   -11,    -6,    -8,    -1,     2,     0,    -2,     3,     2,     1,     3,    -5,    -5,     1,     4,     0,     4,    -5,    -3,    -3,     1,    -3,     0,     0,    -4,    -1,     1,     0,   -10,    -4,    -5,    -5,     0,     3,     4,     1,     1,     8,     6,    -4,    -7,    -2,    -4,    -4,    -4,    -3,    -2,    -3,    -4,     0,    -1,     1,     1,    -1,     0,     0,    -8,    -1,    -9,    -5,    -8,     1,     3,     5,     2,     8,     2,    -2,    -3,    -2,    -5,    -4,    -2,    -7,    -5,    -5,     0,    -1,    -2,    -1,     1,     0,     0,     2,    -2,    -1,    -7,    -4,    -7,     0,    -3,     2,     1,     4,     2,    -2,    -1,    -5,     1,    -6,    -5,    -7,    -4,    -3,     1,     0,    -1,    -1,    -1,     1,    -1,    -1,    -1,    -3,    -5,    -5,     2,     5,     1,     0,    -2,     1,     0,    -4,    -5,    -1,    -2,    -6,    -2,    -7,   -10,    -4,    -2,    -2,    -1,    -2,     1,     2,     0,     0,    -1,    -1,    -7,     3,     5,     5,     6,    -3,    -4,     0,    -1,    -6,    -2,     3,    -2,    -4,    -5,   -14,    -7,    -6,    -5,    -4,    -4,     0,     0,     0,    -1,     0,     1,     0,    -6,     5,     4,    -1,    -2,    -8,   -11,    -6,    -4,    -3,     2,     2,     0,    -4,    -6,   -10,    -8,   -10,    -6,    -4,    -2,    -4,     0,     1,    -1,     1,     0,     2,    -1,    -5,    -3,    -3,    -6,    -7,    -9,   -10,   -11,    -1,     5,     1,    -1,    -4,    -6,   -13,    -7,    -8,    -6,    -6,   -14,    -2,    -1,    -2,     1,     0,     2,    -3,    -3,    -3,    -4,    -4,   -10,    -5,    -6,   -10,    -9,    -1,     6,     5,    -1,    -5,    -5,   -10,    -8,   -10,    -4,    -7,    -5,    -2,    -1,    -2,    -1,    -1,    -1,    -5,    -1,    -2,    -4,    -7,    -7,    -7,    -8,   -17,   -10,    -8,     3,    -3,    -2,    -3,     0,    -4,    -5,    -4,     0,    -4,    -8,    -8,    -1,    -3,    -2,     1,     1,    -1,    -1,    -6,   -12,    -7,   -12,    -8,    -9,   -22,   -19,   -11,     0,    -4,    -2,     2,    -2,    -2,     4,     3,     6,    -3,   -14,    -3,    -3,    -3,     0,     0,    -1,    -3,    -4,   -11,    -6,    -1,    -1,    -4,    -6,   -10,    -7,    -5,    -4,     3,     5,     1,    -5,     0,     2,     0,    -1,     3,    -1,    -1,    -5,    -1,     1,    -1,    -3,     4,     0,    -8,    -4,     1,     2,     4,     7,     1,    -2,     1,     3,     2,     7,     4,    10,     7,     6,     0,     2,     3,     2,     1,    -4,     1,     3,     1,    -4,     4,     5,     2,     6,     5,     6,     6,     3,     3,     0,     2,     2,     6,     1,     6,     9,     3,     3,    -1,    -5,    -3,     2,     4,    -5,     1,     3,     1,   -12,    -7,     4,     9,     3,     1,     1,     3,     3,     2,     1,     2,    -1,     2,    -2,     2,     1,     5,     5,     3,    -9,    -6,     1,    -1,     0,     0,     1,     1,    -1,    -3,     2,    -2,     3,    -1,    -1,    -2,    -3,     1,     0,     4,    -4,    -7,    -9,    -8,    -3,     2,     4,     5,    -2,    -5,    -5,    -6,     3,     1,     0,     0,    -1,     0,    -2,    -3,    -5,    -1,     1,     3,    -1,    -1,    -9,    -6,   -11,    -9,    -9,    -5,    -3,    -1,     1,     2,    -3,    -4,    -6,    -1,     0,     1,     0,    -1,     1,    -1,     0,    -1,    -2,    -1,    -1,    -6,    -2,    -4,    -5,    -6,    -4,    -8,    -6,    -6,    -8,    -6,    -8,    -6,    -5,    -2,     0,     1,     0,    -1,    -1,     1,    -1,     0,    -2,    -2,    -2,    -2,    -1,    -5,     0,    -1,    -3,    -4,    -3,    -5,    -1,    -5,    -3,    -4,    -3,    -3,    -2,     0,    -1,    -1,     1,    -1,     1,    -1,     0,    -1,     0,     1,     0,     0,     0,    -1,    -2,    -2,     0,    -2,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,     1),
		    82 => (    0,     0,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,    -1,     0,     2,     1,     0,     0,    -1,     1,     0,    -1,     1,     0,    -1,     1,     0,     0,     0,     1,     1,     0,    -1,     1,     1,    -3,    -5,    -2,    -4,    -4,    -5,    -9,    -4,     1,     4,     1,    -5,    -9,    -6,    -3,    -5,    -2,     0,    -1,     0,     0,     1,     1,     0,    -7,    -7,     1,     0,    -1,     0,     8,     7,     3,     2,     2,     1,     3,     0,    -1,    -4,    -6,    -4,    -3,    -2,     0,     1,     1,     0,     0,     0,    -1,     0,    -7,    -9,    -1,     0,     2,    -3,     3,     1,     1,    -2,     2,     5,     3,     3,     1,    -3,    -4,    -3,     1,    -5,   -12,     1,     2,     1,     0,     0,     1,    -2,     2,     2,    -3,     1,    -1,    -6,     3,     6,     1,     1,     4,     5,     2,     3,     1,     6,     1,     0,    -2,    -6,    -3,    -4,    -1,    -3,     0,     0,    -1,     2,    -1,    -1,     2,     2,    -6,    -1,     2,    -4,    -3,     2,     0,     0,    -1,     4,    -2,     1,    -3,    -2,    -2,    -4,    -2,    -8,     0,    -3,    -3,     0,     0,     1,    -3,    -3,     1,     0,     5,    -4,    -4,     1,    -2,    -5,     5,     0,     1,     6,     1,     2,    -5,    -3,     0,    -3,    -4,   -10,     4,    -2,    -1,    -1,     1,    -1,    -3,    -3,    -1,     3,     0,    -4,    -4,     3,     1,     0,    -4,     0,     3,     0,     1,    -7,    -1,     3,     4,    -1,   -10,    -4,     1,    -5,    -2,    -2,     2,    -2,    -4,    -2,    -6,    -4,     0,     3,     2,     5,     3,    -6,    -3,    -7,     0,     0,     1,     2,     5,     0,     1,     0,    -5,    -8,   -10,    -4,    -2,     0,    -2,    -1,    -3,    -2,    -8,    -7,    -9,   -11,    -3,     0,    -6,    -9,     0,    -1,    -5,    -1,     2,     3,    -4,    -2,     5,     0,    -4,    -4,    -5,    -3,    -3,    -1,     0,    -1,    -6,    -6,    -8,    -9,   -17,   -24,   -22,   -18,   -14,    -4,    -5,    -1,    -6,     0,    -2,     2,     0,     0,    -2,     0,    -2,    -7,    -6,    -3,    -1,     0,    -3,    -3,    -7,    -7,    -8,   -12,   -15,   -20,   -17,   -14,    -8,    -6,    -8,    -2,    -5,    -4,    -9,    -9,     0,     0,     1,     3,    -2,    -7,    -1,    -3,    -2,     1,    -4,    -8,    -6,   -10,    -8,    -7,    -9,    -3,    -2,    -1,     2,    -1,    -2,     1,    -4,    -6,    -8,    -6,    -3,    -2,     2,     5,    -6,    -6,     7,     1,    -2,    -1,    -4,     0,    -2,    -5,    -4,     1,     9,     4,    -1,    -2,     2,     9,     6,     2,     1,     0,     0,    -3,    -4,    -1,     3,     7,    -1,    -1,     3,     0,     0,     0,    -4,    -5,     6,     4,    -1,     6,     9,     8,     5,     8,     6,     5,     8,     7,    -1,     4,    -7,    -4,    -1,     3,    -1,     1,     1,    -1,     4,     4,     3,     0,    -2,     1,    15,     6,     8,     5,     4,     4,     4,     7,     2,     4,     2,    -3,     2,    -1,     1,    -3,     0,    -4,    -2,    -1,     4,    -1,     6,    11,     7,     0,     0,     1,     6,    -2,     8,    12,     5,     2,     4,     4,     1,    -4,     3,     3,     2,     2,     2,    -1,     0,    -4,    -4,    -2,    -2,    -5,     8,    11,     4,     1,    -2,     1,    -3,     3,     2,     8,    -2,     4,    -3,    -4,     2,     0,    -1,     6,     4,     4,     1,     0,    -4,    -1,    -9,    -6,    -7,    -9,     1,     3,     7,     1,    -1,    -5,     1,     0,     6,     6,     0,     0,    -3,    -4,    -2,     0,     2,    -1,     0,     4,     1,     4,     5,     3,    -2,    -4,    -4,     1,     6,     3,     7,     0,    -4,    -4,    -2,     4,     3,     4,     4,     2,     1,    -3,     1,     0,    -1,    -4,    -1,     1,     0,     4,     5,     1,     4,     4,     2,     7,     6,     5,     4,    -1,    -5,     0,    -1,     3,     8,     3,     0,    -1,    -4,    -3,    -5,    -7,    -6,    -6,    -1,     0,    -5,    -3,    -1,    -2,     0,    -2,     1,     8,    -1,     2,     0,    -1,     3,     0,     2,     3,     2,     2,     2,     3,    -4,    -5,    -1,    -1,    -6,    -4,    -4,    -4,    -1,    -4,     0,     3,     5,     2,     4,     2,    -4,    -3,    -1,    -1,    -1,    -1,     2,     4,    -4,    -3,    -2,    -1,    -4,    -1,     1,    -2,    -5,    -7,    -3,    -5,    -5,    -7,    -1,     0,     1,    -2,    -2,    -3,    -7,    -8,    -1,    -1,    -1,     2,     6,     6,     1,    -6,    -1,    -4,    -8,    -2,    -5,    -1,    -9,    -5,    -8,    -3,    -4,    -6,   -10,    -5,     0,     4,    -6,    -6,    -4,    -5,     1,     0,     1,    -3,    -2,    -2,    -1,    -2,    -5,    -6,   -10,   -12,    -9,    -7,   -11,    -8,    -7,    -7,    -3,    -4,   -10,   -12,    -7,   -11,    -7,     2,     3,     3,     0,     0,     0,    -2,     0,    -2,    -2,    -2,    -3,    -7,    -9,    -3,    -2,    -3,    -8,    -6,    -4,    -6,    -8,    -5,   -10,    -8,    -5,    -6,    -2,    -2,     2,     4,     0,     0,     1,    -1,     0,    -2,    -3,    -3,    -2,    -3,    -1,    -1,    -1,     0,     0,    -3,    -2,    -8,    -6,    -5,    -3,    -2,    -2,    -1,    -2,     1,     0,    -1,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,     0,     1,    -2,    -1,    -1,    -2,     0,    -1,    -1,     0,    -2,    -2,    -3,    -4,    -2,    -1,     0,     0,    -1,    -1),
		    83 => (    1,     0,     1,     1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -2,    -2,     0,     0,     1,     0,     1,     0,     1,     1,     0,    -1,     1,     1,     0,     1,     0,    -1,     1,    -1,     0,    -1,    -1,     0,    -2,    -1,    -2,    -5,    -4,    -4,    -2,    -6,    -3,    -3,    -2,    -1,    -1,     0,     1,     1,    -1,    -1,     0,     0,     0,     0,    -3,    -2,    -3,    -3,    -6,    -8,     3,     0,    -3,    -5,    -7,    -6,    -4,    -1,     1,    -6,    -8,   -10,    -9,    -7,    -1,     1,    -1,     0,    -1,     1,    -1,    -2,    -1,     3,     5,    14,    13,     5,     6,     6,     4,     2,    -1,     7,     9,     6,     5,    12,    21,     2,   -13,   -13,    -7,    -4,     0,     0,     1,    -1,    -8,     0,     3,     4,     2,     9,    11,     0,     6,     3,     3,    -1,     2,     0,     4,     6,     5,     5,     2,    -7,    -7,   -26,   -20,    -8,    -5,     1,     0,     1,    -1,    -1,    -1,     4,    10,    12,     1,     3,     5,    -2,    -4,     1,    -2,    -1,     6,    -3,    -1,     4,     1,    -2,    -2,     2,     2,   -10,    -5,     1,     1,     1,     3,     0,    -1,     9,    13,    11,     5,     5,     2,     0,    -3,     2,    -1,     4,     3,     1,     1,    -1,     1,    -2,     0,     1,     4,   -12,    -5,    -2,     0,     1,     0,     2,    -1,     2,    12,    16,     8,     1,     1,     7,     1,    -4,     1,     0,     3,    -2,    -4,     2,    -2,    -2,    -3,    -1,     4,   -10,    -7,    -3,    -4,    -1,    -5,     0,     2,     9,     2,     4,     1,    -2,    -2,    -6,    -7,    -4,    -2,     7,     3,     4,    -5,     3,     1,    -4,     3,     0,    -3,    -7,    -6,     0,     0,    -3,   -12,    -3,    13,    12,     5,     6,     6,    -3,     2,    -4,    -3,    -2,    -3,    -3,     1,     7,     3,    -1,     2,    -3,     7,     6,   -14,    -6,    -4,     1,    -1,     0,   -13,     1,     3,     6,     8,    10,     0,    -3,    -6,    -7,    -4,    -6,    -2,    -3,    -1,     4,     5,     2,    -6,    -4,     2,     9,    -6,    -7,    -5,     0,    -1,    -5,    -6,     7,    11,    10,     6,     2,     5,    -3,    -1,    -6,    -6,    -2,     0,    -5,     1,     1,     3,    -5,    -7,    -3,     0,    -3,   -17,   -12,    -6,    -1,    -1,    -1,    -6,     3,     7,    10,     7,     4,     1,    -4,     2,    -3,    -4,    -4,    -4,     1,     1,     0,     1,     2,    -4,    -8,    -3,     1,   -11,    -7,    -3,    -1,     1,    -2,    -5,     0,    11,     8,     5,     4,     8,    -1,     3,    -3,    -4,    -1,    -2,     5,   -12,    -3,     5,     5,    -4,    -4,    -5,     3,    -2,   -12,    -3,    -1,     0,     3,    -1,     3,     5,     8,     8,    -1,     3,     0,    -2,    -1,     0,    -3,     2,    -5,    -6,    -1,     3,     3,     2,     2,    -2,     3,    -2,   -16,    -7,     1,    -1,     3,    -3,     2,     4,    10,     6,    -6,    -3,    -6,    -1,    -4,    -2,    -5,    -4,    -2,    -5,    -6,    -2,     6,     1,     2,     4,     7,     8,   -17,     3,    -3,     1,     0,     1,    11,    10,     8,     1,     3,    -8,     0,     1,    -6,   -10,    -2,     1,    -3,    -6,    -4,     5,     8,     1,    -3,     4,     1,     5,   -19,    -8,    -4,     0,     2,    -2,     5,     7,     2,    -2,     1,    -3,    -2,    -4,    -4,     0,     0,    -6,    -4,     2,     2,     4,     7,    -1,     1,    -4,    -3,    -4,   -15,    -5,    -2,    -3,     2,    -1,     3,     8,     6,     0,     0,    -2,    -6,     0,    -2,    -5,     5,     0,     5,     0,     3,     8,    -4,     2,    -3,    -2,    -9,    -3,   -15,    -1,    -4,    -1,    -2,     3,     2,     3,     6,    -3,    -4,    -5,    -9,    -5,    -5,    -1,     2,     6,     5,     0,     5,     4,    -2,     2,    -1,    -2,    -4,     2,    -8,    -6,    -5,    -1,     2,    -6,     1,     3,     4,     0,    -2,    -5,     0,    -4,    -4,    -2,     0,     5,     3,    10,     7,    -1,    -2,     4,     3,     4,     4,    -1,   -10,    -5,     0,    -1,    -1,     3,    -1,     1,    -5,     4,     7,     0,    -2,    -4,     0,     2,     5,     7,     8,     5,     2,     3,     7,    -1,     4,     6,    -2,    -8,   -10,    -5,    -1,    -1,     0,     5,     4,    -6,     3,     7,     8,    -2,     1,     4,     2,    -3,     2,     4,     2,    -3,     3,    -2,     5,     1,     5,    11,     2,    -6,    -7,    -4,    -1,     1,     1,     2,     1,    -3,    -2,     3,     7,     3,     2,     1,     4,     0,    -2,    -2,     3,     3,    -1,    -3,    -5,     0,    11,    10,     5,     9,     4,    -6,     1,     0,     0,     6,    10,     9,     0,     7,     6,     4,     8,     3,    -2,    -2,     1,     3,    -2,     0,     1,    -5,     2,    14,     9,     5,     6,    -9,    -5,    -2,     0,     1,     0,     1,    -3,     0,     8,     7,    -1,     3,     3,    -4,    -2,     3,     9,     1,    -1,    -1,     2,     4,     5,    -4,   -11,   -12,   -12,   -10,    -3,    -2,    -1,     0,     1,     0,    -2,   -12,     5,     3,     1,     4,    -3,    -2,    -5,    -5,    -3,    -4,     0,    11,    12,    11,     2,    -2,    -5,   -13,    -6,    -1,    -1,     0,     1,     0,    -1,     1,     1,    -2,    -4,    -3,    -2,    -3,    -8,    -7,    -6,    -5,    -7,    -7,    -4,    -1,    -2,    -1,    -6,    -7,    -2,    -2,    -2,     1,     1,     1,     1),
		    84 => (    0,     0,     1,     1,     1,     0,     0,     0,     1,     0,     0,     0,    -4,    -2,    -1,    -2,     0,     0,     1,    -1,     1,     0,     1,     0,     0,     1,     0,    -1,     1,    -1,     0,    -1,    -1,    -2,    -4,    -5,    -3,    -5,    -5,    -5,    -6,    -6,    -1,    -6,    -5,    -1,    -3,    -3,    -5,    -4,    -2,    -5,     0,     1,     1,    -1,     1,     1,    -3,    -5,    -6,    -8,    -7,    -7,   -11,   -10,   -14,   -15,     1,     3,     0,    -8,    -7,    -9,   -13,    -7,   -15,    -7,    -7,    -5,    -3,    -3,     1,     1,     1,     0,    -1,   -13,    -9,    -9,    -5,    -8,    -6,   -12,   -11,   -11,    -7,   -15,    -2,    -1,    -7,    -4,    -4,    -1,     5,     0,    -7,    -8,    -4,    -3,    -1,     0,     1,     1,    -6,   -13,    -1,     0,     3,     0,    -6,     0,    -2,    -9,    -1,    -2,    -4,    -6,    -3,    -1,    -2,     1,     0,    -4,     1,     2,     3,    -2,    -9,    -1,    -1,    -1,    -7,    -1,     0,    -2,    -1,    -1,     3,    -2,     5,     0,     5,    -4,    -3,    -6,    -4,     3,    -1,     1,    -6,    -2,     1,    -1,    -3,     3,    -3,     0,     0,     1,    -3,    -5,     3,     7,     4,    -6,    -2,    -7,    -1,     2,     0,    -4,   -10,   -10,    -8,    -6,    -8,    -5,   -10,     0,    -1,    -1,    -2,    -1,     0,    -4,     1,   -12,    -4,     0,     3,     5,    -5,    -6,    -9,    -4,    -2,    -1,    -7,    -5,    -7,    -9,    -8,    -2,    -5,    -6,    -5,    -4,    -4,    -3,     2,     6,     5,    -7,    -4,   -10,     7,     2,     5,     2,    -9,    -9,   -10,    -4,    -9,    -6,    -4,    -1,   -12,    -7,    -7,    -2,    -3,    -1,    -5,    -6,    -4,    -1,     5,     5,     0,    -2,     0,    -8,     6,     2,    -4,     0,    -6,    -4,    -5,    -5,    -8,    -2,     0,    -3,    -7,    -3,    -4,    -2,     0,     3,     2,     6,     3,     4,     6,    -4,    -8,    -2,     1,    -5,     4,     1,    -3,     4,    -2,    -6,    -3,    -1,     0,     0,     5,    -2,    -3,     5,     4,     8,    -2,     0,     3,     2,     2,    -1,    -1,     1,    -4,    -2,    -1,    -6,    -1,     0,     0,     7,     0,     0,     2,     8,     6,     4,     8,    -2,     1,     5,     8,     2,    -3,    -2,     0,     1,     3,     3,    -1,    -2,    -8,    -8,     0,    -1,     4,     4,    -1,     5,     4,     3,     5,     6,     6,     5,     7,     3,    -2,    -1,     1,    -1,    -4,    -1,    -1,     3,     6,     3,     9,     5,     4,    -9,     1,    -1,    -1,     7,     3,     6,     3,     5,     0,     3,     4,     9,     8,     5,     0,    -3,     4,     3,    -5,     1,     1,     6,     4,     5,     4,    11,    11,    -5,     1,     2,   -11,     3,    10,     7,     4,     3,     6,     4,     3,     3,     6,     0,    -2,    -3,     5,     8,    -4,     6,    -3,     7,     4,    -3,     0,     7,     7,    -1,    -1,     2,    11,     5,     0,     6,     2,    -3,     1,     3,     4,     3,     2,     1,    -1,     4,     7,     1,     0,     6,    -1,     0,     7,     4,    -3,     5,    13,    -2,     0,     1,    -2,     7,     2,     5,     7,     5,     4,     1,    -1,    -2,     2,     0,    -1,     8,     3,     4,     7,    10,     3,     1,     0,     0,    -1,     4,     8,    -3,    -1,    -2,     3,    -3,     9,     7,     3,     4,     1,     1,     0,     0,     0,     3,     2,     2,     4,     1,     1,     4,    -4,     0,     2,     2,     2,     1,     5,     0,    -7,     0,     7,     3,     7,     0,    -2,    -2,     2,     4,     0,     3,     1,     5,     6,     1,     1,     2,     3,    -2,    -2,     0,    -1,    -4,    -2,    -7,    -2,    -3,     0,    -5,    -4,     9,    -1,     7,     1,    -6,     3,     1,    -3,     1,     0,    -2,     4,     1,    -3,    -3,    -4,    -8,    -6,    -5,    -8,    -9,    -2,    -6,    -3,    -3,     0,    -1,    -6,     6,     3,     0,     1,     0,     1,    -5,   -12,    -6,    -8,    -4,    -2,    -5,    -2,    -6,    -8,    -7,   -12,    -9,    -6,    -8,    -3,   -13,    -2,     0,     0,    -2,   -10,     3,     4,     1,    -6,    -9,    -3,    -5,    -8,    -5,    -7,    -5,    -8,    -4,     0,    -3,    -5,    -8,    -3,    -7,    -3,    -6,     1,    -8,    -8,    -1,    -1,     0,     0,    -7,   -11,    -2,     0,    -9,   -10,    -9,    -2,    -3,    -6,    -7,    -4,    -2,    -5,    -6,    -4,    -2,    -6,     1,     1,     4,    -4,    -3,    -1,    -2,    -1,     0,     0,   -10,    -5,   -12,     0,     3,     1,    -7,     3,    -3,    -3,    -3,    -4,    -2,    -3,     0,    -4,    -1,    -4,     2,    -2,    -6,    -8,     1,     0,     1,     0,     0,     0,    -1,    -9,    -1,     3,     4,     4,     2,    -5,    -1,    -8,     3,     4,    -4,     0,    -4,   -10,    -6,    -1,     3,    -1,    -5,   -14,    -2,    -3,     1,     0,    -1,    -3,    -2,     2,    -7,     2,     0,    -3,    -6,    -2,    -3,    -8,    -7,    -3,   -10,    -2,    -4,    -5,    -8,    -2,    -1,     3,    -1,    -9,    -4,    -3,     0,     1,     1,     0,    -7,    -3,    -2,    -8,    -9,    -4,    -4,   -13,    -9,    -6,   -13,   -12,    -8,   -11,    -4,    -3,   -12,   -17,   -16,   -15,    -4,    -4,    -1,    -1,    -1,     1,     0,     1,    -1,    -1,    -2,    -1,    -2,    -3,    -3,   -10,   -11,    -6,    -8,   -10,    -3,    -5,   -11,    -7,    -8,   -10,    -7,    -7,    -2,     1,    -1,     1,    -1),
		    85 => (    0,     0,     1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,     0,     1,     1,    -1,     0,     0,    -1,    -1,     0,     0,     1,     0,    -1,    -1,    -1,     1,     0,    -1,    -1,    -1,    -1,     1,     0,     1,    -2,    -5,    -4,    -5,    -4,    -4,    -5,    -5,    -6,    -8,    -4,    -4,    -2,    -1,    -1,     0,     0,     0,     0,     1,    -2,    -2,    -2,    -2,    -3,    -2,   -12,    -9,   -14,   -12,   -10,   -10,   -10,    -2,    -1,     2,     3,    -2,     3,     1,    -1,     3,    -5,    -2,     1,     1,     0,     1,    -4,     4,     6,    -4,   -13,   -11,    -2,     1,     4,    -7,    -8,    -1,    -5,     7,     5,     3,    10,     8,     8,    16,    13,     9,    -4,     4,     3,     0,     0,     0,    -4,     4,   -14,   -12,    -7,    -4,   -13,    -4,     4,    -3,    -3,    -6,     2,     6,     6,    10,    18,     9,     9,    11,    19,     9,    -6,     1,    -4,    -3,     0,     1,    -6,     6,   -15,    -5,    -4,    -4,     0,     4,     5,     1,    -4,    -7,     3,     3,     6,     9,    11,    11,    14,     3,     9,     3,    -4,    -4,    -6,    -7,     0,     0,    -1,   -14,    -2,     7,     7,     3,     6,     3,     3,     0,     0,    -6,    -1,     0,     2,     0,     8,    13,     8,     0,     7,     6,    10,     9,     2,     2,     0,    -2,    -1,   -16,    -9,    -3,     3,     1,     1,     0,     0,     6,    -5,    -3,    -3,   -10,    -2,    -3,     6,    10,     3,     5,    15,    12,    11,     3,     5,     9,    -4,    -5,    -7,   -16,    -5,    -6,     2,     4,    -1,     0,    -5,     2,     4,     0,    -4,    -7,    -9,    -2,    -3,     9,     7,     7,    13,    11,     7,     1,     4,     6,     1,     0,    -7,    -9,    -4,    -4,    -2,     3,     2,    -4,     1,     1,    -1,     0,    -6,   -10,   -10,    -7,    -2,     8,     1,     2,     7,     9,     9,     5,     1,     0,    -1,    -2,    -4,   -14,     3,     0,    -6,    -6,     0,     3,    -6,     4,     4,    -3,    -6,    -4,   -11,    -9,     3,     1,     2,     7,     6,    10,    12,     2,    -3,    -3,    -1,    -1,     0,   -10,     2,    -5,     0,    -5,     1,    -2,    -3,     0,     1,    -3,    -7,    -4,     4,     2,     0,     1,    -5,    -2,     5,     8,    11,     7,    -4,    -3,     0,     0,    -2,    -7,     9,    -1,    -2,     4,     3,     5,    10,     1,     7,    -2,    -2,    -6,    -1,    -3,    -1,    -6,    -6,    -5,     0,     2,     3,     8,    12,    -4,     1,    -1,    -1,    -9,     1,     1,    -2,     6,     0,     0,     3,     4,     6,    -2,    -4,    -1,    -2,    -5,    -7,     2,    -2,     5,    -5,    -8,    -8,    -5,     9,    -4,     0,     0,    -3,   -10,     5,     3,     8,    -1,     0,     5,     5,     4,    -3,     1,     2,    -1,     0,    -3,     2,     0,     5,    -1,     4,     0,    -2,   -10,   -10,    -4,     2,     0,    -6,    -2,     7,     9,     1,     4,    -2,     2,     4,    -1,    -2,     1,    -2,    -9,    -3,     1,    -2,    -1,    -2,    -1,     1,     3,     2,    -4,    -8,    -2,     0,    -1,    -7,    -2,     3,     8,    11,     4,     1,     2,    -3,    -3,    -5,     0,    -2,    -5,    -8,     0,     5,     1,    -4,     4,     6,    -1,    -6,   -12,   -11,    -3,     0,    -2,    -9,    -2,     6,    11,     4,    13,     7,     0,    -1,    -2,   -10,    -2,     2,    -5,    -3,    -4,     1,     1,     4,     1,     5,     0,    -4,   -13,   -19,   -12,    -2,    -1,    -9,     0,     2,     3,    11,     9,     9,     4,    -6,    -2,    -8,    -9,     3,     2,    -2,    -7,    -2,    -2,     5,    -1,    -1,     1,    -6,   -12,   -11,   -10,     1,    -3,     5,     7,     1,     7,    10,     5,     0,     1,     1,     2,    -4,    -7,     2,     4,     2,     2,    -3,     0,    -5,     3,    -1,     4,     4,    -2,   -13,    -7,    -1,    -2,     8,     6,     7,    14,     6,     0,     3,     6,     1,     3,    -2,     2,     0,     7,     2,     2,     2,     2,    -2,     0,     0,     4,    -5,     2,   -15,     1,     0,    -2,    -7,    -1,     4,     9,    14,     3,    -3,     1,    -2,    -3,     1,     1,    -1,    -3,     0,     0,     3,    -1,     1,     3,     2,     1,    -3,     2,     2,     0,     0,    -1,   -12,    -6,    -1,     1,    -2,     6,     0,     2,    -1,     3,    -2,    -3,     5,     3,     3,     5,    -1,     6,     3,    -1,    -4,     1,     1,     4,     9,    -1,    -1,    -1,     4,    -2,     2,     0,     3,     2,    -2,    -2,     7,     3,     4,     6,     4,     4,     3,     2,   -10,    -4,     1,    -2,    -6,    -1,     6,     5,    11,    -1,     0,    -1,    -7,    -4,    -8,    -1,     0,     0,     4,     5,     2,     2,     4,     6,     6,     4,     6,     2,     3,     0,    -2,    -2,    -2,    -7,     2,   -11,    -5,    -1,     0,    -1,    -2,     6,   -12,   -12,     0,    -2,     1,    -2,    -1,    -1,     0,     2,    -4,     6,     7,     6,     2,     7,     6,     6,    11,    10,     8,    -3,    -1,    -1,     0,     1,     0,    -4,    -7,    -9,   -11,   -16,    -8,    -3,    -2,     3,     6,    16,     8,    11,     3,     1,    -3,     3,     0,     0,     0,    -9,    -3,     0,     0,     0,    -1,    -1,    -1,     0,     1,     2,    -1,    -2,    -3,    -2,     1,     0,     1,    -1,   -13,    -6,    -2,    -1,    -4,    -3,    -8,   -10,    -7,    -6,    -1,     1,    -1,     1),
		    86 => (    0,     0,    -1,     1,     1,     0,     1,    -1,     0,     0,     1,     1,     4,     3,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     4,     5,     4,     5,     5,     2,     6,     4,    -7,     0,    -1,     4,     3,     5,     6,     2,     1,    -1,    -1,     1,     0,    -1,     0,    -1,     2,    -1,     3,     1,     5,     3,     5,     7,     4,     3,     6,     3,     2,     0,     4,     4,     6,     7,    11,     9,     7,     3,     1,     3,    -1,    -1,    -1,    -1,    -4,    -1,     1,     4,     8,    10,     9,     9,    10,     8,     5,     7,     5,    -2,     1,     7,     6,     0,     2,     8,     9,     9,     6,    -2,     0,     0,     0,     1,    -9,    -4,     4,     8,    10,     7,     3,     6,     9,     5,     7,    -1,     2,    -3,     4,     5,     1,     3,     8,    -3,     0,     4,     4,     4,    -1,     3,    -1,     0,    -6,    -5,     5,     6,     4,     5,     6,     7,     9,     3,     5,     0,     1,     0,     5,     2,    -5,    -3,     1,    -2,     4,     4,     5,     8,     3,     2,    -1,     0,     0,    -2,     5,     1,     6,     2,     1,     7,     9,     3,    -3,    -3,    -3,    -2,     1,    -2,     2,     1,     1,     6,     2,     3,     3,     3,    -1,    -2,     0,     1,    -1,    -4,     2,     2,     1,     7,     5,     8,     4,     1,     0,    -4,    -1,    -3,     0,     2,     8,     2,     5,     2,    -2,    -4,     2,    -1,    -3,    -6,    -1,    -1,    -4,    -6,     6,     2,    -2,     2,     4,     4,     4,     0,     2,    -4,     2,    -3,    -4,     8,    -4,     2,     4,     8,    -6,    -8,    -8,   -12,    -7,   -10,     1,    -1,    -6,    -6,     2,    -1,    -2,     1,     3,     0,     0,     3,     1,    -1,     0,    -3,    -5,    -8,    -5,     3,     4,    -2,    -7,    -6,    -2,   -10,    -4,    -9,     0,     0,    -5,    -7,     2,    -3,    -3,    -3,    -2,     1,     1,    -3,     2,     1,     1,    -6,    -8,    -9,    -5,     3,     0,    -4,    -8,    -8,    -8,    -3,    -4,   -12,     0,     0,    -4,   -10,    -1,    -1,     0,    -5,    -8,    -3,    -1,     2,     3,    -2,    -5,    -4,    -3,    -3,     3,     3,     0,    -3,    -6,    -3,    -5,    -3,    -9,    -4,    -1,     0,    -1,    -6,    -1,     1,    -2,    -5,   -12,    -1,    -1,     1,     0,    -1,    -2,     0,     3,     9,     8,     2,    -3,     2,    -4,     7,     3,    -3,    -9,    -3,    -1,     0,    -2,    -6,    -1,    -3,    -4,   -12,   -15,    -5,    -2,    -1,    -3,     1,    -3,     2,     5,    -3,    -1,     3,    -3,     2,     0,     9,    -5,    -5,    -8,    -1,    -1,     0,    -1,    -7,    -6,    -3,    -8,    -7,    -9,    -5,    -1,     0,     0,    -1,     0,     2,     1,    -3,    -6,    -3,    -3,     0,     3,     7,    -1,    -1,    -1,     0,     1,    -1,    -2,    -6,    -9,    -5,    -5,    -2,   -13,   -11,    -5,     0,    -1,    -2,    -3,     3,     2,    -5,    -4,     1,    -2,     0,     1,     0,     0,     3,    -6,   -10,     1,    -1,    -3,   -11,    -2,     3,    -5,    -1,   -10,    -5,    -2,    -1,    -3,    -6,    -3,     0,     2,     0,     2,    -1,    -1,     1,     1,     1,     2,     2,    -6,    -9,     0,     0,    -3,   -10,     2,    -3,     0,     2,    -1,     1,     2,     4,    -3,    -7,    -5,    -2,     1,    -1,     3,     1,    -1,    -2,     0,     5,     6,     4,    -5,   -11,     0,    -1,    -2,   -12,    -2,    -4,    -1,     1,     1,     5,     8,     7,     4,    -2,    -1,     2,     2,     5,     5,     2,     4,     4,    -2,     3,     4,     6,    -5,    -5,     1,    -3,   -10,    -9,     0,    -3,     4,     5,     6,     1,    11,    10,     7,     2,     3,     0,     0,    -2,    -1,     2,     2,     0,    -1,    -1,     1,     0,    -3,    -2,     1,    -3,    -3,    -7,    -3,    -3,    -4,    10,     8,     8,    13,    10,    11,     6,     8,     8,     0,    -5,    -1,    -5,     1,    -1,    -2,    -3,    -7,    -2,    -8,     0,     1,     0,    -7,    -3,    -4,    -7,    -4,     6,    18,    11,     9,     4,     6,     6,     7,     2,    -1,    -2,    -2,     4,     2,    -1,    -2,    -2,   -12,   -10,    -7,    -1,    -1,    -1,    -2,    -4,    -8,   -11,    -8,     1,     5,     8,     6,     5,     4,     1,     1,    -1,    -4,    -3,    -3,     0,     3,     3,    -1,    -4,   -15,    -9,    -5,     0,     1,     0,     0,    -6,    -4,    -6,    -6,    -6,    -6,     0,    -1,    -1,     0,    -1,    -1,     2,     2,    -6,    -2,     6,     4,    -2,    -6,   -10,   -12,    -4,    -4,    -1,     0,     1,     1,     0,    -3,    -3,    -1,    -7,   -12,   -12,   -12,   -16,    -8,   -11,    -7,     0,     6,     8,     5,    -5,    -3,   -10,    -6,    -6,    -3,    -1,     1,     1,     1,     1,    -1,     1,    -1,    -4,    -5,    -9,    -6,    -5,    -5,     0,     4,     2,    -3,    -4,    -5,    -5,    -5,    -2,    -9,    -5,    -5,    -7,    -2,     0,     1,     0,    -1,    -1,     0,     0,    -2,    -3,    -1,     0,     0,     1,    -2,    -3,    -1,     1,    -2,    -2,     0,     1,     0,     0,    -3,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,    -1,     0,     1,    -1,    -1,     1,     0,    -1,     0,    -1,     1,    -1,     0,     0,     0,     0,     1,    -1,     0,    -1,    -2,     0,     1,     1,    -1,    -1,     1),
		    87 => (    1,     0,     1,     0,     1,    -1,    -1,     0,     1,    -1,     1,     0,     1,     0,     0,     0,     1,     1,    -1,     1,     0,     1,     0,     1,     1,    -1,     0,    -1,     1,     0,    -1,     1,     0,     0,    -1,    -1,     0,     0,     0,    -3,    -4,    -3,     0,    -5,   -10,    -9,     0,    -1,     0,     1,     0,    -1,     0,     1,    -1,     0,     0,    -1,     1,     0,    -2,     0,     1,    -1,    -1,    -2,    -6,   -11,    -2,    -1,     0,    -8,    -3,    -4,    -3,    -2,     0,    -1,     0,     0,     0,     1,     1,     1,     1,     0,     1,    -2,    -1,    -2,    -5,    -9,    -7,    -6,    -3,    -5,    -7,    -6,    -4,    -6,    -6,    -4,    -3,    -7,    -2,    -3,    -4,    -1,     0,    -1,     0,     1,     1,     1,     0,     1,    -7,    -4,    -3,   -12,   -12,   -10,   -21,    -8,    -4,    -1,    -2,    -3,    -9,    -7,    -7,    -7,    -8,     6,     0,    -7,    -8,    -4,    -2,    -1,     1,    -1,     1,   -10,    -4,     9,     1,     6,     3,     5,    -4,   -11,   -12,     0,    -5,    -8,    -4,    -8,   -10,    -5,    -4,    -3,    -5,   -11,    -5,    -7,    -1,     0,     1,    -1,     5,     7,     6,     9,     6,     6,     4,     5,    10,    -1,     1,    -6,    -6,    -7,    -3,    -1,    -5,     0,    -1,     0,     3,    -9,    -2,    -6,    -3,    -3,     0,     2,     7,     0,    11,    10,    12,    14,     2,    13,    12,     5,     5,     3,     2,    -2,    -4,     0,     2,     0,     1,     0,    11,     2,    -2,    -7,    -2,    -3,    -4,    -2,     0,     1,     1,     5,     2,     9,     2,     6,     6,     5,     8,     2,     3,     3,     0,    -1,    -2,     1,    -1,    -1,     8,     0,    -6,   -10,    -6,    -5,    -1,     0,     9,     4,     3,     1,     0,     3,     3,     0,     0,     2,     9,     5,     8,     4,     1,     0,    -1,     0,     2,     0,     5,     2,   -10,     1,     8,    15,    -1,    -4,     4,    -1,    -4,    -3,    -2,    -3,     2,     0,    -2,    -5,    -5,     1,    -1,    -1,     1,     5,     3,    -2,     3,    -4,    -3,    -3,    -4,     6,     8,    14,     1,    -3,     3,    -3,    -4,    -7,    -4,    -3,    -3,    -2,    -8,    -2,    -7,   -10,    -3,    -1,    -2,    -1,    -4,    -2,     1,    -6,     0,     2,    -8,   -10,    -7,     2,     0,     3,    -4,    -6,    -4,    -8,    -7,    -8,   -10,   -13,   -15,    -6,    -8,    -6,    -4,     2,     3,     0,     1,     2,     1,    -2,    -4,    -5,   -17,    -2,    -9,     2,     0,     0,     2,    -7,   -12,    -5,    -4,    -6,    -7,    -5,    -7,    -5,    -3,    -5,    -2,     6,    -2,     2,     3,     0,    -7,     4,    -3,    -1,    -9,    -5,    -7,    -4,    -1,     1,    -1,    -2,    -4,    -2,     0,     0,    -4,    -4,     2,     1,     3,     2,     3,     2,    -4,     7,     3,     6,    -1,     4,    -1,     3,     1,    -6,    -5,    -1,     1,    -1,    -1,     0,    -1,     0,     0,    -2,    -6,    -1,    -4,    -2,     0,     2,     1,     2,    -4,     4,     5,     0,    -6,     8,     0,     4,    -1,    -5,    -2,    -4,     1,    -2,     0,    -4,    -1,    -1,    -2,    -1,    -3,     0,     4,    -2,     3,     5,     0,    -1,    -1,    -1,     2,     1,     2,     1,    -2,    -4,     1,   -12,    -9,    -1,     0,     1,    -7,    -7,    -8,    -5,     4,     5,     1,     5,     6,     2,     3,     0,     0,    -2,     3,    -1,    -6,    -3,     2,     0,     1,    -1,     1,    -5,     2,    -5,     1,     1,    -1,    -4,    -5,    -1,    -4,     5,     1,     1,     1,     0,     0,    -1,    -3,    -4,    -5,    -2,    -6,    -3,    -1,    -6,    -2,    -2,    -3,    -6,     5,    -5,     0,     1,    -1,    -1,    -5,    -8,    -2,     1,     1,    -1,    -5,     1,    -1,     1,     1,    -2,    -6,    -4,   -10,    -6,    -7,   -11,    -4,    -1,     6,    -1,    -7,    -3,    -1,     5,    -2,    -4,   -13,   -11,    -6,     0,     1,    -1,    -4,     2,    -1,     0,    -2,    -4,    -3,   -11,   -13,    -8,    -8,    -8,   -11,     1,     1,    -8,    -7,    -1,    -1,    -1,    -3,    -9,    -5,    -6,    -7,   -11,    -8,    -7,    -3,    -3,     0,     1,    -3,    -3,    -4,    -8,   -10,    -7,    -9,    -6,    -9,     0,    -1,    -4,    -1,     1,    -2,    -1,    -2,   -11,     1,    -2,    -3,    -2,    -9,    -7,    -2,    -1,    -1,    -3,    -5,     0,    -2,     0,    -4,    -3,    -6,   -18,   -15,   -10,    -5,    -1,    -7,    -1,    -1,    -1,    -4,   -14,    -2,     0,     2,     3,    -9,    -4,     0,    -1,     1,     0,     0,     1,    -3,    -1,    -9,    -3,    -6,    -7,   -14,    -6,    -6,    -3,    -7,     1,     0,     0,     3,    -1,     4,     4,    -1,    -2,    -2,    -4,    -6,     0,    -1,     1,    -1,    -2,    -4,     5,    -6,    -2,     2,     3,    -7,    -6,    -5,    -2,    -1,     0,     1,     1,    -4,     3,    -3,    -4,    -4,     8,     4,    -3,    -6,    -4,    -2,    -1,    -1,    -5,     0,     0,    -2,     0,    -4,    -2,    -2,    -2,    -7,    -1,    -2,     1,     1,     1,    -1,    -5,   -16,   -12,   -14,    -4,     0,    -3,    -5,    -8,    -6,    -2,     1,     7,     0,    -3,     0,    -7,     1,    -1,    -3,    -5,    -1,     0,     0,     1,    -1,     1,     1,     0,     1,     1,     0,    -3,     2,     6,     8,     5,    -2,    -3,    -4,     5,     6,     8,     7,    -2,    -1,    -1,    -3,     0,    -1,    -1,     0,    -1),
		    88 => (    0,    -1,     0,    -1,    -1,     0,    -1,     1,    -1,     0,     1,     1,     1,     1,     1,     1,    -1,     0,     1,     0,    -1,     1,    -1,     0,     1,     1,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -3,    -5,   -13,   -14,   -11,    -2,    -2,    -2,    -2,    -2,    -1,     0,     1,    -1,    -1,     0,     1,     0,     0,     0,     0,    -2,    -1,    -5,    -5,    -7,    -8,    -5,    -3,     0,    -6,    -8,     3,     4,     0,    -5,    -8,    -8,    -1,    -2,    -2,    -1,     0,     0,     1,    -1,    -3,    -2,   -10,    -8,   -11,    -7,    -4,     2,     3,     4,     1,    -1,    -6,    -9,   -12,    -6,    -2,     2,     5,     1,     3,     3,    -3,    -1,     1,    -1,     1,     2,     0,    -5,   -11,    -8,    -8,     4,     2,     9,     9,     2,    -8,     0,    -4,    -4,     1,     0,    -5,    -4,     1,    -5,     2,     3,     3,     2,    -2,     0,    -1,    -4,    -3,   -10,    -9,    -9,     1,    -3,     3,     7,     5,     1,     4,     1,     5,     5,     7,     3,     0,     0,    -2,    -7,    -6,     4,     1,    -3,    -5,     1,     1,    -8,    -7,     2,    -7,    -9,    -5,    -1,    -1,     2,     1,    -2,     0,     3,     5,     5,     2,     3,    -4,    -2,     0,     3,     2,     1,     3,     0,    -1,     0,    -8,    -4,     2,     4,    -3,    -5,    -1,     2,     3,     1,     0,    -2,    -1,     0,     7,     7,     2,    -1,    -3,     3,     3,     6,     7,     3,     2,     1,    -5,    -4,    -5,    -4,    10,     5,     0,     3,     3,    -6,     1,     3,     0,    -1,     1,     1,     4,     3,     2,     2,    -2,    -2,    -3,     0,     4,    -2,     2,     4,     1,     1,    -4,    -6,     6,    11,     0,     1,    -3,    -2,     1,     1,    -4,    -2,    -3,     1,     3,    -1,    -4,    -1,     2,     0,     0,    -3,     1,    -1,     7,    10,    -8,    -1,    -4,    -8,    -5,     5,    -1,    -2,     0,    -4,    -6,    -5,    -6,    -3,     4,     5,    -2,    -9,    -7,    -5,    -4,    -1,    -4,     2,     2,     4,     3,     8,    -7,     1,    -2,    -6,    -3,     4,    -1,     4,    -2,    -3,    -2,    -8,    -4,    -1,     4,     0,   -11,   -10,    -6,    -4,    -1,    -2,    -2,    -2,     6,     2,    -5,     4,    -6,     0,    -1,    -1,     1,    -5,     0,    -7,    -9,    -5,    -6,    -2,     4,     4,     3,     3,     0,    -4,    -6,    -2,    -3,     1,     1,     3,     0,    -4,   -13,   -15,    -8,    -1,     0,     0,    -3,    -7,    -4,    -6,    -5,    -3,     7,     7,     6,     9,     4,     0,     2,     0,    -3,     1,    -2,     3,     6,     3,     1,    -9,   -12,   -11,     1,    -2,    -1,    -2,    -5,    -6,    -1,     2,    -3,     3,     8,     9,    10,     8,     5,     1,     3,    -1,    -2,     0,     4,     5,     5,    -2,    -5,    -5,     1,    -6,    -3,    -1,     0,    -3,    -1,    -7,    -1,     6,     6,     7,    11,    12,     6,     5,     7,     3,     1,     2,     0,     4,     4,     5,     2,     2,    -6,    -5,     9,   -10,    -3,    -1,     0,    -4,    -4,    -5,    -4,    -2,     5,     2,     8,    10,     9,     3,    -1,    -1,     0,     4,     9,     8,     2,     6,     4,     0,    -1,     0,     4,   -13,    -4,    -1,    -2,    -6,    -3,     1,    -6,    -7,     0,     1,     1,     3,     1,    -2,    -4,    -2,     5,     0,     2,     3,     3,     1,    -1,    -2,     2,     3,    -3,    -1,    -6,    -1,    -2,    -6,   -10,    -5,    -6,    -2,    -4,    -4,     0,    -2,    -5,    -5,    -1,     4,    -1,     0,    -5,     1,    -3,    -8,    -7,    -2,     4,    -2,    -8,    -1,    -2,     0,     1,    -3,   -11,    -6,   -10,    -8,    -9,    -8,    -7,    -4,    -5,     1,     5,     5,     2,     5,    -2,    -2,    -5,    -4,     0,     3,     1,    -4,    -9,    -5,    -4,    -1,     0,    -5,   -11,    -6,    -5,    -5,    -1,     0,    -6,    -3,    -3,     4,     5,     8,     6,     3,     1,    -4,     0,     2,     1,     1,     0,    -9,    -7,    -7,    -1,    -3,    -3,    -6,    -2,    -5,     0,     1,    -1,     0,     0,    -3,     6,    14,     6,     4,     8,     5,     4,    -1,     0,     2,    -5,    -3,     0,    -5,    -4,    -7,    -1,    -2,    -2,    -3,     0,     5,     3,    -1,    -3,    -4,     1,     1,     7,     4,     2,    10,     8,     3,    -1,    -1,    -4,     3,    -3,     2,     3,    -3,    -7,    -7,    -2,    -1,     0,    -2,    -1,     3,     1,    -3,    -6,    -3,     5,     6,     1,     4,    10,     7,     5,     3,    -4,    -1,     0,     4,     1,     3,     4,   -10,    -8,    -4,     0,     0,     1,    -3,    -3,    -2,    -4,    -5,    -6,    -4,     1,    -1,     2,     8,    11,     8,     1,    -2,    -4,     1,    10,     8,     2,    -7,    -4,   -12,    -6,    -3,     0,     0,     0,    -3,    -1,   -12,    -9,     0,    -4,    -8,    -8,    -1,     6,     5,     7,     3,     2,    -8,    -3,     1,     2,    -4,   -11,   -11,    -7,    -6,    -2,    -4,    -1,     1,     0,     1,    -5,    -4,    -5,    -8,    -6,     6,     4,    -5,    -2,    -1,     3,    -1,   -10,    -5,    -3,    -7,    -7,   -14,   -11,    -5,    -4,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -2,    -2,     0,    -7,    -9,    -5,    -1,    -2,    -6,   -11,    -8,    -8,    -7,    -4,    -2,    -1,     0,    -2,    -1,     1,     1,     0,    -1),
		    89 => (    0,    -1,     1,     1,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,     0,     1,    -1,     1,    -1,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,     1,     1,     1,     1,     1,     0,     0,    -1,     0,     1,     0,    -3,    -6,    -4,     0,    -1,    -2,    -1,    -4,    -4,     0,    -2,    -1,     0,     1,     0,     1,     1,     1,     1,    -1,    -5,    -2,     0,     0,    -2,    -2,     0,    -1,    -5,     0,    -1,    -7,    -3,    -2,    -2,    -3,    -3,    -4,    -2,    -2,     0,    -2,     0,     0,    -1,     0,     1,     1,    -3,    -5,    -6,    -5,    -6,    -2,    -2,    -1,    -4,    -3,    -5,    -7,    -6,    -5,    -5,    -8,    -5,    -3,    -3,    -3,    -1,    -1,    -1,     0,     1,     0,     1,    -1,    -1,    -3,    -1,    -7,     1,    -4,    -2,    -2,    -6,   -10,    -7,    -5,    -4,    -2,    -2,    -5,    -8,    -9,    -4,    -3,    -2,    -1,    -6,    -1,     1,    -1,     0,     1,    -3,     0,    -1,    -2,    -3,    -3,    -4,    -9,    -3,    -3,    -3,     0,    -1,     1,    -4,    -2,    -4,    -1,    -1,    -5,    -3,    -1,    -2,    -3,    -1,     0,     0,    -1,    -4,     0,    -1,    -5,    -5,   -12,    -5,    -4,    -5,    -2,     3,     8,     5,     3,     4,     0,     1,     3,     0,    -4,    -5,    -2,    -4,    -2,    -2,     0,     0,    -3,     0,    -3,    -7,    -9,    -8,   -12,    -1,    -2,     3,     3,     0,    -2,     4,     0,     0,    -3,    -1,    -1,    -1,    -4,    -4,    -7,    -3,     0,    -2,    -4,    -3,    -1,    -4,    -1,    -8,    -6,   -12,    -4,    -5,     3,     0,    -3,     0,     0,   -10,    -4,    -1,    -1,    -1,     1,    -4,    -3,    -6,   -10,    -3,    -2,     0,     1,    -1,    -2,    -3,    -8,    -9,    -6,    -9,     0,     2,    -1,     3,    -2,    -2,     2,    -5,    -5,    -2,     6,     2,     2,    -5,    -4,    -2,    -4,    -9,    -1,    -4,     1,    -2,    -4,     0,    -1,    -3,    -5,     2,     2,     1,    -6,    -4,    -9,    -7,    -4,    -5,    -9,    -6,     5,     1,    -1,    -7,    -3,     0,    -5,    -1,    -1,    -3,     0,    -8,    -1,     4,    -1,    -3,    -3,    -1,     2,    -2,    -4,   -11,    -6,    -1,    -3,    -4,    -5,     0,    -3,     0,     0,    -3,    -1,     4,    -6,    -2,    -1,    -4,    -1,    -1,     1,     3,     2,     2,     1,    -1,     4,    -3,    -4,    -9,    -2,    -6,    -9,    -6,    -3,    -3,    -7,    -1,     0,     3,     0,     1,   -11,    -4,    -1,    -2,    -1,    -5,    -4,     5,     5,     2,     1,     0,    -1,    -7,    -4,    -5,    -8,    -7,    -3,    -2,     2,    -6,    -7,    -1,    -1,     4,     0,    -4,    -8,    -5,    -2,    -1,    -1,    -4,    -6,    -1,     3,     2,     2,     1,     5,    -7,    -3,   -11,    -8,    -5,    -3,     2,     1,    -4,     3,     3,     0,     1,     2,    -8,    -5,    -3,     2,    -1,     0,    -1,    -5,    -2,     0,     0,     4,     3,     3,    -6,    -2,   -10,    -9,    -8,    -4,    -4,    -4,    -7,     3,     2,     5,     2,     1,   -13,    -9,    -2,     1,     0,     1,     0,    -6,    -4,     3,    -4,     6,     0,     1,    -3,     3,    -2,     0,    -2,    -5,    -6,    -7,    -4,     6,     2,     4,    -3,    -2,   -10,    -4,    -5,    -1,     0,     0,    -1,    -5,    -4,     4,    -4,     0,     5,    -5,     0,    -1,    -1,    -1,    -6,    -3,     0,     0,     0,     2,     2,     3,    -3,    -2,    -6,    -1,    -2,    -4,    -2,     0,     1,    -5,    -3,     4,     3,     3,    -1,    -3,    -1,     6,     2,     4,     1,     2,    -2,    -4,     3,     4,     1,    -2,     2,     3,    -4,    -9,     0,    -5,    -4,    -1,     0,    -3,    -2,     2,     8,     6,    10,    -3,     1,     6,    12,     3,    -1,    -4,    -1,    -1,     1,     5,    -4,    -1,    -3,    -1,    -5,    -3,     2,    -5,    -1,     1,    -1,    -2,    -2,    -1,     4,     2,    -1,     1,     2,    -1,     0,    -1,    -4,    -8,    -4,    -3,     2,     6,    -3,    -2,     1,    -1,    -2,     7,     3,    -5,     0,     1,     1,    -5,    -3,    -7,    -2,     1,     4,     3,     1,     0,    -1,    -4,    -3,    -3,     0,     1,     0,     3,     1,     2,    -5,     0,     1,     8,    -2,    -9,     1,    -1,     1,    -2,    -3,    -4,    -4,    -5,    -5,     0,    -1,    -3,    -5,    -2,    -6,     4,     1,    -2,    -1,     0,     1,     2,    -1,     3,    -2,     7,     2,    -7,     0,     0,     0,    -1,     1,    -4,    -5,    -4,    -6,    -6,   -11,   -11,   -10,    -8,    -2,     2,     5,    -4,    -2,    -5,     4,     1,     3,     8,    -1,     7,     2,    -5,     0,     0,     0,    -2,     1,    -1,    -1,    -2,    -2,    -4,    -5,   -10,    -9,    -2,     7,    -1,     0,     0,    -2,     1,     3,     5,     6,     8,     5,     6,     2,     0,     1,    -1,    -1,     4,    -3,    -3,     1,    -1,    -3,    -3,    -5,     0,     2,     5,     7,    -1,    -4,    -5,    -6,    -2,     8,    10,     6,    10,     5,     4,    -2,    -2,     1,     0,     1,     1,     1,     3,     0,     0,     1,     0,    -1,     0,    -1,    -2,    -5,    -3,    -9,   -11,    -6,    -1,     1,     7,     4,     3,     4,    -1,     0,     1,     1,     0,    -1,     0,     1,    -2,    -1,     0,     0,     0,     0,     1,     1,    -1,     0,    -3,    -1,    -4,    -7,    -5,    -5,    -3,    -4,     1,    -2,     1,     0,     0,     1),
		    90 => (   -1,     0,    -1,     1,     1,    -1,    -1,     0,     0,    -1,     1,     1,     0,     1,     0,    -1,    -1,     1,    -1,     1,     0,     0,     0,     0,    -1,     1,     0,    -1,    -1,     0,    -1,     1,     0,     1,    -1,    -1,    -1,     0,    -1,    -1,     1,     1,    -2,    -1,     0,     1,     0,     1,     0,     0,    -1,     0,     1,     0,     0,    -1,     1,    -1,     0,     1,     0,     0,    -3,    -1,    -2,    -3,    -3,    -2,    -2,    -3,    -2,    -1,     0,     1,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     1,    -2,     0,    -1,     0,     1,    -1,    -2,    -3,    -4,    -2,    -1,    -1,     1,     3,     3,     0,     0,     0,    -1,    -2,     1,     1,     0,     0,     1,     0,     1,    -2,    -2,    -5,    -3,     2,     1,     0,    -1,    -4,    -2,    -2,    -2,    -2,     3,     4,     2,     4,     4,     0,    -1,    -1,     0,    -1,    -1,     1,     1,     1,    -1,     1,     0,    -1,     1,    -4,    -2,    -2,    -2,    -1,     0,     1,    -2,    -2,     0,    -2,     0,     5,     5,     1,    -1,    -1,    -1,    -1,    -1,    -4,     1,     0,    -2,    -2,    -1,    -3,     1,     2,     1,    -2,    -2,    -1,    -2,    -3,    -1,    -2,     3,     1,     0,     2,     3,     2,    -2,    -2,    -2,    -5,    -1,     0,     0,    -2,    -2,    -3,    -1,     1,     4,     1,    -2,     2,     2,     1,     2,     1,     0,     5,     1,     3,     6,     2,     0,     1,     4,     0,    -1,     0,    -3,     0,     0,    -1,     3,    -2,     2,     2,     2,     3,     2,    -3,    -2,     1,     3,    -2,    -1,    -2,     0,     2,     1,     2,     4,     4,     2,     2,    -2,    -1,    -3,    -2,    -1,     0,     1,    -1,     6,     1,    -2,     0,     2,     2,    -2,    -6,    -7,    -5,    -5,    -5,    -2,    -1,     0,     0,     0,     5,     3,    -1,     1,    -2,     0,    -1,     1,     1,     1,     0,     0,     5,     4,     4,     3,     1,    -6,    -5,    -6,    -4,    -3,     0,    -5,    -4,    -4,    -2,    -2,    -3,     4,     1,    -1,    -2,    -3,     0,     1,     4,     1,    -1,     3,     5,     2,    -3,     1,    -5,    -6,    -8,    -6,     0,     1,     2,    -3,    -3,    -5,    -8,    -7,    -4,     0,     1,     4,     0,     0,    -1,    -1,     0,     1,    -1,     3,     2,     1,    -2,    -1,    -4,    -7,    -8,    -5,     0,    -1,    -2,    -8,    -9,    -5,    -6,    -6,    -2,     0,    -1,     2,     2,    -1,     1,     1,    -1,     0,     1,     6,     1,     5,    -3,    -3,    -6,    -9,    -9,    -5,    -3,    -1,    -3,    -7,    -6,    -7,    -6,    -6,    -3,     0,     3,     3,     1,     0,    -2,     1,     0,     0,    -4,     7,     4,    -1,    -5,    -7,    -8,    -7,    -6,    -6,    -5,    -3,    -7,    -6,    -5,    -5,    -6,    -6,    -3,    -4,    -1,    -3,     2,    -2,    -1,    -1,     1,     0,     1,     6,     3,    -1,    -3,    -5,    -7,    -5,    -6,    -3,    -3,    -3,    -1,    -3,    -5,    -4,    -5,    -6,    -3,     1,     0,    -2,     1,    -2,     0,     1,     0,    -2,     0,     3,     4,     3,    -1,    -2,    -3,    -4,    -3,    -4,    -3,     3,    -3,    -3,    -8,    -7,    -7,    -3,    -5,    -1,     5,     0,     2,    -3,     1,     1,    -1,    -2,     3,     5,     4,     4,     4,    -3,    -3,     1,     0,    -3,    -3,    -2,    -4,    -8,    -7,    -7,    -7,    -4,     0,     3,    -1,    -1,     2,    -7,     1,     1,     0,    -1,    -1,     7,     2,     2,     4,    -1,    -1,     0,    -3,    -1,    -2,    -6,    -3,    -6,    -6,    -9,    -5,    -3,     2,     0,     1,     0,    -1,    -1,    -1,     1,     0,     1,     0,     5,     0,     1,     2,    -1,     0,     1,    -1,     0,    -2,    -2,    -3,    -5,    -2,    -2,    -1,     3,     0,     0,    -2,     1,    -4,    -2,     0,    -1,     0,     1,     0,     4,    -2,     4,     2,     1,    -3,    -2,     1,    -2,     0,     1,     0,     3,     3,    -4,    -1,     1,    -1,     2,    -2,     0,    -3,    -1,     0,     1,     0,    -2,     0,     0,    -4,     0,     5,     0,     0,    -1,     2,    -2,     0,    -1,     0,    -2,     1,     0,     2,     2,     1,    -3,     0,    -2,     0,     1,     1,     1,    -1,    -1,    -2,    -3,    -2,    -4,     4,     1,    -1,     1,     2,    -2,     1,    -1,    -3,     2,     3,     0,     1,     1,    -2,    -1,    -2,    -3,     0,     1,     1,     1,     0,     0,    -2,    -2,    -2,     2,     3,    -1,    -2,    -1,     0,     1,    -3,    -1,    -1,    -3,    -1,    -2,     1,     0,     0,     0,    -3,    -4,    -3,    -3,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     4,     3,     2,    -3,     0,    -1,    -2,     1,     3,     2,     1,     1,     2,    -2,    -2,     0,    -1,    -1,     0,     0,    -1,     1,    -1,     0,     1,     0,    -1,    -1,     3,     5,     5,     1,     0,     0,    -2,    -2,    -3,     0,     0,    -2,    -6,    -7,    -6,    -4,    -4,    -3,    -1,    -1,     0,     0,     1,     1,     1,     0,     0,    -3,    -4,     0,    -1,     0,    -1,     0,     0,    -3,    -3,    -2,    -3,   -10,    -5,    -5,    -5,    -4,    -2,    -4,     0,    -1,     1,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,    -2,    -1,     0,     0,     0,     0,    -1,     1,    -3,    -3,    -3,     0,     0,     0,    -1),
		    91 => (   -1,     0,     1,     0,     1,    -1,    -1,     0,     1,     0,     0,     0,     1,    -1,     0,     1,     1,     1,     1,     0,    -1,     0,     1,     1,     1,     1,     1,    -1,     0,     0,     0,     1,     0,     1,     0,     0,     1,     0,     0,    -1,     0,    -2,     6,     3,     4,    -4,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     1,    -1,     1,    -1,     1,     1,    -1,     0,     1,    -4,    -4,    -3,    -4,    -1,     2,     2,     5,    10,     6,     6,     2,     3,    -7,    -5,    -6,    -1,     0,    -1,     0,     0,    -1,     8,     4,    -1,    -4,    -7,     4,     1,     1,    -5,    -9,    -4,     0,    -1,     1,     2,     0,     1,    -6,    -2,    -4,    -3,    -4,    -3,    -1,     0,    -1,     1,     0,     8,     7,     6,     0,    -2,     3,     5,     4,     3,     1,    -6,     1,    -2,     2,    -1,     0,     0,    -6,    -6,    -3,     6,     5,     4,    -3,    -2,    -3,     0,    -1,     3,     2,     9,     7,     1,     1,     5,     1,    -1,    -1,    -2,    -3,    -6,    -1,    -2,    -2,    -3,    -2,    -7,     2,     6,     8,     6,    -5,    -3,    -4,    -1,    -1,    -4,     0,     9,     3,     3,    -1,    -5,    -4,    -1,    -2,     2,    -3,    -2,    -4,    -5,    -4,    -3,   -10,    -3,     4,     7,     6,     2,     0,    -2,    -2,     1,     0,    -4,    -5,    -4,    -4,    -5,     3,   -10,    -2,     9,     7,     5,    -1,     2,    -3,    -8,    -4,    -2,    -7,    -2,     5,     6,     7,     1,    -3,    -5,    -2,    -1,     0,    -6,    -4,    -4,    -5,    -4,     6,    -8,    -2,     8,    -1,     5,     0,    -2,    -3,    -4,    -6,    -6,    -6,     3,     3,     3,     1,     1,    -3,    -5,    -2,     0,     0,    -5,     0,    -4,    -5,    -3,     7,    -3,     1,     3,     0,    -4,    -5,    -4,    -3,    -5,   -10,    -6,    -8,     1,     1,     3,     3,     1,    -1,    -5,    -2,    -1,    -1,    -3,     0,    -3,    -2,    -5,     3,     2,    -3,     5,     1,     1,     0,    -1,    -3,    -8,    -7,    -2,    -2,     0,     0,     3,     5,    -3,    -1,     1,     2,    -1,     1,     0,     0,     0,    -4,    -7,     3,    -5,    -2,    -1,    -3,    -1,    -3,     3,     0,    -7,    -2,    -2,    -2,    -2,    -3,     4,     2,    -3,     1,     0,     6,    -1,     1,    -4,     0,     1,    -2,    -3,    -3,    -6,    -5,     0,     0,    -2,    -4,     2,    -2,    -2,    -2,    -1,    -2,    -2,    -4,     0,     1,    -5,     2,     4,     7,     1,    -1,    -3,     0,    -1,    -3,    -1,    -1,     0,    -2,    -2,    -3,     1,    -3,     0,     1,    -3,    -2,    -6,    -2,    -4,    -5,    -4,   -10,    -5,     4,     1,     1,     0,     1,     1,     2,    -2,    -4,     1,    -2,    -3,    -4,    -9,   -12,    -4,     4,     3,     3,     0,    -1,    -2,    -8,    -6,    -7,    -8,    -4,    -3,    -5,     0,     0,     1,     0,    -1,     0,    -3,    -9,    -4,    -4,    -6,    -9,   -13,   -11,    -4,     2,     5,    -4,    -5,     2,     1,    -6,    -7,    -4,    -7,    -4,    -9,    -8,    -7,    -2,     1,    -1,     0,     0,    -3,    -2,    -4,    -4,    -6,    -1,    -5,    -4,    -6,    -2,     6,     1,    -3,     2,     1,    -2,    -2,    -1,     0,    -3,     6,    -8,    -6,    -2,     1,     0,    -1,    -2,    -1,    -1,    -2,    -3,     1,     0,     3,     1,    -4,    -2,     4,    -1,     3,    -3,     2,     1,     4,     3,     3,    -1,     0,    -6,    -4,    -4,     1,    -1,    -1,    -4,    -3,     0,    -5,     0,     3,     6,     4,    -6,    -7,    -5,     2,     1,     1,     4,     1,     2,    -4,    -2,     2,     0,     1,     0,    -4,     0,    -1,     0,     3,    -4,    -3,    -1,     7,     8,    10,     9,     7,     1,    -7,     0,    -1,     3,     5,     1,     2,    -3,     0,     0,     5,    11,     4,     3,    -4,    -2,     1,     0,     0,    -2,     3,     5,     7,     8,     6,     5,     4,     0,    -3,    -1,     3,     0,     3,     0,     1,     1,     7,     6,     8,     4,     2,     0,    -3,    -1,     2,     2,    -1,    -1,    -3,    -5,    -3,     0,    -1,    -3,    -3,    -6,    -2,     1,    -4,     0,    -5,    -3,     1,     3,     3,    -1,     4,     1,     0,     4,    -2,     0,     4,     2,    -3,    -2,    -2,     4,    -1,    -3,    -7,    -6,    -5,    -7,     1,     1,     0,     2,    -5,    -2,    -1,    -1,     1,     0,    -6,    -4,    -1,     0,     1,    -1,    -1,    -1,    -1,    -3,     1,     5,     6,     3,    -1,    -1,     1,     0,     5,     1,    -4,    -4,    -4,     3,    -2,    -2,     5,     1,    -3,    -4,    -3,    -4,     6,     0,     1,     0,     1,    -2,     0,     0,     0,    -2,    -2,    -2,     1,     1,    -1,     0,    -4,    -9,    -4,    -5,    -3,    -7,    -1,    -7,    -3,    -3,    -6,     4,     5,     1,    -1,     0,     0,    -2,    -2,    -3,    -1,    -3,    -4,    -2,    -4,    -1,     0,     4,     5,    -3,    -7,    -5,    -5,    -5,    -9,    -6,    -3,    -2,     1,     0,    -1,     0,    -1,     0,     0,    -2,    -2,    -6,    -5,    -4,    -2,    -2,    -1,     0,    -2,    -4,    -5,    -4,    -3,    -5,    -1,    -1,    -2,    -2,    -1,    -1,     1,     1,     1,     1,     0,    -1,     0,     1,    -1,     0,    -1,     0,    -1,     1,    -2,    -4,     1,    -1,    -1,     0,    -1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0),
		    92 => (    1,     1,     1,     1,     0,     0,    -1,    -1,     0,    -1,     1,    -1,    -1,    -1,     2,     2,     1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     1,     0,     1,     0,     1,    -1,     1,    -2,    -4,    -6,    -8,    -2,    -2,    -1,     3,     4,     0,    -3,   -10,    -6,    -7,    -5,    -1,     1,    -1,     0,     1,     1,    -1,    -1,    -3,    -3,     0,     1,     1,     1,     8,     8,     9,     1,     3,     7,    11,     9,     4,    -4,    -9,    -5,    -2,    -5,    -1,     0,     0,     1,     1,    -1,     0,     0,    -6,    -8,     4,     5,     7,     0,    -6,    -8,   -11,   -14,     0,    -2,     0,     1,    -4,   -11,    -7,    -6,    -1,     0,    -7,    -7,    -1,    -1,     0,    -1,     0,    -2,    -5,     0,     3,    12,     9,     7,    11,     3,    -3,    -4,    -4,    -3,     2,    -3,    -1,     2,    -2,    -2,    -5,     1,    -5,    -9,    -1,    -6,    -2,     0,    -1,    -5,    -3,     0,    -5,    -4,     1,     7,     2,     5,     0,     2,     2,     3,     1,     0,     1,     3,     4,     2,     6,    -2,    -4,    -8,     3,   -11,    -3,     0,    -1,     1,     0,     3,    -1,    -1,    -2,     5,    -1,     1,    -5,     1,    -4,     0,     0,     3,     2,     5,     2,    -1,     2,    -1,    -3,   -13,    -2,   -10,    -2,    -1,    -1,     4,     0,     5,    11,     3,     1,     3,    -1,    -7,    -4,     0,     2,    -2,     2,     4,    -3,     1,    -2,     1,     6,     5,    -9,     2,     6,    -6,    -4,    -6,     7,     4,     1,    -1,     9,     3,    -2,     3,     2,    -2,     2,     2,     0,    -1,    -5,    -3,    -1,    -4,     1,     0,    -4,     0,     6,    -2,    -4,   -10,    -3,     1,    -4,     1,     5,    -6,     1,     0,    -3,     0,    -3,     0,     3,     4,     3,    -2,     0,    -2,    -1,     0,    -2,     0,    -2,     5,    -1,    -5,   -14,    -2,    -2,     1,     1,    -3,     3,    -3,     6,    10,     1,     1,    -3,     6,    -2,     0,     0,    -2,     0,    -3,     7,    -4,    -4,    -1,     1,    -3,    -9,    -5,    -4,    -3,    -4,     0,    -5,     1,     1,    -2,     3,     5,     4,     1,     3,     4,    -1,    -5,    -6,    -1,    -5,    -1,    -4,     0,     2,     2,    -1,    -7,    -5,     2,     3,    -3,    -6,     0,    -3,    -9,     0,    -3,     1,     9,     4,     0,     6,    -1,    -6,    -4,    -3,    -7,    -5,    -5,    -3,     4,     7,    -3,     6,     5,    -5,     6,     2,     0,    -2,    -1,    -5,    -3,    -1,    -1,     4,    15,     5,    -2,     1,    -2,    -1,    -2,     2,    -6,    -4,    -5,    -2,     3,     5,    -1,     1,     5,    11,     8,     9,     9,    -1,     1,    -1,    -2,     1,     4,     5,     9,    10,    -5,     3,     1,    -8,    -4,    -5,    -4,    -3,    -2,     0,    -1,     4,    -7,     3,     9,    16,    14,     7,     6,     3,     0,    -4,     7,     8,     0,     2,     4,     4,     6,     1,    -3,    -2,    -2,    -4,    -1,     0,    -2,    -4,    -1,    -3,     2,     5,     5,     5,    -1,     5,    11,     9,     0,     0,     9,     8,    -5,    -4,     1,     9,     4,     9,     4,     1,     4,    -1,    -2,    -2,    -1,    -4,    -3,     2,    -2,    18,    14,     9,     2,    10,    12,     7,     0,    -2,     9,     6,    -2,    -3,     2,    -1,    -2,    -1,     1,     0,     1,     0,     3,    -2,    -3,     0,    -1,    -1,     5,    18,    10,     4,     3,     5,     5,     4,    -1,     0,     1,     3,    -2,    -1,     1,    -4,     2,    -2,    -3,     1,     2,    -1,    -6,    -3,    -4,    -6,    -1,     4,    16,    14,    11,     8,     6,     5,    -2,     2,     1,    -5,     2,    -2,     0,     0,    -3,     0,     3,     2,     3,     4,    -2,    -3,     1,     4,    -3,    -7,     3,     9,    10,    13,     9,     4,     0,    -3,     2,     7,    -1,    -3,     8,    -4,    -2,     0,     0,     0,     0,     4,     6,     6,     0,     0,    -5,     1,    -5,    -2,     3,    11,    13,    16,     7,     5,     2,     1,     1,    -1,    -1,    -1,     8,    -3,     5,    -1,     2,     0,     6,     9,     5,     0,     3,     3,    -5,     0,    -1,    -5,    12,    18,    14,    12,    15,     2,    -2,     1,    -2,    -1,     0,     0,    -3,    -6,    -2,     2,    -4,     0,     5,     5,     2,     3,    -3,     0,    -3,    -2,     1,     4,    16,    15,    14,    11,    10,     4,    -6,     2,    -1,    -1,    -1,     1,     0,    -8,     0,     2,     4,     1,     2,     9,     4,     2,     2,     1,    -3,    -3,    10,    19,    15,    11,    15,    14,    10,     6,    -5,     0,     0,    -1,     1,     0,    -6,    -2,    -5,    -9,     4,    -3,     0,     4,     5,     2,    -8,   -12,    -2,     1,    12,    16,    21,    15,     9,    12,     9,    -2,     3,     1,     3,     0,     1,     0,    -2,    -1,    -7,   -14,     5,    -4,    -4,    -5,    -8,    -7,   -10,    -9,     1,     2,     2,     8,    13,     4,     1,     2,    -5,    -5,    -3,     0,     2,    -1,     1,     1,     1,    -1,    -2,    -4,    -9,   -13,    -6,   -14,   -17,   -13,   -11,   -17,   -17,   -13,   -13,   -12,   -10,   -16,    -5,    -3,    -6,     1,     0,     0,     0,     0,     1,     1,    -1,     1,    -2,    -2,    -2,    -2,    -1,    -2,    -6,    -7,    -5,    -7,    -7,    -3,    -4,    -3,    -2,    -3,    -2,    -2,    -3,     0,    -1,     1,     1,     1),
		    93 => (    0,     0,    -1,     1,    -1,    -1,     1,     0,     1,    -1,     1,     0,    -1,    -2,     0,    -1,     1,    -1,    -1,     1,     1,     1,     0,    -1,     1,    -1,     0,     1,     1,    -1,     0,     0,     1,     0,     0,    -1,     1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -1,     0,    -1,     0,     0,    -1,     1,     1,    -1,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -5,    -6,     7,     2,    -2,    -5,    -8,    -5,    -5,    -3,    -4,    -3,    -9,    -7,    -8,    -5,    -1,     0,     1,    -1,     0,     0,    -1,    -1,     0,    -2,     1,     3,    -5,    -7,   -10,    -8,    -9,   -12,   -15,    -8,    -6,    -7,   -10,    -7,    -6,    -4,    -3,    -6,    -2,    -2,     0,     0,    -1,     0,     1,     0,     2,     7,     8,    -3,    -2,   -10,    -2,    -2,    -3,    -7,   -12,   -11,   -11,   -10,   -10,   -10,    -8,    -2,    -4,    -3,    -2,    -5,     0,     1,     1,    -1,     0,     2,     3,     7,     1,    -3,    -1,     3,     6,     5,     5,    -2,    -4,    -2,    -4,    -3,    -7,   -10,    -7,    -6,    -6,    -3,    -1,    -6,    -2,     1,     0,     0,     0,     4,     2,    -4,     2,     5,     0,     4,    -2,     3,     1,    -3,    -5,    -5,    -7,    -6,    -5,    -9,    -7,    -6,    -6,    -6,    -4,    -1,    -4,     0,     0,     2,    -1,     4,     1,    -1,     5,     2,     4,    -1,    -1,    -6,     0,     1,    -2,     3,    -5,    -8,   -11,   -12,    -7,    -7,    -5,    -6,    -4,    -1,    -3,    -1,     1,     1,    -4,     2,     0,     0,    -2,    -5,    -1,    -1,    -6,     0,     7,     7,     8,     5,    -1,   -10,   -12,   -13,   -10,    -4,    -5,    -6,    -4,    -2,    -2,     1,    -1,    -3,    -3,     1,    -2,     2,    -4,    -3,    -5,    -2,    -3,     5,     6,     7,     8,     1,    -5,   -14,   -13,   -13,    -9,    -5,    -4,    -2,    -3,    -4,    -3,    -1,     0,    -6,    -2,     7,     1,     4,     0,    -3,    -5,     0,     1,     3,     5,     4,     1,    -5,    -7,   -15,   -16,   -13,   -10,    -9,    -5,     0,    -2,    -3,    -2,     0,    -1,    -8,     0,     9,     5,     1,    -1,     0,    -2,     2,     4,     2,     4,     0,    -4,    -5,    -5,    -7,    -6,    -8,    -6,    -9,    -7,    -2,    -1,    -6,    -4,     0,     0,    -6,    -7,     6,    -2,     0,    -6,    -4,     3,     2,     6,     5,     5,     1,     1,     1,    -5,    -5,     2,     0,     0,     3,     7,     5,    -5,    -4,    -2,    -1,     0,    -2,    -6,     7,     4,     1,    -1,    -3,     3,     5,     5,     4,     4,     3,     1,    -3,    -1,    -1,     2,    -1,    -2,     2,     4,     6,     6,    -5,    -3,     0,    -1,     2,    -1,     3,    -6,    -4,    -4,    -3,     1,     4,     2,    -1,    -1,     0,    -3,    -1,     2,    -3,    -1,     5,    -1,     1,     1,    11,     4,    -6,    -2,    -1,     0,     3,     0,     2,    -6,    -5,    -4,    -1,     3,     1,    -2,    -5,    -4,    -4,    -1,    -4,     1,     0,     0,     4,     7,     5,     4,     4,     1,    -5,    -1,     0,     1,     1,     0,     0,    -6,   -10,    -4,    -7,     1,     5,    -4,    -5,    -5,    -9,   -11,    -3,    -5,    -4,     0,     2,     6,     6,     6,     0,    -1,    -4,    -4,    -2,     1,     0,    -1,     5,    -2,    -5,    -4,    -8,    -3,    -4,    -9,    -5,    -5,    -5,   -10,   -10,    -5,    -5,    -8,     3,     3,     9,     4,     3,    -1,    -4,    -2,    -1,    -1,    -1,     1,     0,     0,    -3,    -6,    -4,     0,    -3,   -10,    -4,    -2,    -5,    -4,    -8,    -4,     0,    -2,     0,     3,     4,     3,     0,     2,    -3,    -2,    -4,     1,     0,    -2,    -3,    -3,    -2,    -3,     2,    -1,    -2,    -5,    -3,     1,     3,     1,    -2,     1,     4,    -2,     0,     1,     2,     1,    -3,     2,    -1,    -5,    -3,     1,     0,    -3,    -5,    -4,    -5,    -6,     0,     2,     3,    -2,     1,     2,     3,     4,     5,     6,     0,    -3,    -2,     4,     4,     1,    -1,     3,    -2,    -2,    -1,    -1,     0,     0,     0,     3,    -1,    -8,    -6,    -3,    -2,    -4,    -3,    -5,    -2,     1,     0,     1,    -2,    -4,     0,     0,    -5,    -2,     2,    -3,     0,    -3,    -1,     0,     0,     0,     0,     0,    -1,    -7,    -7,    -7,    -6,    -4,    -5,     0,     0,    -5,    -2,    -5,    -5,    -2,    -2,    -2,    -2,    -1,     2,    -3,    -3,     0,     1,     1,     1,     2,    -4,    -1,    -2,    -1,     0,    -3,    -3,    -4,     0,     2,    -2,    -4,    -2,    -4,    -3,    -6,    -3,    -3,    -3,    -3,    -5,    -1,    -2,     0,     0,     1,     0,     3,    -2,    -4,    -3,     3,     4,     2,     0,     0,     9,     2,    -3,    -1,    -2,    -5,    -6,    -4,    -1,    -4,     0,    -1,    -7,    -3,    -2,     0,     0,     1,     0,     1,    -5,     0,    -2,     1,     2,     1,     0,    -2,    -2,    -2,     3,     2,    -2,    -4,    -3,     0,    -1,    -9,    -6,    -5,    -8,     0,     0,     1,     1,     0,     1,     0,    -2,    -2,    -3,    -3,    -3,    -6,    -6,    -2,    -5,    -4,     0,    -7,    -3,     1,     0,    -4,    -3,    -3,    -1,    -6,    -1,     1,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -3,    -2,    -3,    -3,    -4,    -3,    -6,    -1,     1,     0,    -5,    -2,    -3,    -2,     1,     0,     0,     1,     0),
		    94 => (    0,    -1,     0,    -1,     0,     1,     0,     0,     1,     1,     1,    -1,    -2,    -1,    -2,    -2,     0,    -1,    -1,    -1,     1,     1,     0,     1,    -1,     0,     0,    -1,     1,     1,     0,     1,     0,     0,    -2,    -5,    -1,    -4,    -5,    -5,    -5,    -4,    -1,    -6,    -6,    -3,     0,     0,    -5,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -6,   -10,    -2,    -5,    -7,    -4,    -5,    -9,   -14,    -9,    -6,    -9,    -4,    -1,    -3,    -6,    -6,    -6,    -1,    -5,    -4,    -6,    -3,    -1,     0,     0,    -1,     0,    -7,   -12,    -3,    -9,    -9,    -5,    -7,    -8,    -4,    -5,   -10,    -7,    -5,     4,    -5,    -7,     0,    -1,     1,     1,     2,    -7,    -4,     1,     1,     1,     1,    -3,    -6,     1,    -4,    -7,     1,     1,    -2,    -7,    -1,     3,    -4,    -4,   -10,    -3,    -6,    -5,     6,     4,     3,     0,    -4,    -7,     1,    -2,     0,     0,     0,    -3,    -7,    -7,    -4,    -5,    -1,     2,     2,     7,    -2,    -2,    -4,    -7,   -10,    -4,     2,    12,     2,     1,     2,    -4,    -4,    -7,     3,    -4,     1,     0,     0,    -1,    -1,    -4,    -4,    -1,     1,    -2,    -1,    -8,    -4,    -4,    -1,   -11,   -18,    -3,     1,     5,     7,    10,    10,    -5,    -3,    -5,    -4,    -1,    -4,     1,    -3,    -5,     0,    -4,    -1,    -2,     6,    -2,    -5,    -7,     1,     5,    -3,   -14,   -12,    -2,     3,     5,     4,     3,     3,    -3,    -4,    -7,    -6,    -2,    -4,    -5,    -6,     5,     0,    -3,     0,     2,     3,    -4,    -6,    -5,     3,     0,    -5,    -8,    -6,    -6,    10,     1,     4,     0,    -6,    -6,    -8,    -7,    -3,    -6,    -3,     0,    -5,     3,    -2,    -3,    -4,     1,    -1,    -3,    -2,    -8,    -1,    -2,    -2,    -5,    -9,    -1,     6,     3,    -2,     0,     5,     1,    -6,    -6,    -2,    -2,    -3,     0,    -4,     4,     6,    -1,    -4,    -6,     1,     1,    -4,     3,     0,    -2,    -1,    -6,   -12,    -3,     4,     1,    -2,    -3,     4,    -5,   -10,    -9,    -2,     0,    -2,     1,    -8,    -2,     5,    -5,     0,    -2,    -2,     3,     0,     2,     4,     2,    -3,   -12,    -9,     1,     5,     0,    -1,    -4,    -9,    -8,    -8,   -13,    -5,    -1,    -6,     1,    -4,     2,    -1,    -5,     0,     6,     2,     0,    -1,     6,     2,     3,    -9,    -9,    -9,     0,     1,     1,    -2,    -5,    -7,    -8,     1,     3,     2,    -4,    -5,     0,    -4,    -1,    -1,    -2,     0,     6,     1,     0,     2,     4,     4,    -2,    -8,   -10,    -8,    -3,     2,     3,    -4,    -6,     1,     5,     4,    -4,    -3,    -6,     1,     1,     0,    -7,    -2,     8,     5,     0,     3,    -2,     6,     8,     6,    -1,    -2,    -3,    -6,     0,     1,     2,     2,     2,     5,    -1,     1,    -2,    -6,    -5,     0,     0,    -1,    11,     0,     6,     2,    -2,    -2,     1,     1,     5,     4,     4,     1,    -4,    -6,    -2,    -1,    -1,     4,    -1,     3,     9,    -3,    -8,    -9,    -4,     1,     0,    -1,     0,    -6,    -3,    -6,     2,     0,    -3,    -1,    -1,    -9,    -5,    -3,    -5,    -2,    -1,     1,     2,    -2,     5,     2,    -1,   -10,    -2,    -5,    -6,    -3,    -1,     1,     3,    -9,     0,    -1,     0,     3,     4,    -1,     0,    -1,    -9,    -1,     0,     3,    -1,     2,     3,    -3,     1,     4,    -5,    -3,    -6,     4,    -1,    -4,    -3,     1,     3,    -5,     2,     4,     3,     5,     0,    -1,    -3,    -3,    -9,    -2,     2,     6,    -1,     2,     1,     2,     5,     1,    -7,    -2,    -6,    -5,    -2,    -1,     1,    -1,    -5,     0,    -2,     1,     6,     0,     1,     1,    -1,   -10,   -10,    -3,    -2,     6,     1,    -4,     5,     3,     3,     5,    -5,    -3,    -6,    -8,     0,    -1,     0,     1,    -3,    -1,     1,    -3,     0,     2,     0,    -4,    -7,    -2,    -1,     0,     0,     1,     0,     3,     4,     4,     4,     5,    -5,    -2,     0,    -3,     0,     0,    -1,     1,    -6,    -1,     1,    -2,     1,     2,     2,    -6,    -5,    -6,    -1,     0,     0,     2,    -3,     4,     3,     1,     4,     5,     4,    -3,     4,    -1,    -4,    -1,     1,     1,     0,    -6,    -9,     4,     1,    -1,    -6,    -9,   -14,    -7,    -5,     0,    -1,    -2,    -3,    -4,     2,     4,     5,     6,     2,    -2,    -1,     8,     2,    -1,     0,     0,    -1,    -4,    -7,    -5,    -1,    -3,    -1,   -10,   -12,    -7,    -6,    -4,    -1,     0,     3,    -5,     0,     3,     6,     9,    -5,    -4,     1,     2,     2,    -1,     1,     1,    -1,    -1,    -3,    -1,     0,    -1,    -4,    -6,    -7,    -7,    -4,    -1,    -6,    -3,     1,    -2,     0,    -2,     1,    -1,    -7,    -1,    -6,    -4,    -3,     0,    -1,     1,    -3,    -1,    -4,     0,    -1,     0,    -3,    -6,    -9,    -3,     0,    -4,   -11,     0,     2,    -2,    -6,   -11,    -6,    -8,   -10,    -5,    -7,    -5,    -3,     1,     0,    -1,     0,    -1,    -5,     0,    -1,    -1,    -2,    -6,   -11,    -1,    -3,    -7,   -11,    -7,   -12,    -9,    -9,    -8,   -12,    -9,   -10,    -1,    -1,     1,    -1,     1,     1,    -1,     1,     1,    -1,     1,    -1,    -3,    -2,    -4,    -6,    -5,    -5,    -3,    -5,     1,    -7,    -9,    -6,    -5,    -5,    -3,    -6,    -2,     1,     0,     1,    -1),
		    95 => (    0,     1,     1,     0,    -1,     1,     1,     0,     1,     1,     0,    -1,     1,    -1,     0,     0,     0,    -1,     0,     1,    -1,    -1,    -1,     0,    -1,     1,     0,    -1,     1,     0,    -1,     0,    -1,     1,     0,     1,     0,     1,    -1,    -1,     0,     0,    -1,    -2,    -2,    -3,    -1,    -1,     0,    -1,     1,     1,     0,    -1,     0,     1,     0,     0,    -1,     1,     1,    -1,    -2,    -3,    -3,    -5,    -4,    -4,    -5,    -3,    -2,     3,    -1,    -1,    -1,     2,     4,     2,     2,     5,    -1,    -1,     0,    -1,     0,     0,    -2,     1,     0,    -1,    -5,    -7,    -2,     0,     5,     1,     5,     7,     9,     3,    -2,    -5,     7,    -2,    -2,     2,    -3,    -3,    -4,     1,     2,    -1,     1,    -1,    -3,     0,    -4,    -4,     4,     0,    -7,     5,     0,     4,     5,    -5,    -5,    -2,     2,    -3,     2,     6,    -4,     1,     5,     6,    11,    10,     3,    -3,     1,     1,    -2,     1,     0,     1,    -3,    -6,     1,     8,     7,     0,    -6,    -6,    -4,    -2,     3,     0,     2,     1,     2,     5,     5,     5,     8,     6,     6,    -2,     0,    -1,    -1,    -2,     3,     2,    -4,    -2,     7,     1,     2,    -6,    -6,    -1,     2,     7,     3,     6,     4,    -2,     2,     4,     7,    -1,     4,     4,     6,     0,     0,     0,     0,    -4,     0,    -1,    -3,     4,     4,     5,     5,    -1,    -6,    -3,     7,     6,     9,     7,     2,     2,     2,     2,    -2,    -4,    -3,     5,     5,     2,     0,    -1,    -7,    -5,    -6,    -3,     0,     2,     8,     6,     6,    -4,    -3,    -6,    -1,     2,    -2,     1,     2,    -4,    -1,    -6,    -4,    -4,    -3,    -5,     7,     1,    -1,    -2,    -7,    -7,    -4,    -2,     1,     1,     4,     5,     3,     4,    -9,   -11,   -13,   -16,   -17,   -22,   -12,   -16,   -16,   -15,   -10,    -7,    -7,    -5,     7,     4,     1,    -1,    -2,    -5,    -2,    -1,    -3,     1,     3,     3,     2,    -2,    -8,   -11,   -13,    -9,    -9,   -19,   -20,   -18,   -22,   -21,   -19,    -9,    -5,    -3,     2,     4,    -1,    -1,    -1,    -1,    -1,    -3,     0,    -1,     3,     2,    -4,    -2,    -3,    -4,     0,     3,     3,     0,    -5,    -6,   -11,   -12,   -14,   -11,    -9,    -2,     0,     1,     0,    -1,     0,     4,     0,     4,     4,     2,     6,     1,     5,     1,    -2,    -3,    -3,     2,     2,     2,     2,    -2,     1,     1,    -5,    -3,    -6,    -4,     0,     0,    -1,     1,     0,     2,     5,     2,    -3,    -3,    -1,     2,     0,     3,    -3,    -3,    -5,    -5,     0,     0,     1,     1,     0,     0,     1,     4,    -1,    -3,    -3,    -6,     0,    -2,    -2,     0,     6,     3,     5,     0,    -1,     4,     0,    -2,    -2,    -5,    -4,     1,    -1,    -4,    -2,    -5,    -1,    -2,     4,     2,    10,    -5,    -7,    -4,     0,     2,    -1,    -8,    -5,    -7,     3,    -6,     0,    -2,     4,     4,    -2,    -3,    -3,    -4,    -2,    -9,    -5,     0,     1,    -3,    -1,    -1,     8,     0,    -5,    -6,    -1,    -1,    -1,    -4,    -9,    -7,    -4,    -2,    -3,     1,     3,     0,    -2,    -5,    -1,    -1,    -1,    -4,    -9,    -4,    -2,     1,     2,     1,     0,    -5,    -9,    -8,    -1,    -2,    -4,     5,     0,    -5,     2,     1,    -4,    -1,     1,     1,     0,    -3,    -6,    -8,    -4,    -5,    -2,     3,     2,     2,     3,     1,     1,    -1,    -9,    -9,    -1,     0,     4,     6,    -3,     2,    -2,     0,    -1,    -6,     0,    -2,    -4,    -7,   -13,    -7,    -6,    -6,    -1,     0,     0,     5,    -4,    -4,    -1,     0,   -10,    -8,     1,     0,     7,     6,     3,     0,    -3,    -7,   -11,    -6,    -3,    -8,    -4,   -13,    -7,    -9,    -7,     2,     2,     4,     6,     3,     1,    -4,     6,     0,    -2,    -6,    -1,    -1,     4,     5,     5,    -1,    -5,    -4,    -3,    -1,    -2,    -2,    -3,     1,    -2,     3,     1,     5,     3,     3,     0,     1,     0,    -1,    -3,    -1,    -7,     1,    -1,    -1,    -2,     2,     4,    -1,     1,     0,    -4,    -8,     0,    -2,    -2,     0,    -4,     5,     2,     7,     1,    -2,     0,     3,     4,     6,     2,     7,    -1,     0,    -1,     1,    -5,     2,    -2,     2,     0,    -1,    -2,    -4,    -5,    -2,    -2,    -2,    -4,     5,     5,     1,     1,    -1,     1,     0,     2,    11,     2,    10,    10,     0,     0,    -1,     4,     4,     0,     1,    -1,    -3,     4,     1,    -2,    -1,    -2,     0,     1,    -3,    -3,    -3,    -3,    -4,     5,     1,     5,     5,     3,     7,    12,    -1,    -1,    -1,     0,     5,     7,     3,     5,    -3,    -2,     4,    -2,    -5,    -1,     3,     2,     6,    -5,    -1,    -1,     1,     1,     3,    -2,    -7,    -1,    -3,    -1,     0,    -1,     0,     1,     6,    -5,    -3,     8,     4,     7,     8,     6,    -1,     8,     5,     6,     5,    -4,     0,     4,     7,     6,     5,     9,     6,     4,    -1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     1,     0,     2,     1,     7,     4,     1,   -10,    -5,    -2,     1,    -6,    -4,     1,    -3,    -2,     1,     1,    -1,     1,    -1,     0,     1,     1,    -1,     0,     0,    -1,     1,     0,    -1,     0,     0,    -2,    -2,    -1,     0,     0,    -2,    -5,    -6,    -5,     0,     0,     1,     0,    -1),
		    96 => (   -1,     1,    -1,     0,    -1,     0,    -1,    -1,     1,     0,    -1,    -1,     5,     5,    -1,     0,     1,    -1,     0,     1,     0,     0,     1,     0,     0,     1,     1,    -1,     0,     1,     0,     0,     1,     2,     2,     5,     7,     5,     4,     2,     7,    11,    -3,     2,     5,     7,     6,     2,     5,     3,     3,     2,     1,     0,     1,    -1,     0,     1,     0,     0,     7,     8,     5,     5,     3,     3,     6,     8,    13,     9,     5,     4,     5,     6,     2,     0,     2,    -2,    -1,    -2,     2,     2,     1,     0,    -1,     1,    -1,    10,     0,     1,     9,    10,     6,     4,     6,     1,     3,    10,     6,     4,    -2,    -6,    -4,    -1,     3,    -4,    -2,    -2,    -1,    -2,     0,     1,    -1,     0,    -2,    12,     1,     9,     7,     0,    -1,     2,     2,     2,     5,     1,     0,    -3,    -5,    -1,    -2,    -3,   -10,    -5,    -7,    -8,    -7,    -6,    -1,     2,     0,     0,    -2,    -2,     4,     3,     0,    -3,    -4,     1,     2,     0,     6,     1,    -8,     0,    -8,    -3,    -3,    -7,   -11,   -11,   -13,    -9,    -5,    -3,     2,     2,     1,    -1,    -1,    -6,     3,    -2,    -4,    -8,    -7,     6,     3,     5,     4,     1,    -3,    -9,    -6,    -7,   -15,   -15,   -10,   -15,   -13,   -13,    -6,    -2,     1,    -4,    -1,     0,    -1,    -8,     3,     2,    -6,    -9,     0,     0,     3,     3,     1,     0,    -5,   -10,   -14,   -14,   -17,   -12,    -8,    -2,   -14,   -14,   -10,    -4,     2,    -6,    -1,     0,     1,    -7,     5,     0,    -3,    -2,     4,     3,     1,     0,    -2,     0,   -12,   -20,   -15,    -8,    -9,     0,     1,     3,    -4,    -7,   -10,    -9,     1,    -6,     0,    -1,     0,    -2,     5,    -1,    -5,    -2,     3,    -1,    -1,     2,     0,   -13,    -9,    -7,    -2,    -1,    -1,     7,     8,     7,     4,     2,     0,    -8,    -6,    -3,    -1,    -2,     0,    -2,     2,     2,    -3,     0,     3,    -3,     2,    -2,    -2,   -15,    -9,     0,     2,     7,     6,     3,     4,     2,    -1,    -1,     2,    -3,    -8,    -9,     1,     1,    -1,    -4,     4,     4,    -5,     2,     1,    -2,    -3,    -4,    -6,   -13,    -7,     0,     4,     3,     3,     3,     4,     0,     0,    -1,     1,     1,    -4,    -5,     0,     0,    -2,    -7,     2,    -1,    -1,     0,     2,    -2,    -3,    -3,    -7,    -4,     4,    -4,     5,    -2,     3,     4,     5,     2,     5,     5,     6,     3,    -6,    -5,     0,     0,    -2,    -7,    -2,     4,     2,    -3,     0,    -2,     1,    -6,    -9,    -3,    -1,     0,     3,     0,    -6,     4,     0,     3,     4,     8,     6,     2,    -5,     1,     1,     0,    -2,    -6,    -4,     2,     6,    -2,     4,    -1,     2,     1,    -5,     0,     1,     3,     1,     0,     5,    -4,     2,     2,     5,     7,     1,    11,    -1,     0,    -1,     0,    -2,    -4,    -5,    -2,     5,    -1,     0,     1,     0,    -1,    -1,     4,     4,     1,    -1,    -2,     1,    -3,     2,     3,    -1,    -1,     2,     8,     0,    -7,     0,     0,    -3,    -6,    -2,     1,     4,     1,    -2,     0,     3,     6,    -3,    -1,     3,     0,     1,    -1,    -6,     2,    -3,    -1,    -3,     1,     5,     8,     0,    -4,    -1,     0,     1,    -5,    -3,    -3,     0,    -1,     4,    -3,     0,    -3,    -2,     2,     5,     3,    -2,    -5,    -4,     0,    -7,    -1,    -3,     0,     9,     8,    -1,    -4,     1,     1,     0,    -5,     3,    -3,    -7,     3,     0,    -3,    -9,    -6,    -4,     0,     2,    -2,    -1,     1,    -1,    -2,    -1,    -2,     1,     5,     5,     1,    -3,    -2,     0,    -1,     0,    -2,     5,    -4,    -3,     2,     2,     0,     0,    -7,    -6,    -3,     5,     5,     4,    -2,    -7,    -3,     0,    -2,    -2,     0,     0,     4,    -3,     0,     1,    -1,     0,    -3,     5,     0,    -7,    -2,    -6,    -2,     1,    -4,    -6,    -3,     3,    10,     5,     2,     5,    -3,     4,    -3,    -5,    -5,    -3,     3,     1,     0,     1,    -1,    -1,    -2,     1,    -1,     0,     2,    -5,    -2,    -3,    -5,    -6,     2,     4,     3,     1,     3,    -4,    -7,     1,    -4,    -2,    -5,    -6,    -1,     2,     1,     1,     0,    -1,    -2,    -2,     0,     2,    -7,   -11,    -7,    -5,    -9,    -5,     1,    -1,    -4,    -5,    -3,    -5,    -7,    -4,   -10,   -10,   -11,   -11,    -3,     2,     0,     0,    -1,     0,    -2,    -3,    -1,    -1,    -3,    -5,    -9,   -13,   -10,    -7,    -2,    -2,    -9,   -16,   -17,   -14,    -8,    -2,    -8,    -8,    -5,   -10,     0,    -1,    -1,     1,    -1,    -1,     0,    -1,     0,     0,    -2,    -2,    -1,     0,     2,     0,    -4,    -7,    -7,   -10,    -5,    -8,   -10,    -3,    -2,    -3,     0,    -1,    -1,     0,     0,     1,     1,    -1,     0,     1,     0,    -2,    -2,    -2,    -2,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -3,    -7,    -3,    -5,    -4,    -1,     1,     0,     1,     1,     1,     0,    -1,    -1,     0,     1,    -2,    -1,    -1,    -1,    -3,    -2,    -1,    -3,    -2,    -1,    -1,    -2,     0,    -2,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,    -1,     0,     1,     0,     1,    -1,    -3,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     1,    -1,    -1,     0,    -1),
		    97 => (    0,     1,     1,    -1,     1,    -1,     1,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     1,     0,     0,    -1,     1,    -1,     0,     0,     0,     0,     1,     0,     1,    -1,    -1,    -1,     1,    -1,     0,    -1,    -5,    -3,    -3,     1,    -2,    -6,    -8,     0,    -2,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     1,     0,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -5,    -5,   -10,    -1,    -1,    -2,    -4,    -2,     0,    -1,     0,    -2,    -2,    -3,    -3,     0,     0,     0,     0,     0,    -1,     1,    -2,    -1,    -6,    -6,   -13,   -11,   -10,   -11,   -14,   -12,   -14,    -7,    -3,    -3,    -3,     0,    -4,    -5,    -6,    -9,    -3,    -2,    -3,    -1,     0,     0,     0,    -1,    -2,    -7,    -9,   -10,   -11,   -17,   -17,   -16,    -9,    -9,    -9,    -8,    -6,   -12,    -9,    -6,    -6,    -7,    -4,    -7,   -13,   -14,    -7,    -3,     1,     0,     0,     1,    -8,   -14,     3,    -7,    -2,     2,     3,    -5,    -3,     1,     4,     5,    -1,     5,     2,     0,    -6,   -11,    -7,    -5,   -15,   -10,   -13,    -6,     0,     0,     0,     5,     5,     4,    -4,    -3,    -3,    -4,     0,    -1,     0,     2,     1,     2,     5,    -1,    -3,    -1,     1,     6,     4,     5,    -6,   -10,    -8,    -8,    -5,    -1,     6,     6,     2,     5,    -5,    -3,     1,    -2,     0,    -2,     2,     3,     1,     2,    -3,    -3,     9,     1,    -2,     1,    -1,    -1,    -2,     0,    -8,   -11,    -6,    -6,    13,     3,    -1,     3,     0,    -4,     2,     3,     5,     5,     3,     0,    -2,    -3,     0,    -2,     3,     6,     2,     4,     0,    -3,    -4,    -4,   -13,   -15,    -4,     1,     6,    -2,     1,     4,     3,     4,     1,     4,     8,     7,     1,    -6,    -3,     3,     3,     0,     4,     4,     0,     5,     0,     3,    -3,    -6,    -1,    -1,    13,     1,     5,     3,     0,     4,     3,    -1,     4,     7,     4,     4,    -5,    -8,    -2,     4,     8,     4,     0,     3,     2,     6,     0,    -2,    -5,    -5,     3,     0,    11,    -1,     1,     8,     2,    -2,    -1,    -1,     2,     4,     3,    -4,    -4,     3,     6,    11,     7,     5,     0,     4,    -3,     2,    -3,     0,     3,     2,    -9,    -5,     7,     0,     4,     8,     2,    -4,    -4,    -1,    -1,     3,     1,     2,     6,     5,     6,    11,    10,     6,     3,     1,    -6,    -2,     0,     8,     0,     3,     6,     4,     6,     0,     2,     8,     0,    -6,    -4,     2,    -1,     0,     2,     0,     4,     5,     4,    13,     8,     5,     2,    -5,    -5,    -9,    -3,     1,    -3,     0,     6,    -2,    -5,    -1,     3,     3,    -5,    -8,    -1,    -2,    -4,    -1,     1,    -3,     2,     1,     2,     7,     2,     2,     3,    -3,    -3,    -4,    -8,    -2,     1,     5,    -5,    -6,     0,    -1,     0,     2,    -5,    -6,    -1,     1,    -2,    -9,    -8,    -3,    -2,    -3,     1,    -2,    -4,     0,     3,     7,    -2,     1,     1,     7,     5,     4,     2,    -3,    -4,     0,    -2,    -1,    -4,    -2,    -1,     0,    -1,     0,     5,     4,    -3,    -8,    -5,    -4,    -2,    -2,     9,    13,    10,     3,     8,     5,     8,     6,    -6,    -5,    -5,     0,    -2,    -2,    -3,     0,     1,     0,    -4,     0,     0,     0,    -6,    -9,    -3,     0,     0,     6,     9,    11,     2,     6,     4,     8,     6,     1,     4,    -1,    -7,     2,     1,     2,    -2,    -1,     5,     4,    -2,    -4,    -6,    -2,    -5,    -5,    -3,    -2,     1,     2,    13,     7,     4,     2,     1,     4,     2,     0,     1,     1,    -5,    -1,     2,     1,    -1,     2,     3,     3,     1,     3,    -5,    -3,    -3,    -5,    -7,    -3,    -3,     7,    13,     5,     4,     1,     2,     1,    -1,     4,    -1,    -5,    -2,     1,     3,    -1,    -3,    -8,     2,     0,     3,     3,     1,    -2,    -2,    -3,     0,     0,     2,     0,     3,    -1,     0,    -1,    -1,    -3,    -3,     3,    -3,    -6,     1,     0,     1,    -1,    -3,    -5,     5,     4,     4,     3,     5,     5,     1,     2,     1,    -2,     3,     1,    -4,    -6,    -5,    -3,     2,    -2,    -2,    -5,    -4,    -2,     1,     0,     0,    -3,    -5,    -6,     3,     8,     4,     1,     1,     3,    -1,     3,     2,    -2,    -5,    -1,    -7,    -5,    -6,    -6,    -5,    -9,    -9,    -6,     1,    -6,    -1,    -1,     1,    -2,   -10,    -5,     4,     7,     5,     3,     0,     5,     0,    -2,     0,   -10,    -8,    -3,    -7,    -9,    -7,    -5,    -5,   -10,    -9,    -3,     1,    -5,     1,     0,     1,     0,    -1,    -1,     5,     2,     5,     0,     0,     0,     1,    -1,     0,    -6,    -7,    -5,    -4,   -10,    -9,    -8,    -2,    -9,   -10,    -6,    -5,    -1,     1,    -1,    -1,    -3,     6,    -1,     0,     1,     2,    -4,     2,     2,    -1,    -2,     1,    -9,    -8,     0,    -6,    -8,   -10,    -7,    -2,     0,    -7,    -3,    -1,    -1,     0,    -1,    -1,    -1,    -7,    -4,    -6,    -3,    -3,     1,     7,    -1,    -2,    -1,    -1,     0,     1,    -2,    -6,    -2,    -2,     0,     3,     0,     0,    -1,     0,     1,     1,     0,     1,    -1,     0,     3,     3,     0,    -3,    -2,     0,     0,    -5,    -2,    -3,    -5,     2,     0,     7,     3,    -3,     0,     4,     0,     5,    -1,     0,     0,    -1),
		    98 => (    1,    -1,    -1,     0,     1,    -1,     0,     1,     0,     0,     0,    -1,     1,    -1,     0,    -1,    -1,     0,     1,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     1,    -1,     0,     1,     1,     1,     1,     0,     1,    -1,    -2,    -2,    -5,    -4,    -5,    -2,     1,    -2,    -1,     0,    -1,    -1,    -1,    -1,     1,     1,     1,    -1,     0,     0,     0,     1,     0,    -3,    -7,   -10,    -9,    -3,    -1,    -2,    -6,    -6,    -2,    -1,     0,    -1,    -2,    -4,    -2,     0,     0,     0,     0,     1,     1,    -1,    -1,    -2,    -4,    -3,   -12,     4,     6,     8,     3,     7,     8,     5,     3,     1,     3,    -2,    -6,    -5,    -7,    -4,     0,    -2,    -2,    -1,    -1,     0,    -2,     1,    -1,    -8,    -9,    -2,     2,     3,     3,    -2,    -6,     1,    -2,    -1,    -2,    -1,     0,    -1,     2,     0,     2,    -8,    -4,    -2,     0,     1,    -2,     0,    -1,     0,    -6,    -8,   -14,    -4,     2,     3,    -3,     0,     1,    -7,    -4,     3,    -1,     2,     5,     3,     0,     4,     0,    -3,    -5,    -4,    -1,     2,    -1,     1,     0,    -7,    -4,    -3,    -4,     0,    10,     5,     3,     3,     2,     0,     2,     3,     4,     3,     0,    -4,     3,    -3,    -1,    -4,    -1,    -4,    -3,     0,     0,    -1,    -5,    -3,    -6,    -2,     0,     6,     9,    -5,    -2,     2,    -4,    -1,    -4,    -3,    -3,    -4,    -1,     0,     2,    -1,    -6,    -3,    -5,    -2,    -2,    -2,    -2,    -1,    -3,    -5,    -3,    -8,    -7,     2,     9,    -3,    -2,     5,     3,    -3,    -6,    -6,    -3,    -9,     1,     0,     1,    -2,    -2,    -1,    -6,     0,     3,     3,     0,     1,    -1,    -2,    -2,    -9,    -7,    -1,    -3,    -3,     1,     6,     7,     3,    -3,    -4,    -2,    -1,     5,    -5,    -1,     0,     3,    -1,    -3,    -2,     1,    -8,    -7,     1,    -2,    -4,    -4,    -4,    -9,     3,    -4,   -12,    -3,     4,    13,    12,     8,     3,    -1,     1,     2,     2,    -6,     5,     3,     1,    -5,    -9,   -10,    -8,    -8,     0,    -1,    -1,    -5,    -3,    -4,     0,    -1,    -4,    -1,    -9,     1,     6,    10,     7,     0,    -2,    -5,    -2,    -2,    -1,    -2,    -4,    -4,    -9,    -7,    -2,    -3,     0,     1,    -2,    -1,    -2,    -5,    -3,    -7,   -10,   -10,   -12,   -12,     1,     1,     2,     8,     2,    -1,     2,     3,     1,     2,     2,    -1,    -1,    -5,    -4,    -3,    -1,     0,    -3,    -1,    -3,    -2,    -1,    -6,   -10,   -14,   -11,    -8,    -6,     0,     0,     5,     2,    -2,    -1,    -3,    -7,     0,     2,    -7,    -6,    -5,    -4,    -1,    -1,    -1,     0,    -6,    -3,     1,     0,    -4,    -5,    -7,    -1,     3,     2,     1,    -1,    -4,     0,     1,     0,    -5,    -3,     3,    -2,    -7,    -7,    -4,    -8,    -4,    -1,     1,    -4,    -4,    -6,    -3,    -4,     0,    -2,     1,     0,     3,    -2,    -5,    -3,    -1,     4,    -3,    -5,     0,     0,     3,    -6,    -4,    -5,    -4,    -9,    -3,     0,    -1,    -2,    -2,    -4,    -1,     5,     4,     1,     6,     1,     0,    -5,    -1,    -8,     0,    -8,     5,    -4,     5,     5,     2,    -3,    -1,    -3,    -2,   -11,    -4,     1,    -1,    -3,    -9,     3,     1,    -3,     5,     4,     1,    -3,    -1,    -2,    -9,    -8,    -2,    -6,    -2,     2,     6,     2,     7,     5,     0,    -5,    -4,    -2,    -5,    -1,    -1,    -2,    -3,     8,     0,     2,     5,    -1,    -5,    -3,     2,    -3,    -8,    -3,    -3,   -11,    -4,     2,     4,     3,     3,     3,     2,    -7,    -4,     0,    -3,     0,    -2,    -5,     5,     6,     8,     6,     3,    -6,    -3,     1,     2,    -8,    -5,    -6,    -2,    -3,    -1,    -3,     0,     2,     3,     1,    -5,    -7,    -3,    -9,    -3,    -1,     0,    -4,     1,     5,     3,     4,     3,    -2,    -7,    -1,     1,    -6,    -1,    -1,     2,     3,    -3,    -4,    -3,     4,     3,     2,    -4,    -3,    -1,    -8,    -1,    -3,    -2,    -5,    -5,     1,     0,     0,    -1,    -4,     0,    -3,    -1,     1,    -3,     4,    -2,    -3,    -5,    -8,     2,     4,     4,    -1,    -3,    -5,    -3,    -7,    -1,    -3,    -2,    -4,    -6,    -5,     1,     7,     5,    -4,    -3,     1,     2,     3,    -5,    -1,    -6,    -4,    -2,    -4,    -2,     1,    -2,    -7,    -3,     0,    -1,    -4,     0,    -1,     1,    -1,    -2,    -7,     4,     1,     6,     1,    -5,    -3,    -5,     1,    -1,     0,    -2,    -2,    -5,    -2,     0,    -3,   -10,    -4,    -2,     0,     4,    -7,    -1,    -1,    -1,    -3,    -2,    -5,    -6,     3,     2,     2,     0,    -4,    -4,    -1,     0,     3,     4,     6,    -4,     1,    -1,     0,    -4,    -4,    -1,    -5,    -1,    -2,     0,     0,     1,    -1,     0,    -1,    -4,     0,    -2,    -6,    -4,    -6,    -7,    -6,    -7,    -7,    -8,    -6,    -3,    -1,     0,     0,    -3,    -1,    -1,    -1,     0,    -1,     1,     0,    -1,    -1,    -3,    -2,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -5,    -6,    -7,    -4,    -3,    -2,    -2,    -5,    -8,    -8,    -4,     1,     0,    -1,     1,     0,    -1,     0,     1,     0,    -2,    -1,    -3,    -1,    -2,    -2,    -1,    -1,     0,    -4,    -1,    -1,    -2,    -2,    -2,    -1,     0,    -1,     1,    -1,    -1,    -1,    -1,     0),
		    99 => (    0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     0,     0,    -1,     1,     1,     0,     1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     1,     1,     0,    -1,     0,    -2,    -3,    -4,    -4,     1,    -1,     0,    -1,    -2,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -2,     0,     1,    -3,     0,     0,     0,    -1,     0,    -2,    -2,    -3,     0,     0,     0,    -1,     0,     1,     0,     0,    -3,    -1,    -2,    -2,    -1,    -4,    -3,    -2,     0,     1,    -1,    -2,     0,    -1,    -2,    -2,    -2,    -4,    -1,    -4,    -2,    -4,    -3,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -7,    -1,     1,     0,     0,    -2,    -5,    -5,    -2,    -6,    -3,    -5,    -3,    -7,    -9,    -1,    -1,    -1,     0,    -6,    -2,    -1,     1,     1,    -1,    -3,    -1,     0,     0,    -2,    -2,    -3,    -2,    -4,    -5,    -7,    -8,    -9,    -6,    -2,    -1,     3,    -4,    -3,    -3,    -2,    -1,    -2,    -3,     1,    -1,     1,     0,    -3,    -1,    -3,    -4,    -3,    -6,    -2,    -4,     0,    -1,    -1,     0,     0,    -4,    -7,    -2,    -4,    -5,    -4,    -4,    -2,    -2,     0,    -2,    -3,     1,    -1,    -1,    -2,    -2,    -4,    -7,    -9,    -9,    -5,    -4,     1,     0,     3,     1,     2,     3,    -5,    -2,    -5,    -4,    -8,    -4,     3,    -3,    -1,    -1,    -2,    -4,    -4,    -2,    -2,    -5,    -6,    -7,   -10,    -7,    -5,     0,     1,     1,    -2,     1,     0,     5,    -4,    -2,     2,    -1,     0,    -5,     0,    -1,    -6,    -1,     0,     0,    -5,    -4,    -4,    -6,    -4,    -7,    -2,     1,    -2,     0,     2,     3,     2,     2,     8,     2,    -2,     1,     5,     1,     0,     0,    -1,    -3,    -4,    -3,    -2,    -1,    -5,    -4,     0,    -3,    -4,    -6,    -3,     1,    -4,    -6,     3,     3,     2,     5,     1,     3,    -3,     5,     4,    -1,     1,    -1,    -5,    -4,    -4,    -2,    -3,     0,   -10,     6,     0,    -2,    -3,    -3,     0,     0,    -3,    -8,     0,     1,     4,     2,    -1,    -4,    -5,     0,     1,     1,    -2,     0,    -2,    -6,    -6,    -1,    -2,     0,    -5,     2,     6,     5,     0,     3,     0,    -3,   -10,    -6,    -1,    -2,    -3,     0,     0,    -2,     0,    -1,     3,     0,     4,    -1,    -1,    -6,    -3,    -5,    -1,     1,    -5,    -2,     3,     3,     2,     3,    -1,    -4,   -12,    -3,    -2,    -8,    -8,    -5,     1,     0,    -5,     1,     1,    -3,     4,     1,    -3,    -7,    -5,    -2,     0,     0,    -3,    -4,     4,     3,     3,    -1,    -1,    -8,    -7,    -2,    -2,    -5,    -6,    -7,    -1,    -2,    -4,     0,     1,     3,     3,    -2,    -5,    -6,    -4,     0,     0,    -1,     1,    -6,     4,     6,     2,     2,     0,    -5,    -8,    -2,    -4,    -5,    -1,    -1,     0,     0,    -7,     1,    -1,    -1,     2,     2,    -6,    -7,    -4,     0,    -2,     0,    -2,    -4,     4,     7,     5,     8,     3,     1,     2,     1,    -5,     1,     0,     1,     0,    -7,    -5,    -4,    -5,     0,    -1,     5,     3,    -6,    -1,    -3,    -1,     0,    -1,   -10,    -1,    -1,     0,     3,     5,     7,     5,     4,     6,     4,    -1,    -2,    -4,    -6,    -7,    -1,    -3,    -3,    -1,     4,    -1,    -6,    -2,    -4,    -4,    -1,     0,    -9,     3,    -3,    -5,    -1,     2,    -1,    -1,     6,     1,    -1,    -7,    -2,     0,    -2,    -2,    -1,    -6,    -1,    -3,     4,     3,    -3,    -1,    -5,    -3,    -1,    -1,    -5,     4,     0,    -5,    -5,    -3,    -7,    -6,    -2,    -2,     1,    -8,     2,     0,    -3,    -3,    -2,    -8,     0,    -5,    -1,     5,     5,     4,    -4,    -1,    -1,     0,    -2,     4,     3,    -1,    -4,    -5,    -7,    -4,    -6,    -3,    -9,    -6,     3,     2,    -4,    -7,    -2,    -4,     1,     0,    -2,     5,     6,    10,    -5,    -1,     0,     1,    -3,     1,     2,    -1,    -3,    -3,    -4,    -7,    -4,    -2,    -1,    -4,     4,    -3,   -13,    -3,    -1,    -2,    -2,     4,    -4,     0,     2,     6,    -6,    -1,     0,     1,    -4,    -3,    -5,    -2,    -3,    -4,    -3,    -4,    -2,    -4,    -1,    -1,     6,    -7,    -8,    -1,     0,    -2,     0,     1,    -1,     1,    -2,    -6,    -1,    -1,     0,     0,    -3,    -3,    -3,    -1,    -2,    -2,    -2,    -1,    -3,    -1,     0,     0,     2,    -3,     1,     2,    -1,    -3,     5,     0,     6,     2,     0,    -3,    -2,    -1,     0,    -1,    -3,    -1,    -4,    -2,     0,     2,    -5,    -5,    -3,    -2,     0,    -1,     2,     2,     4,    -2,    -1,    -1,     4,     3,     4,     2,     0,    -1,    -1,     1,     0,    -1,     7,    -5,     0,     3,     1,     0,    -6,    -2,    -2,     0,    -2,    -4,     4,     3,     2,    -1,    -2,     2,     5,     3,     4,     1,    -2,    -1,    -1,    -1,     0,     0,     1,     7,     4,     3,     3,     0,     1,     4,    -4,    -1,    -2,    -5,     0,     2,    -1,    -1,    -1,     3,     5,     8,     4,     0,     2,     1,     1,     0,     0,    -1,    -1,     0,    -3,    -1,     2,     5,     4,     4,     0,     1,    -1,    -4,    -1,    -1,    -1,    -1,    -3,    -2,    -2,    -1,     2,    -3,     1,    -1,     0,     0)
        );

 ---------------------------------INFO-
 -- COEF =10.784521

 -- MIN =-31.999998
 -- MAX =21.19651

 -- SUMMIN =-2273.605
 -- SUMMAX =1653.0385
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
