----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,     0,     1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -1,     1,     1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,     1,     1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,     1,     1,    -2,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,    -1,     0,     1,    -1,     0,    -1,    -2,     0,    -1,     0,    -2,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,    -1,    -1,     0,    -1,     0,     2,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     0,     0,     0,     1,     0,    -1,    -2,     0,     1,     2,     0,     0,     1,     0,    -2,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,    -1,    -3,    -2,     0,     1,     1,     0,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,     0,     0,     1,     1,     0,    -2,    -2,     0,     0,     1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,     0,     1,     2,     0,    -3,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -1,    -1,    -1,     1,     1,    -1,    -3,     0,     0,     2,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,     1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -2,     0,     0,     1,    -1,    -2,    -1,     0,     1,     0,     0,     1,    -1,     0,     0,    -1,    -1,    -2,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     1,     1,    -1,    -1,    -3,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     1,     1,     0,    -1,    -1,     1,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,    -2,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,     1,     1,     1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,     1,     0,     1,     1,    -1,    -1,    -1,    -2,     0,    -1,    -1,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,    -2,    -1,    -1,     0,     2,     0,     0,    -1,    -1,     0,    -1,    -1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0),
		     1 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,     0,     1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     2,     1,     0,     0,     0,     2,     1,     1,     1,     0,     0,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,     0,     1,     0,     0,     0,     1,     0,     1,    -1,    -3,    -1,    -2,    -1,    -1,     0,     0,     1,     2,     1,     0,    -1,    -1,    -3,    -1,    -1,    -2,    -3,    -1,     0,     2,     0,     0,     0,     1,     1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     1,     1,    -1,     0,     0,    -2,     0,     0,    -2,    -2,    -1,    -1,    -1,     0,     1,     0,     1,    -1,    -1,     0,    -3,    -2,    -1,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,    -1,    -3,    -1,    -1,    -2,    -2,     0,     1,     0,     1,     0,     1,     0,    -1,    -1,     0,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -3,    -3,     0,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -4,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -1,     0,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,     0,    -2,    -2,    -1,     0,     1,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -2,     0,     2,     0,     0,     0,     1,     1,     0,    -1,    -1,    -2,    -3,    -1,    -2,    -1,    -1,     0,     2,     0,    -2,    -1,    -1,    -1,     0,     0,    -1,    -2,    -2,     0,     2,     0,     0,    -1,     1,     0,     0,     0,     0,    -3,    -2,    -1,    -1,     0,    -1,     1,     0,     1,    -3,    -3,    -1,     1,     2,     2,     1,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,    -3,    -1,    -1,     0,     0,     1,    -1,     0,    -2,    -3,     0,     1,     0,     0,    -2,    -1,     0,     1,     0,     0,     0,     1,     1,     1,    -2,    -1,    -1,     0,    -2,    -1,     0,     0,    -1,     1,     0,    -1,    -2,     0,     1,     2,     2,     1,    -1,    -1,     2,     2,     0,     0,     0,     1,     2,     1,     0,     0,     0,     1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,     0,     2,     1,    -1,    -3,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,     1,     1,     1,     1,    -1,     0,     0,    -2,    -2,    -2,     0,     2,     1,     2,     2,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     2,     2,     2,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,    -1,    -2,    -2,     0,     1,     1,     1,     0,     0,     0,     1,     1,     0,     1,     0,     0,     1,     1,    -1,     1,     1,     0,     0,    -1,     0,     1,     0,     1,    -1,    -2,    -3,     0,     1,     0,     0,     0,    -1,     0,     1,     2,     0,     1,     0,     0,     1,     0,     0,     2,     1,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -2,    -2,    -1,    -1,     0,     1,    -1,    -1,     0,     1,     1,     1,     0,     1,     1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     1,    -1,     0,    -1,    -2,    -2,    -2,    -1,     1,     0,     0,     1,     1,     1,     0,     0,     1,     1,     0,     0,     0,    -1,    -3,     0,     0,    -1,     1,    -1,     0,     0,     1,    -1,    -1,    -2,     0,     1,     2,     1,     1,     1,     1,     2,     3,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     1,    -1,     0,     1,     0,     0,     1,     0,     0,     0,     1,     2,     2,     0,     0,     0,     1,     1,     2,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -2,     1,     1,     0,     0,     0,     3,     2,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,    -2,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -2,    -2,    -2,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		     2 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,     0,    -1,    -1,    -1,    -1,    -3,    -1,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,    -1,     0,     1,     1,     0,    -1,    -2,    -1,    -2,    -2,    -1,     1,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,     1,     0,     0,    -1,     1,     1,     0,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,     2,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -1,     0,     0,     1,     1,     1,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,    -2,    -2,    -1,    -1,     1,     1,     1,     0,     0,     0,    -2,    -2,     2,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,     1,     0,     0,     0,     1,     0,     1,    -1,    -1,    -1,    -1,    -2,     0,     1,     0,     0,    -3,     0,     2,    -1,     0,    -2,     2,     1,    -1,    -1,     1,     0,     0,    -1,    -2,     0,     1,     0,     0,     1,    -2,    -3,    -1,    -1,     0,     1,     0,     0,     0,     0,     1,    -2,     0,     0,    -1,     2,    -1,    -1,     0,     0,     0,    -1,    -1,     1,    -1,    -1,     0,     1,     0,    -1,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,     1,    -1,     0,    -1,     1,    -2,    -1,     1,     1,     1,     0,     0,     0,     0,     1,     2,     3,     1,    -1,    -1,     0,     1,     0,     1,     0,    -1,    -1,    -1,     1,    -1,     0,    -1,    -1,    -1,     1,     0,     1,     2,     1,     1,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -3,    -1,     1,     1,     1,     1,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,     0,    -2,     0,     0,     2,     0,     0,     0,     0,     1,     0,    -1,    -2,    -2,    -3,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,     3,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -2,    -2,    -2,     1,     1,    -1,    -2,    -1,     1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     1,     2,     1,     0,     0,     0,     0,     1,     0,    -1,    -3,    -1,    -1,     0,     0,     1,     1,     0,     1,    -1,     1,     1,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,     0,     0,     1,     1,     0,    -1,     0,    -1,     0,     0,     0,     1,     0,     1,     2,     1,     2,     0,    -2,    -3,    -2,    -1,     0,    -1,     0,     1,     1,     0,     0,     1,     1,     0,     1,     0,    -1,     0,     0,     1,    -1,     2,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     2,     0,     0,    -1,     2,     1,     2,     1,     0,    -1,     0,     0,    -1,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     2,     0,     2,     3,     0,     0,     0,     2,     2,     1,     1,     0,     0,    -1,     1,     1,     1,     0,     0,     0,     1,     1,     0,    -1,    -1,     0,     1,     1,     2,     1,     2,     2,     0,     0,     0,     1,     1,     1,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     1,     1,    -1,     0,     0,    -1,     0,    -1,     1,     2,     1,     2,     0,     0,     0,     0,     0,     1,     2,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     1,     2,     2,     1,    -1,     0,     1,     1,     1,     2,     0,     0,     0,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -3,    -1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,     1,     1,     1,     0,     0,    -1,     0,    -1,    -2,    -1,    -2,    -2,    -1,     0,    -2,    -4,    -1,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,    -1,     1,    -1,    -1,     0,    -1,     0,    -2,    -3,    -2,    -2,    -2,    -1,    -1,    -3,    -4,    -2,     1,     0,     1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -2,    -2,    -2,    -1,    -1,    -2,     0,    -1,    -2,    -1,    -3,    -3,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -3,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -3,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0),
		     3 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -3,    -2,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     1,     1,    -1,     0,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     1,     1,     2,     1,     0,     0,     1,     1,     0,    -1,     0,     1,     0,     0,    -2,    -1,    -4,    -3,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     1,     1,     0,     0,     0,     0,     0,     1,     1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     1,     2,     1,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,    -1,    -1,     2,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     1,     1,     0,     0,     0,     1,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,     0,     2,     1,     0,    -1,     1,     0,    -2,     1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -3,    -4,    -1,    -1,     0,     0,    -1,     2,     2,     0,    -2,    -1,     0,    -1,     0,    -1,    -1,    -2,    -3,    -5,    -2,     0,     0,     0,     1,     1,     0,     0,    -2,    -5,    -2,    -2,     0,     0,    -1,     3,     1,    -1,    -2,    -3,    -4,    -3,    -3,    -3,    -5,    -4,    -4,    -2,    -1,     0,    -1,     0,     0,     0,     1,     1,    -1,    -4,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -4,    -3,    -4,    -5,    -3,    -3,    -1,     1,     2,     2,     0,     1,     0,     1,     2,     1,     1,    -2,    -2,    -2,    -1,     0,     0,     0,    -1,    -2,     1,    -1,    -1,    -2,    -1,    -2,    -1,     0,     2,     2,     1,     0,     0,    -1,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,     0,     2,     1,     0,    -1,     0,    -1,     0,     1,     1,     1,    -1,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     2,    -1,    -1,     2,     1,     0,     1,     1,     1,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,    -1,    -2,    -3,    -1,    -1,    -1,     1,     1,     0,     1,     0,    -2,    -3,    -2,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,    -2,     0,    -1,    -1,     2,     0,     0,     0,     1,     1,     1,     0,    -3,    -3,    -4,    -2,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     1,     0,     1,    -1,    -1,    -2,    -1,     1,     0,     0,     0,     2,     0,    -2,     0,    -2,    -1,    -3,    -5,    -6,    -2,    -3,    -3,    -1,    -1,     1,     1,     1,     0,     0,     1,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,     2,     1,    -1,     1,     0,     1,     0,    -1,    -2,    -1,    -3,    -3,    -1,     0,    -1,     0,     0,     1,     1,     1,     0,    -3,    -4,    -1,    -1,    -1,     0,     0,    -1,     2,     0,     0,     1,     0,     1,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -1,    -1,    -1,     0,     0,    -2,     2,     2,     0,     0,     0,     1,     0,     1,     1,     1,     1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     1,     2,     0,    -1,     0,     1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -2,    -1,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,    -1,     0,     1,     1,     1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     0,    -2,    -2,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     1,     1,     0,     2,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,     0,     2,     0,     0,     2,    -1,    -2,    -3,    -3,    -1,    -2,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -3,    -1,    -2,     1,     2,     1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0),
		     4 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -3,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -2,     0,     0,     2,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -1,     2,     1,     0,     1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,    -3,    -3,     0,    -1,     0,    -1,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     1,    -1,     1,     1,     0,    -1,    -2,    -4,    -4,    -2,    -1,     0,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,     1,     0,     0,     0,     1,     1,    -2,    -3,    -5,    -2,    -1,     2,     2,     2,     1,     0,    -1,    -2,    -2,     0,     0,    -2,    -1,    -3,     0,     0,     1,     1,     1,     0,     1,     2,     0,    -1,     0,    -4,    -3,    -1,     2,     1,     1,    -1,    -1,     1,     0,    -1,    -1,     0,    -2,    -2,     0,    -2,     0,     0,     2,     1,    -2,     0,     1,     0,     1,     1,     1,    -2,    -3,     0,     3,     0,     0,     0,    -1,    -1,    -1,     0,    -2,     0,    -2,    -1,     0,    -1,     0,     1,     1,     0,    -4,    -1,     1,     1,     0,     1,     1,    -2,    -2,     1,     1,     0,     1,     1,    -1,    -2,    -1,    -2,    -2,     1,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     1,     1,     0,    -3,    -3,     0,     1,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,     0,    -1,    -2,     0,    -1,     1,     1,     1,     1,     0,     0,    -1,    -1,     1,     0,     0,    -1,    -2,     1,     0,     0,     0,     0,    -1,     0,     1,     3,     3,     2,    -2,    -1,     0,    -1,    -1,     0,     1,     1,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     1,     3,     1,     0,     0,    -2,     0,     0,     0,    -1,     0,     1,     2,     0,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     1,     1,     0,     2,     1,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,     2,     0,     0,     1,     0,     0,     0,     0,     0,     1,     1,     1,     1,     0,     1,     1,     0,     0,     1,    -1,    -2,    -2,     1,     0,     0,     0,    -2,     1,     2,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     1,     0,     0,     1,    -1,    -2,     0,    -1,    -1,     0,     0,     0,     2,     1,     2,     0,    -2,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     2,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,    -2,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,    -2,     1,    -1,     0,    -1,     2,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -3,    -2,    -2,     0,    -1,    -2,    -1,     1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,    -3,     0,     0,    -1,    -1,     0,    -2,    -1,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,     1,     0,    -2,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -2,     0,    -2,    -2,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     0,     0,     1,     0,     0,     0,     0,    -1,     0,    -1,     1,     1,     0,    -3,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,    -1,    -2,     0,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     2,     0,     1,     1,     2,    -1,     0,     0,     0,     0,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -4,    -2,    -1,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     1,     0,    -1,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,    -2,    -3,    -3,    -2,    -1,    -2,    -3,    -1,    -2,    -2,    -3,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0),
		     5 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -1,     1,     1,     1,     2,     1,     2,     1,     1,     2,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,    -2,    -2,    -1,    -1,    -1,     1,    -1,    -2,    -2,     0,     0,     1,     1,    -1,     0,     1,     1,     1,     0,     0,     0,    -1,     0,    -2,    -2,    -2,    -2,    -3,    -1,    -3,    -2,    -2,     0,     2,     0,     1,     0,     0,     0,     0,     1,     1,     1,     2,     3,     1,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -3,    -2,     0,     0,     1,     0,     0,     0,     1,     1,     1,     0,     2,     2,     1,     2,     2,     3,     1,     0,     0,     0,     1,     0,    -1,    -3,    -3,    -2,    -1,    -1,     0,     0,     2,     0,     0,     0,     1,     1,     2,     0,     2,     0,     0,     2,     1,     2,     1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     1,     1,     0,    -1,    -1,     0,     1,     1,     0,     1,     0,    -1,     0,    -1,     1,     1,     1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -2,     1,     2,     1,    -1,    -1,    -2,    -4,    -2,    -2,    -5,    -2,    -3,    -2,    -1,     0,     0,     1,     0,     0,     0,    -2,    -2,    -2,     0,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -5,    -6,    -7,    -7,    -7,    -5,    -4,    -4,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     0,    -1,    -4,    -4,    -4,    -4,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     1,     0,     1,    -1,    -2,    -4,    -3,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,     0,     1,     2,     1,     0,     1,     0,     0,     0,    -1,     0,     0,     1,    -1,    -1,    -1,     0,     0,    -1,     1,     0,     0,     0,     1,    -1,    -2,    -2,     0,     0,     1,     0,     0,    -1,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     1,    -1,    -2,    -1,    -2,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -2,    -3,    -4,    -3,    -2,     0,     0,    -1,     0,     0,     2,     0,     1,     0,     1,     1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,     0,    -1,    -1,    -1,    -3,    -1,    -3,    -4,    -1,    -2,    -2,    -2,     0,    -1,    -1,     2,     1,     1,     1,     0,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     1,    -1,     0,    -1,    -3,    -2,     0,    -1,     0,     0,     1,    -1,     0,     1,     0,    -1,    -2,     0,    -2,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,     1,     1,     0,     1,     1,     0,     1,     0,     1,     0,     1,     0,     0,    -1,     0,    -1,    -2,     0,     0,    -1,     0,     0,     1,     0,     3,     0,     0,     0,     2,     1,     0,     0,    -1,     1,     1,     0,     0,     0,    -1,     1,     1,    -1,     1,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     2,     2,     0,     0,     0,     0,     1,     1,     1,     1,     0,     0,     1,    -1,    -1,     1,     1,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     2,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,     2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,    -1,    -1,     0,     0,     2,     1,     0,    -1,    -1,    -1,     0,     2,     0,    -2,    -1,    -1,    -1,    -1,     0,     1,    -2,    -3,     0,     0,     0,     0,    -1,     0,     1,     1,     3,     2,     0,     1,     2,     0,     1,     0,     1,    -1,    -2,    -1,    -1,    -2,     0,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,    -1,     0,     1,     2,     0,     1,     1,     1,     0,     0,    -1,     0,    -1,    -2,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0),
		     6 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     2,     1,     1,     1,     1,     0,     0,     1,     1,     0,     1,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,     0,     0,    -1,     1,     2,     1,     1,     2,     1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     3,     2,     0,     1,     2,     0,     0,    -1,     0,     1,     1,     1,    -1,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     1,     1,    -1,     0,     0,     1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,     2,     1,     1,    -1,    -2,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     1,     0,    -1,     1,     1,     0,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,    -1,    -1,    -2,    -2,     0,    -1,     0,    -2,     1,     2,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -2,    -2,     0,    -1,     1,     0,     0,     0,     0,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,     2,     1,     0,     1,    -1,    -1,    -1,    -3,    -2,    -2,    -1,    -2,    -3,    -2,    -1,     1,    -2,     0,     0,     0,    -1,    -1,    -3,     0,    -1,    -1,     1,     0,     0,     1,     0,    -1,    -2,    -2,    -4,    -3,    -3,    -2,    -2,    -4,    -3,    -3,    -2,    -1,    -1,     0,     0,    -1,    -1,    -1,    -3,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -3,    -2,    -4,    -4,    -3,    -2,    -3,    -3,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,    -3,    -2,     0,     1,     0,    -1,     0,     1,    -1,    -3,    -3,    -1,     1,     0,    -2,    -1,    -1,    -1,    -1,     0,     1,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     1,    -2,    -2,    -1,     1,     1,     1,    -1,     0,    -2,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     1,     0,    -1,     0,    -1,    -3,    -1,     0,     1,     0,     0,     1,     1,     0,    -1,    -1,     1,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,     0,     2,     1,    -2,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     2,     1,     0,     1,     0,    -1,    -1,     1,     0,     0,     0,    -1,    -3,    -1,     1,     1,     0,     0,     1,     1,     0,     0,     1,     0,     1,    -1,     1,     1,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,     0,     2,     1,     0,     0,     0,     2,     0,    -1,     1,     0,     0,    -1,     1,     0,     0,     1,     2,     1,     0,     0,    -2,    -2,     0,     0,     0,    -1,    -1,     1,     2,     0,     0,    -2,     1,     2,     0,    -1,     2,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,    -2,    -2,     0,     0,     0,    -1,     0,    -1,     1,     1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     1,     1,     0,     2,     1,    -1,    -2,     0,     0,     0,    -1,     0,    -1,     0,     1,     0,    -1,     0,     0,     1,     0,     1,    -1,    -1,    -1,     0,     1,     0,     2,     1,     1,     1,     2,    -1,    -2,     0,     0,     0,    -1,     1,    -2,    -1,     1,     0,    -1,    -1,     0,     1,     1,     1,     1,     0,     0,    -1,     0,    -1,    -1,    -1,     1,     0,     1,     0,     0,     0,     0,     0,    -1,     1,    -1,    -1,     0,    -2,    -1,    -1,     0,    -1,     0,     2,     2,     0,     0,     1,     0,     0,    -1,     1,     1,     1,     2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,     0,    -1,    -2,    -2,     1,     1,     0,     0,     0,     0,     1,    -1,     1,     2,     1,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,     1,    -2,    -4,    -4,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     1,    -1,    -1,    -1,     0,    -1,    -3,    -2,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,     2,     0,    -3,    -2,    -2,    -3,    -3,    -3,    -3,    -1,    -1,    -2,    -2,    -2,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -2,    -2,    -3,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		     7 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -1,    -3,    -1,     0,     0,    -1,    -2,    -2,    -3,    -2,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     1,     2,     1,     2,     1,    -1,     0,     0,     1,     1,     1,     0,     0,    -1,    -2,    -3,    -2,    -2,    -3,    -4,    -3,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     0,     0,     1,     0,     2,     1,     1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -2,    -2,    -3,    -2,    -2,    -1,     0,     1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,     1,     0,    -1,    -2,    -1,    -1,    -2,    -1,     0,    -1,     0,     1,    -1,    -2,    -2,    -1,    -1,     2,     1,     0,     2,     2,     0,     1,     0,     1,     0,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -3,    -3,    -1,     0,     1,     0,     1,     1,     2,     1,     0,     2,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     0,     1,     1,     1,    -1,    -1,     0,     2,     3,     0,     0,     0,    -1,     1,     0,     1,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     1,     1,     1,     1,     0,     0,     0,     1,     1,     2,     0,    -1,     0,     1,     0,    -1,     2,     2,     2,     1,     0,     0,     0,     0,     0,     0,    -1,     1,    -1,     1,     1,    -1,    -1,    -1,    -1,    -2,     0,     2,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     2,     0,     1,     1,    -2,    -2,    -2,    -1,    -1,    -1,    -2,    -2,    -2,    -3,    -3,     0,     0,     0,     0,     1,     0,     1,    -1,     0,     2,     1,     1,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,    -3,    -3,    -2,    -2,    -3,    -2,     0,     0,     1,     0,     1,     1,     2,    -1,     0,     0,    -1,    -2,    -2,     0,     0,     0,    -1,     0,    -2,    -1,    -1,    -3,    -1,    -1,     0,     0,     0,     0,     1,     1,    -1,     1,     0,     0,     2,     0,     1,     0,    -1,    -3,    -1,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,    -2,     0,     1,     1,     1,     1,     1,     1,    -1,    -1,     0,     0,     0,     0,     1,     1,    -1,    -3,    -3,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -1,     0,     1,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -1,    -2,    -3,    -2,    -1,    -3,    -2,     0,     1,     2,    -2,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -1,     0,     1,     0,     0,    -1,    -3,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,     0,     0,    -1,    -2,     0,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -2,    -2,    -1,     0,     1,     0,    -1,     0,    -2,     0,     0,     0,     0,    -2,    -1,     1,     2,    -1,     0,     0,     0,    -1,     0,     0,    -3,    -2,    -3,    -3,    -2,    -2,    -2,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,    -3,     1,     1,     1,     2,     2,     1,     1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -2,    -2,    -2,     0,     0,    -3,    -2,     0,    -1,     0,     0,     0,    -1,    -3,     1,     0,     1,     3,     0,     0,     0,     1,    -1,    -1,    -2,    -1,    -2,    -4,    -3,    -3,    -2,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     1,     2,     1,     0,     2,     0,    -1,     0,     0,     1,    -1,    -1,    -3,    -3,    -3,    -2,    -2,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0,    -1,     1,    -1,     0,     0,     1,    -1,    -1,     0,     1,     0,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -3,     0,     0,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,     0,     1,     1,     1,    -1,     0,     0,     1,    -1,     0,     0,    -1,     0,     0,    -1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     1,     1,    -1,     2,     1,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0),
		     8 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,     0,    -1,    -1,     1,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,     1,     1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     2,     1,     0,    -1,     1,     2,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     1,     0,    -1,    -1,     1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     1,    -1,    -1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,    -2,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -2,    -2,     1,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,    -2,    -1,     0,     2,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -2,     1,     0,    -2,    -2,    -2,    -1,     0,     1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     2,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,     0,     0,     1,     1,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,     1,    -1,    -1,     0,    -2,     0,    -1,     0,     0,    -1,     0,     1,     1,     1,     0,     0,     1,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     1,     0,    -2,    -2,    -2,     0,     0,    -1,    -2,     0,     1,     0,    -2,     1,     2,     1,     1,     0,    -1,    -1,     0,     0,    -2,    -1,     0,     1,     2,     1,     1,     0,    -2,    -3,     0,     0,     0,     0,    -2,    -1,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -1,     1,     1,     1,     1,    -1,    -2,    -2,    -2,    -3,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     0,    -2,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,     1,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -2,    -1,     0,     0,    -1,     1,    -1,    -1,    -1,    -1,    -2,    -4,    -2,     0,     1,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0,    -1,     1,     1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -2,     1,     1,     0,     0,     1,     0,     0,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     2,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -2,    -1,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -3,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     1,     1,    -1,     1,     1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -3,     0,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		     9 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -1,     0,     1,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,     0,     0,     1,    -1,    -1,    -2,    -2,    -2,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     1,    -1,     0,    -2,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -3,    -3,    -3,    -2,    -1,    -1,    -1,    -2,     1,     0,     0,     0,     3,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -3,    -1,    -2,    -1,     0,    -2,    -1,     0,     1,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,    -1,     2,     0,    -1,    -1,    -1,     0,    -2,     0,     0,    -1,    -1,    -2,     0,     1,     0,     0,     0,     1,    -1,     0,     0,     0,     1,     1,    -2,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,    -1,     0,     0,     1,    -1,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -1,     0,     1,     3,    -1,    -2,     0,    -3,    -1,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,     0,     0,    -1,    -2,    -2,    -3,    -1,    -1,     1,     0,     1,     0,     2,     3,     0,    -2,     0,     0,     0,    -2,     1,    -1,    -1,     0,     1,     0,     1,    -1,    -2,    -1,    -2,    -1,    -1,    -2,     0,     0,     1,     0,     1,     1,     0,    -2,    -2,    -2,     0,     0,    -1,    -1,     1,    -1,     0,     0,     0,     1,     2,     0,     0,     0,    -1,     1,     2,     0,     0,     2,     1,     2,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     1,    -1,     0,    -1,     2,     2,     1,     0,     1,     1,     1,     1,     0,     0,     0,     1,     0,    -2,    -1,    -2,    -2,     0,     0,     0,     0,     0,    -2,    -1,     1,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     2,     0,     0,     0,     0,     1,     0,    -1,    -2,    -2,    -2,    -2,     0,     2,     0,     0,     0,    -1,    -1,     1,    -1,     0,     0,    -1,     0,     0,     1,    -1,     0,    -1,    -1,     0,     1,     0,     0,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     1,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -1,    -1,    -2,    -1,     1,     0,     0,     0,     0,    -1,     0,    -2,    -2,     0,     1,    -1,    -2,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     1,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -2,    -1,    -2,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -2,    -1,     0,     0,     0,     2,    -1,    -1,     0,     0,     1,    -1,    -2,    -1,    -3,    -2,     1,    -1,    -2,     0,     1,     1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,     0,     1,     0,    -1,     0,    -1,    -1,    -2,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,    -1,    -2,    -2,    -2,    -3,    -1,     1,     1,     1,     1,     0,    -1,    -2,    -1,    -1,     0,    -2,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,     0,     1,     1,     0,    -1,     0,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     1,     0,     0,     0,    -2,     0,    -1,    -1,     0,    -1,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     1,     0,     1,     0,     1,     0,    -1,    -1,     0,     1,     1,     0,     0,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     2,     1,     0,     1,     1,    -1,     0,     1,     2,     0,     1,     1,     1,     2,     2,     1,     1,     2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     1,     1,     1,     2,     1,     1,     1,     1,     0,     1,     1,     2,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    10 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,    -2,    -1,    -2,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -2,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,    -2,    -2,    -1,    -2,    -3,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -2,    -1,     0,    -2,    -1,    -2,    -1,     0,     0,    -1,     0,    -1,     0,    -2,    -1,     1,     0,    -2,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     1,     1,    -1,    -2,    -2,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     0,    -2,     0,    -1,    -1,    -3,    -2,    -1,     1,     3,    -2,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -2,     0,     1,     0,     1,     1,    -1,    -2,     0,    -1,    -1,    -3,    -1,    -2,     0,     0,     0,     2,     0,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,     1,     1,     1,     0,     1,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,     0,     0,     3,    -1,    -1,    -1,     0,     0,    -1,    -2,    -2,     0,     0,     0,     0,    -1,    -2,    -2,     0,     1,     1,     0,    -2,    -2,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,     1,     1,     0,    -1,    -3,     0,     0,     0,     1,     0,    -2,    -2,    -1,     0,     1,     1,     0,    -1,    -2,    -1,    -2,    -2,    -1,     0,     0,     1,     1,    -1,     2,     1,     1,     0,    -1,     1,     0,     0,     0,    -1,    -3,    -4,    -2,     0,     0,     1,     2,    -1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,    -2,     0,     1,    -1,     0,     1,     1,     0,     2,     1,     0,    -2,    -2,    -1,    -1,     1,     2,     2,    -1,     0,     1,     0,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     1,     0,     1,     1,     3,    -1,    -3,    -2,    -1,     0,     2,     0,     1,    -2,     0,     1,     0,     0,    -2,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     1,     1,    -2,    -3,     0,     1,     1,     1,     1,    -1,    -2,    -1,     0,    -1,    -1,    -2,     2,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -2,     0,     1,     1,    -1,     1,     0,    -2,    -1,    -1,    -1,    -1,    -1,     3,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     1,     0,    -1,    -2,    -1,     0,     2,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,    -1,    -1,    -1,    -2,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,    -1,     0,    -1,    -1,     0,    -2,    -1,     0,     0,     1,     0,    -1,     0,    -1,    -2,    -1,     0,     0,     1,     1,     1,     1,     0,    -2,    -1,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     2,     0,     1,     1,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,     0,     0,     0,     4,     1,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     1,     0,     0,     0,    -2,     0,     1,     1,    -1,    -2,     0,    -2,    -1,    -1,    -1,     0,     1,     2,     1,     0,     0,     0,    -1,    -2,    -3,    -1,    -1,    -1,     1,     2,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -2,    -1,     0,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     1,     1,    -2,    -2,    -2,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -1,     0,     1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,     0,    -1,    -2,    -3,    -4,    -4,    -4,    -3,    -2,    -2,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -1,    -1,    -2,    -1,    -2,    -1,    -1,     0,    -2,    -1,    -2,    -2,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    11 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -2,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     1,     1,     1,     0,     0,     0,     0,    -1,    -2,    -2,     0,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,     1,     1,     0,     1,     1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     1,     1,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     1,     1,     1,     0,     0,    -2,    -1,    -1,    -1,    -1,     0,    -3,    -3,    -2,     0,     1,     0,     0,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     2,     0,    -1,     0,    -2,     1,     1,     0,    -3,    -3,    -4,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,     0,     1,     0,    -2,    -3,    -3,    -2,    -1,     0,     1,     0,     0,     0,     0,     0,    -2,    -3,    -2,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -2,    -1,    -2,    -3,    -1,     0,     1,     0,     0,     1,     0,     0,     0,    -2,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -2,    -3,    -3,    -4,    -4,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -3,    -4,    -2,     0,     2,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -2,    -1,    -1,     2,     1,     1,     2,     0,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,     0,    -2,    -1,    -2,    -1,    -1,     1,     2,     0,     1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     0,     1,     1,    -1,    -3,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     1,     0,     0,     1,    -1,    -2,    -4,    -4,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -2,     0,     0,     2,     1,     1,     0,     0,     0,     0,     1,     0,    -1,    -4,    -4,    -3,     0,     0,     0,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,    -1,     0,     0,     0,    -1,     1,     1,     0,    -3,    -2,     0,     1,     1,     2,     2,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -1,     0,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     0,     1,     1,     2,     3,     2,     2,     0,    -3,    -1,     0,     0,     0,     0,    -1,    -3,    -2,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     1,     1,     0,     2,     1,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     0,    -1,     1,    -1,    -2,    -2,    -1,     1,    -1,    -2,    -1,    -1,     0,     1,     1,     2,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,     1,    -1,    -1,    -1,    -1,     0,     2,     1,     1,     0,     0,     1,     1,     0,     0,     0,     2,     0,     0,     0,     1,    -1,    -1,    -1,     0,    -1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     1,     1,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     2,     2,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -2,     0,     1,     0,    -1,     1,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -3,    -1,     1,    -1,     0,     1,     0,    -2,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    12 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,     0,    -1,     0,    -1,     0,     1,     2,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     2,     0,     0,     0,     1,     1,     2,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,     2,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     2,     1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     0,     2,    -2,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,    -1,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     1,    -1,    -1,     0,     1,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     1,     1,     2,     1,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     1,     2,     1,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,    -1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     2,     1,     1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,    -2,    -1,     0,     1,     1,     1,     1,     2,     2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,     1,    -1,     0,     1,     1,     1,     1,     1,     1,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     1,     1,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     2,     0,     1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     0,     1,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -3,    -3,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0),
		    13 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -3,    -4,    -3,    -3,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,     1,     1,    -1,    -1,     0,     0,    -1,     1,     0,    -1,    -1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,     2,     2,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     2,     0,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     0,     1,     0,    -3,     0,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     1,    -1,     2,    -1,     2,     1,     0,     1,     0,     1,     0,     1,     1,    -1,    -1,     0,     0,    -1,     0,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     2,     0,     0,     1,     0,     2,     1,     1,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,     0,    -1,    -3,    -2,    -1,    -1,     0,     0,    -1,     1,     1,     1,     0,     2,     2,     1,     1,     0,    -2,    -1,     0,     0,     1,     0,     0,     0,     1,     0,     0,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     1,     2,     2,     1,     1,     1,    -2,    -3,    -4,    -2,    -2,     0,     1,     1,     0,     2,     0,     0,     0,    -1,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     2,     1,    -1,    -2,    -3,    -5,    -3,    -1,    -1,     1,     2,     0,     0,    -1,    -1,     0,     0,     1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     2,     2,    -1,    -2,    -4,    -2,    -2,     0,     1,     1,     1,     1,     0,    -1,    -2,    -1,    -1,    -2,    -2,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -2,    -1,     0,     1,     0,     1,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     1,     0,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -2,     0,    -1,    -1,    -1,     1,     0,    -2,    -1,    -1,     0,     1,     0,     1,    -1,    -1,    -1,     0,     0,     1,     1,     2,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     1,    -1,     2,     0,    -1,     0,    -1,     0,     0,     1,     1,    -1,    -2,    -1,    -1,     1,     2,     0,     0,     1,     1,     1,     0,     0,     0,     0,    -1,     0,     2,     1,     1,     0,    -2,    -2,    -1,     0,     0,     1,     1,    -1,    -3,    -3,    -2,    -1,    -1,    -2,     0,     0,     1,     0,     0,     1,     0,     0,     0,    -1,     1,     1,     0,    -1,    -3,    -1,     0,     0,     0,     1,     2,     0,    -2,    -2,    -3,    -4,    -6,    -5,    -5,    -5,    -4,    -3,    -3,    -1,     2,     0,     1,     1,     1,     2,     1,    -1,    -2,    -1,    -1,     0,     0,    -2,     1,     1,     1,    -1,    -1,    -2,    -3,    -4,    -4,    -4,    -3,    -3,    -3,    -2,    -1,     0,     1,     1,     1,     1,     2,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -2,    -2,     0,     0,     1,     1,     0,     0,     3,     0,    -1,     0,     0,     0,     0,     1,     1,     1,     0,     1,     1,     0,     0,     0,     0,     1,     1,    -1,     0,    -1,     0,     1,     0,     1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     2,     1,     0,     1,     1,     1,     0,    -1,     0,     1,    -1,     0,     0,    -1,     0,     0,     1,     1,     0,     1,    -2,    -2,     0,     0,     0,     0,     1,     2,     2,     0,     0,     1,     1,     0,     0,     1,    -1,     1,    -1,     0,    -1,    -1,    -2,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     2,     1,     0,     2,     1,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     1,     1,     1,     0,    -1,    -1,    -1,    -2,    -1,     0,    -2,    -2,    -2,    -1,    -1,    -1,    -3,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,    -2,     1,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0),
		    14 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -3,    -2,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -3,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     1,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -3,    -2,    -1,     0,     0,    -1,    -2,    -2,    -1,     0,     1,     0,    -2,    -2,     0,     1,     1,     1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     1,     1,     0,    -2,    -2,     0,     0,     0,    -1,    -1,     1,     0,     1,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     1,     0,     1,     1,     0,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,     1,    -2,     0,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,    -1,     0,    -1,     1,     1,     1,     3,     3,     2,     1,     1,     0,     1,    -1,     0,     0,    -1,     0,    -1,     0,    -2,    -1,     0,     0,     1,     1,     1,     0,     0,     1,     0,     1,     1,     1,     2,     2,     2,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -3,     0,     0,     0,     0,     2,     1,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -2,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,     1,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -3,    -3,    -2,    -2,    -1,     0,     0,    -1,     1,     0,    -2,    -2,    -2,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,     0,    -1,     0,     0,     1,     0,     1,    -1,    -3,    -3,    -2,    -1,    -2,     0,     0,     0,     1,    -1,     0,     1,     0,     1,     1,     1,     0,     1,     1,    -1,     1,     1,     0,     0,     0,     1,     2,     1,    -1,    -2,    -1,    -2,    -2,     0,     0,    -1,     0,     1,     0,     0,     0,     1,     1,     0,     1,     1,     0,     0,     2,     1,     1,     1,     1,     1,     1,     0,     0,    -2,    -1,    -2,     0,     0,     0,    -3,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     2,     0,     1,     2,     1,     1,     0,     0,    -1,     0,    -1,     1,     0,     0,     0,     1,     0,     1,    -2,    -1,     0,     0,    -1,    -2,    -1,    -1,     1,     1,     2,     2,     2,     2,     0,     0,     0,     1,    -1,    -1,    -1,     2,    -1,     0,     0,     0,     1,     1,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,     2,     3,     2,     3,     1,     2,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     1,    -1,     2,    -1,    -1,    -1,     0,    -1,     0,     1,     2,     2,     2,     2,     3,     1,     1,    -1,    -1,     0,     0,     0,    -1,     0,     1,    -1,    -2,     0,     0,     0,     2,    -1,    -1,    -1,    -3,    -1,     0,     1,     1,     0,     2,     2,     2,     1,     0,    -1,     0,     0,     0,     2,    -1,    -2,    -1,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     1,     1,     2,     0,    -1,     1,     1,     0,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,     0,     1,     1,     1,     1,     1,     1,     0,     0,     2,     0,     1,     1,     1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -2,    -1,    -2,     0,    -2,     0,     1,     0,     0,    -1,    -2,    -2,     2,     1,     1,     0,     0,     1,     0,     0,     1,     0,    -1,    -3,    -2,     0,     0,     0,     0,    -1,    -4,    -2,     0,     0,     0,    -2,     0,    -1,    -1,     0,     0,     1,     0,    -1,    -1,     1,     0,     1,     0,     1,    -1,    -2,    -1,    -1,     0,     0,     0,    -2,    -4,    -3,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -3,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     2,    -1,    -1,     0,     0,    -2,     1,    -1,     0,     0,     0,     0,     0,     2,     1,    -1,    -2,    -1,     0,    -2,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,     1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     2,     0,    -1,    -2,    -1,    -1,    -2,    -1,    -3,    -2,    -2,    -3,    -2,    -2,    -2,    -1,    -3,    -4,    -4,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -2,     0,    -1,    -2,    -1,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     0),
		    15 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -2,    -2,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     1,     1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     1,    -1,    -1,     0,     0,    -1,    -2,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     1,     1,     0,    -1,    -1,    -1,     0,    -1,     0,     1,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,     0,    -1,    -2,    -2,    -3,    -3,    -3,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     1,     0,     0,    -2,    -1,     1,    -1,     0,     0,    -1,    -3,    -1,    -1,    -3,    -2,    -1,    -1,    -1,     0,     0,    -1,    -2,     0,     0,     0,     0,    -1,    -1,     1,    -1,    -2,    -1,     0,     0,     0,     0,    -2,    -1,    -2,     1,     1,     1,    -1,    -1,     0,    -1,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     1,     0,     0,     1,     1,     2,     2,     1,     1,     1,     3,     2,     2,     1,     0,     0,     0,     0,     0,    -1,    -1,     1,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     1,     0,     1,     1,     2,     2,     3,     3,     1,     1,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     2,     1,     2,     1,     0,     1,     3,     0,     0,     0,     0,     0,    -2,     0,    -1,    -1,     1,     0,     1,     0,     0,     0,    -1,    -2,     0,     0,    -3,    -2,    -1,    -2,     0,    -1,     0,     0,     2,    -1,     0,     0,    -1,    -2,     1,     1,     0,     0,     1,     0,     1,     2,     1,     1,    -2,    -2,    -2,    -2,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     2,     0,     0,     0,     0,     1,     0,     0,     2,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -2,     0,    -1,     0,    -1,    -1,     0,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,    -2,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,    -3,    -2,     0,    -2,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,     1,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,     1,     1,    -1,    -1,    -2,     1,     1,     0,    -1,     0,    -1,    -1,     1,    -1,    -1,    -1,    -1,     0,     0,     1,    -1,     0,    -1,     1,     1,    -1,    -1,     0,     0,     0,     0,     1,     0,     1,     0,     1,     0,     0,    -1,     0,     1,     0,    -2,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,     1,     1,     0,     1,     1,    -1,     0,     0,    -1,     0,     1,     1,     0,     0,    -1,     0,     1,     0,     0,     0,    -2,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     0,    -1,    -1,     1,    -1,     0,     0,     0,     1,     0,     1,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     1,     1,     1,     0,     1,     1,     0,     1,     0,     1,     1,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,     0,     0,     1,     0,     1,     0,     1,     2,     1,    -1,     0,     0,    -1,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     1,     1,     1,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,     0,    -1,     0,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0),
		    16 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,     1,     0,    -1,     0,    -1,    -1,     1,     0,     2,     2,     0,    -1,    -1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     1,     2,     1,     0,     0,     2,     1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     2,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     1,     1,     0,     0,    -1,     0,     2,     2,     0,     0,     0,     0,    -2,    -3,    -1,    -2,     0,     0,     1,     1,     0,     0,    -2,    -2,     0,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,     1,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     1,     0,    -1,     1,     1,     0,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     1,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,    -2,    -1,    -2,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     1,     1,     0,     0,    -1,    -1,    -2,    -3,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     1,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     1,     1,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     2,     0,    -1,    -1,     0,     0,    -1,     1,     0,     0,    -2,    -1,    -1,    -3,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     2,     2,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     1,     1,     0,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     1,     1,     0,    -1,    -1,     0,     0,     0,    -1,     1,     1,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,    -2,     0,     0,     0,     0,    -1,     0,     1,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -2,     0,     0,     0,     1,     0,     1,     1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,     2,     1,    -1,     0,    -1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     1,     2,     1,    -2,    -2,    -1,     0,    -1,     0,     1,     0,    -1,    -1,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,    -2,    -1,     0,     1,     0,     1,    -2,    -1,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     2,     1,     1,     0,    -1,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,     1,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -2,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     2,     1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    17 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -2,    -2,    -1,    -2,    -3,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,    -2,    -2,    -4,    -5,    -5,    -4,    -3,     0,    -2,    -1,    -1,     0,     0,     0,     0,     1,     2,     0,     0,     0,    -1,    -1,    -1,    -2,     1,     1,     1,    -1,    -3,    -2,     0,     0,     0,    -1,     2,     1,     0,    -1,    -1,    -2,    -1,     0,     3,     3,     2,     0,     0,     0,     1,     0,     0,     0,    -1,     1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,     0,    -2,    -1,    -2,     3,     1,     0,    -1,    -1,    -1,     0,    -1,     0,     1,     0,     1,    -1,    -1,    -1,    -1,     1,     1,     0,     0,    -1,     0,     1,     2,     1,    -1,    -1,     0,     2,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,     0,     1,     0,    -1,     0,     1,     1,     0,     0,     0,     1,     2,     0,    -2,     0,     0,     1,     1,     0,     1,     0,     1,     0,     1,     0,     0,     1,     1,     2,     0,    -1,    -1,     0,     0,     1,     1,     1,    -1,    -1,    -1,    -1,    -2,     1,     0,     0,     1,     1,     1,     2,     0,    -1,    -1,     1,     0,     2,     2,     0,    -2,    -1,    -1,     0,     2,     1,     1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     1,     1,     0,     1,     0,     1,     1,     1,     1,     1,     1,    -4,    -4,    -1,     1,     1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,     1,     1,     0,     0,     1,     1,     1,     1,     0,     0,     0,    -1,    -5,    -4,    -2,     1,     0,     1,    -1,     0,     1,    -1,    -2,     0,    -2,     0,     0,     0,     1,     3,     1,    -1,     2,     0,     0,     0,     1,     2,     0,    -2,    -7,    -3,    -1,     1,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,    -2,     1,     1,     1,    -1,    -1,     2,    -1,    -6,    -4,    -2,    -1,     1,     1,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     2,     0,     0,     2,    -3,    -6,    -1,     0,     0,     0,     0,     1,     1,    -1,     0,     1,    -1,    -1,    -1,     0,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -2,    -3,    -4,    -3,     0,     0,     0,     0,    -1,     1,    -1,     0,     0,     1,    -3,    -4,    -1,     0,    -1,     1,     0,     2,    -3,    -1,     0,     1,     0,    -1,    -3,    -5,    -1,     0,     1,     1,     0,     1,     1,     1,    -1,     1,    -1,    -1,    -4,    -4,     0,     0,     0,     0,     1,     1,    -2,     0,     0,     0,    -3,    -3,    -4,    -4,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,    -2,    -2,    -3,    -2,     1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -4,    -1,     1,     1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,    -2,    -2,    -3,    -1,     0,     0,     0,     0,     0,     0,    -1,    -3,    -1,    -3,    -2,    -2,    -1,     2,     1,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,     0,    -1,     0,     0,     4,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,    -1,     1,     1,     1,     1,     0,     1,    -2,     0,     1,     0,     0,    -1,    -1,     1,    -1,    -1,     0,    -3,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -2,     1,     0,     0,     1,     0,     0,     1,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -2,    -2,     0,    -2,     0,     0,     0,     0,     0,     0,    -2,    -3,    -1,    -1,     0,     0,     0,     0,     1,     0,     1,     0,     1,     1,    -1,     0,    -1,     1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,     0,     1,     1,     0,     1,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     1,     1,     0,     1,     0,     0,     0,     0,    -1,    -1,     1,     1,    -1,     1,     2,     1,     1,     0,     0,     0,     0),
		    18 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -3,     0,     0,     0,    -1,    -1,    -2,    -3,     0,     0,     0,     1,     1,     2,     2,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,    -2,    -1,    -2,     0,     0,    -1,    -2,     0,    -1,    -2,    -2,     1,     0,     0,     0,     0,     1,     2,     2,     1,     1,     0,     2,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     2,     1,     0,     2,     2,     1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     1,     0,     0,    -1,     1,     0,     0,     0,    -1,    -2,    -1,     1,     0,    -1,    -2,     1,     0,     3,     0,    -1,     0,    -2,    -1,     0,     0,    -1,     1,     2,     0,    -1,    -1,     0,     0,     0,     0,     1,    -1,     0,     1,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,    -1,     1,     2,    -1,     1,     1,    -1,     1,     0,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,    -2,     0,     1,     1,     0,     0,     1,     1,     0,     0,     0,     0,     1,     1,    -1,    -1,     0,    -1,    -1,     1,     1,     0,     0,    -1,    -2,     0,     0,    -1,     1,     1,     0,     0,     1,     0,     0,    -1,    -3,     0,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     1,     0,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     0,    -1,     0,     1,     0,    -2,    -1,    -3,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     1,     0,     1,     1,     0,     0,    -1,     0,    -1,     0,    -2,    -1,    -2,    -1,     1,     2,     0,     2,    -2,     0,     0,    -1,     2,    -1,     1,     0,     0,    -1,    -1,     0,    -1,     1,     1,     0,    -1,    -1,     0,     0,     1,    -1,     0,     1,     3,     3,     1,     1,    -3,     0,     0,    -1,     1,     0,    -1,    -3,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,    -2,     0,     0,     1,     1,     2,     3,     3,     1,    -1,    -1,     0,     0,     0,     0,    -2,     0,    -2,    -1,    -1,    -2,    -2,     0,    -1,     0,     1,     0,     0,    -2,     1,    -1,     1,     0,     1,     0,     2,     1,    -1,    -2,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -2,    -1,     0,     1,     0,     0,    -1,     1,    -3,    -1,     0,    -1,    -2,     0,     2,     2,     0,    -2,    -1,     0,     0,    -1,     1,    -2,     1,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -1,     0,    -2,    -2,    -2,    -1,     1,     0,     1,    -2,    -1,     0,     0,    -1,     1,    -2,     0,     0,     1,    -1,    -1,     0,     1,     1,    -1,     1,     1,     0,     0,    -2,    -2,    -1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,     1,     1,     2,    -1,    -3,    -1,     1,     0,     0,    -1,     1,    -1,    -3,    -1,     0,    -2,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,    -1,    -2,     1,     0,     1,     1,    -1,    -3,    -1,     0,     0,     1,    -1,     0,    -1,    -2,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -3,     0,    -1,     1,     1,     1,     1,     2,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -2,    -3,     0,     1,     1,     1,     0,     0,     0,    -1,    -1,     1,    -1,    -1,     0,    -1,    -3,    -2,     0,    -1,     0,     1,    -2,     0,     0,     0,     0,    -1,    -2,    -3,    -2,     0,     0,     0,     0,     1,     0,     1,    -1,     0,    -3,     0,     0,    -2,    -4,    -2,    -1,    -1,     0,     1,    -2,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,    -1,    -2,     0,     1,     0,     1,    -1,     0,     1,    -2,    -4,    -3,    -1,    -2,    -1,     1,     1,    -2,     0,     0,     0,     0,     0,    -2,    -3,    -2,     0,     1,     0,     0,     0,     1,     1,     1,     0,     1,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -1,    -2,    -2,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -1,     1,    -2,    -2,    -1,     0,     1,    -1,     0,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,    -1,    -2,    -2,    -1,    -2,    -3,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    19 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     2,     1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -3,    -3,    -2,    -2,    -3,    -2,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -3,    -3,    -4,    -4,    -3,    -3,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,    -1,     1,     0,    -1,    -1,    -1,    -2,    -2,    -4,    -4,    -2,     0,     0,     0,     1,     1,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -3,    -4,    -2,    -1,     1,     1,     2,     2,    -1,     1,     0,     1,    -1,    -1,     1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     2,    -1,     0,    -1,    -2,    -1,     1,     1,    -1,    -1,     0,     0,     0,     1,    -2,     0,     1,     1,    -2,    -2,    -1,     0,     0,    -1,     1,     1,     1,     0,     0,    -1,    -2,    -1,     0,     1,     1,     0,    -2,     0,    -2,    -3,    -1,     0,    -1,    -1,     2,    -1,    -1,    -2,     0,    -1,     0,    -1,    -2,     1,     1,     0,    -1,    -2,    -1,     1,     1,     1,     0,     0,     0,     0,    -1,    -2,     0,     0,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,    -1,     1,     0,     0,     0,     3,     2,     1,     0,     0,    -2,    -3,    -1,    -2,    -1,    -1,    -2,    -2,    -2,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     1,     2,     1,     1,     1,     1,     0,     0,     0,    -4,    -4,    -1,    -2,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     1,     0,     0,     1,     1,     1,     2,     1,     1,    -4,    -3,    -1,    -1,     1,     1,     0,     2,     0,     0,     0,    -1,     0,     0,    -3,    -2,    -1,     0,     0,     2,     1,     1,    -1,    -1,     0,     0,     0,    -4,    -5,    -2,     1,     0,     0,     2,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -1,    -1,    -1,     1,     0,    -1,     0,     1,     0,    -1,    -1,    -2,    -2,     1,     2,    -1,    -1,     2,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -3,    -3,    -1,     0,    -1,    -2,     0,     1,     1,    -2,    -1,    -2,    -2,     1,     1,     0,     0,     0,     0,    -2,    -1,     0,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -4,    -3,    -2,    -2,     0,     0,     0,     0,    -2,    -1,    -2,     0,     1,     2,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -3,    -2,    -1,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,    -2,     1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -1,     1,     1,     0,     0,     1,    -2,     1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     1,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     1,     2,     0,    -1,     1,     2,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -2,    -1,     1,     2,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,     0,     1,     0,     0,     1,     0,    -2,    -1,     1,    -1,     1,    -1,    -1,     3,     1,    -1,    -1,     0,     1,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     2,     2,     0,     0,     1,     0,     1,    -1,     1,     2,     1,     2,     0,     3,     3,     0,    -2,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     2,     2,     1,     1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    20 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     1,     0,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     1,     2,     1,     2,     1,     0,     0,    -2,    -1,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     1,     1,     1,     1,     1,     1,     1,     0,     0,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,     1,     0,     0,     1,     0,     1,     1,     0,     1,     0,     0,     1,    -1,     0,     1,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -2,     0,     0,     0,     1,     0,    -1,    -2,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,    -1,     0,    -1,     0,     1,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,    -2,     1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,    -2,     1,     0,    -1,     0,     0,    -1,    -2,    -2,    -1,    -3,    -3,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,    -2,    -1,     0,     0,    -1,     0,     1,     0,    -1,    -1,     0,    -2,    -2,    -2,    -2,    -3,    -2,     0,     0,     1,     0,     0,     1,    -1,    -1,     0,     1,     1,    -2,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     1,     0,     1,     0,    -1,     0,     1,     0,     0,    -2,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,    -1,     0,     1,     0,    -1,    -2,    -1,     0,     1,     1,     0,     1,    -2,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     1,     1,     0,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -1,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0),
		    21 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     2,     1,     0,    -1,     0,     1,     1,     1,     0,    -2,    -1,     2,     0,    -2,    -1,    -1,    -1,    -1,     0,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     0,     2,     2,     0,    -1,     0,     2,     2,     2,     1,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     2,     0,     1,     1,     1,     2,     1,     1,     2,     2,     1,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     1,     0,    -4,    -2,    -2,     0,     0,    -1,     0,     1,     0,     1,     2,     1,     1,     3,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,    -2,    -2,    -1,     0,    -2,    -2,    -2,    -3,     1,     2,     3,    -1,    -1,     1,     0,     1,    -1,     1,     0,     1,     0,    -1,    -1,     1,    -1,     1,     1,     0,    -1,    -3,    -2,     0,    -2,    -2,    -3,    -3,     0,     2,     2,    -1,    -2,     1,    -1,     0,     1,     1,     1,     0,     1,     1,     0,     0,     0,     1,     0,    -2,    -1,    -4,    -1,     0,    -1,    -2,    -3,    -2,    -1,     0,     1,    -1,    -1,    -1,    -2,    -1,     2,     0,     0,     0,     1,     2,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -2,     0,    -1,    -2,    -3,    -2,    -1,    -1,     0,     1,    -1,    -1,    -2,     0,     1,     0,     0,     2,     2,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -2,     0,     0,     0,    -1,    -2,     0,     0,    -1,     2,     1,     0,    -1,    -1,     0,     0,     0,     0,     2,     3,     1,     0,     1,    -2,    -2,    -2,    -2,    -2,    -2,     2,     0,     0,    -3,    -1,     0,     0,     1,     2,     0,    -1,    -1,     0,     1,     0,     1,     1,     1,     2,     1,     0,     0,    -2,    -2,    -1,    -2,    -1,     0,     2,     0,     0,    -1,     0,    -1,     1,     1,     1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     2,    -1,     0,     0,    -1,    -1,    -3,    -2,     1,     1,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,     0,    -3,    -1,     0,    -1,    -1,    -1,    -2,     1,     3,     0,     0,     0,     0,    -1,    -2,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,    -1,    -2,    -3,    -2,    -1,     0,    -2,    -2,    -3,    -1,     0,    -1,     0,     0,     0,    -2,    -2,     0,     0,    -1,    -1,     1,     0,    -1,     0,     1,     1,    -2,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,    -3,    -1,     1,     0,    -1,    -1,    -2,    -1,     1,     1,     1,     1,    -2,    -2,    -3,    -2,     0,     0,     1,     2,     2,     1,     0,    -1,    -2,     0,     0,    -1,    -3,    -2,    -2,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     2,     2,     2,     2,     0,     0,     1,     1,    -1,     1,     0,     0,     0,    -3,    -2,    -1,     0,     0,     0,     0,     1,     1,    -1,    -1,     1,     0,    -1,     0,     0,     1,     3,     2,     0,     1,     2,     1,    -1,     0,     0,     0,    -1,    -3,     0,     0,     1,     0,     1,     1,     2,     1,     0,    -1,    -1,     0,     0,     1,     2,     2,     3,     1,     0,     0,     1,     0,     0,     0,     1,     0,    -2,     0,     0,     1,     0,     0,     0,     1,     1,    -1,    -2,    -1,    -1,     1,     1,     0,     2,     2,     3,     2,     0,    -1,     1,     1,    -1,     0,     0,     0,    -2,    -1,    -1,     1,     0,     0,     1,     0,     1,    -1,    -1,     0,    -1,     1,     0,     1,     4,     3,     2,     2,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -2,     0,    -1,     0,     2,     0,     1,     3,     1,     1,     2,     1,     2,     1,     0,    -1,    -2,    -1,     1,     0,     0,     0,     0,     0,    -2,    -1,    -2,     0,    -2,    -2,     0,    -1,     0,     0,     0,     1,     1,     2,     1,     1,     0,     1,     1,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -3,    -3,    -2,    -5,    -4,    -4,     0,     0,    -1,     0,    -2,    -3,    -3,    -4,    -3,    -3,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -4,    -4,    -3,    -5,    -5,    -3,    -2,    -2,    -3,     0,     0,     1,    -2,    -1,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    22 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,    -3,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     1,     1,     2,     1,     1,     1,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -2,    -2,     1,     1,    -1,     0,     3,     1,     2,     2,     1,     0,    -1,     0,     0,    -2,    -1,    -1,     1,     0,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     1,     1,     1,     2,     1,     1,     1,     1,     0,     0,     1,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     1,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,     1,     2,     1,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,     1,     0,     0,     0,     1,     0,     1,     2,     1,     0,     0,     0,    -2,    -1,    -1,    -2,    -3,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,     1,     1,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -1,    -3,    -1,     0,    -1,     0,    -1,     1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,     0,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,    -2,    -2,    -2,    -2,    -1,    -2,    -2,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -3,    -2,    -2,    -1,     1,     1,     1,     0,    -1,    -3,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -4,    -3,    -3,    -3,    -3,    -3,    -2,    -2,    -3,    -1,     0,    -1,     1,     0,    -1,    -1,     1,     1,     0,    -2,    -1,     0,    -1,    -1,    -1,    -3,    -2,    -2,    -4,    -3,    -2,    -2,    -3,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -2,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,     0,    -1,    -1,    -1,     1,     2,     2,     1,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,     1,     0,    -1,     0,     1,     1,     2,     2,     2,     3,     0,     1,     1,     1,     0,     1,     0,     0,    -1,     0,     0,     1,     0,     1,     1,     0,    -1,     0,     1,     1,     2,     1,     0,     1,     2,     2,     1,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     1,     2,     0,     0,     1,     0,     2,     1,     1,     1,     0,     0,     0,     1,     0,     0,     0,     0,     1,     1,     1,     1,     1,     2,     1,     0,    -1,     2,     2,     1,     0,     0,     1,    -1,     1,     1,     1,     0,     1,     0,     1,    -1,     0,    -1,     0,     1,     0,     1,     1,     0,     0,    -1,     0,    -1,    -2,     1,     0,     1,     0,     0,    -1,    -2,    -1,     2,     1,     1,     2,     1,     0,    -1,    -2,     0,     0,     0,     1,     0,    -1,     0,     1,    -1,     1,     0,     1,     0,     0,     3,     0,    -1,     0,    -3,    -1,    -2,     0,     0,     1,     0,     0,    -2,    -2,    -1,     0,     2,     0,     1,     0,    -1,     0,     0,     1,    -1,     0,    -1,     2,     2,     0,    -1,     1,     0,     0,     0,    -2,     0,     2,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,     1,    -1,     0,    -1,    -1,    -1,     1,    -1,     1,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -1,     1,     0,     0,    -2,    -1,    -3,     0,     0,     0,     1,     2,     1,     0,     0,    -1,    -1,     0,    -1,     0,    -2,    -1,    -3,    -4,    -1,    -2,     0,     0,    -1,    -1,     1,     0,     0,    -2,    -3,     0,     0,     0,     0,     1,     0,     0,    -2,    -1,    -1,     0,     0,    -1,    -1,    -3,    -2,    -3,    -2,    -2,    -1,    -3,    -2,    -2,     0,    -1,    -1,    -2,    -3,     0,     0,     0,    -2,    -1,    -2,    -1,    -4,    -2,    -2,    -3,    -3,    -2,    -3,    -4,    -4,    -3,    -2,    -1,    -4,    -4,    -3,    -1,     0,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -2,    -2,    -2,    -3,    -3,    -2,    -3,    -2,    -1,    -1,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0),
		    23 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -1,    -1,    -2,    -3,    -2,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     3,     1,     1,    -1,     0,     0,     0,    -1,     0,     1,     0,    -3,    -2,    -1,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,     1,     0,     0,     1,     1,     0,     1,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -3,    -1,    -2,    -3,    -2,     0,     0,     0,     0,     0,     1,     0,     0,     1,     1,     0,     0,     0,     1,     1,     0,     1,     0,     0,     1,    -1,    -1,    -1,    -3,    -3,    -3,    -3,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,     2,     2,     0,     1,     2,     2,     0,     0,     1,     0,     1,     0,     0,     1,     0,    -1,    -3,    -3,    -3,    -1,    -1,    -1,     0,     0,     0,     0,     1,     2,     2,     1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     1,     1,     0,     0,    -2,    -3,    -3,    -3,    -2,     0,    -1,    -1,    -1,     0,     0,     1,     0,     2,     1,     1,     0,    -2,    -1,    -4,    -2,    -1,    -1,     1,     1,     0,     0,     1,    -2,    -2,    -3,    -3,    -2,    -1,    -2,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -5,    -4,    -3,    -3,    -1,     0,     1,     1,     1,     0,     0,    -2,    -4,    -3,    -3,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -2,    -3,    -5,    -6,    -3,    -1,     1,     0,     0,     1,     1,     0,     0,     1,    -2,    -3,    -4,    -3,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -3,    -3,    -3,    -2,     2,     1,     1,     2,     1,     2,     1,     0,    -2,    -2,    -1,    -2,    -2,    -2,    -1,     0,    -2,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     2,     1,     2,     1,     0,     0,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,     1,     1,     3,     2,     1,     0,    -1,     0,     0,     2,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     1,     0,     1,     0,     1,     0,    -3,     0,    -1,     0,     1,     0,    -1,     0,     0,    -1,    -2,    -1,    -2,    -1,    -2,    -1,     0,     0,    -2,     0,     1,     0,     0,     0,     2,     0,     1,     1,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -1,    -2,    -2,    -3,    -5,    -3,    -1,    -1,     0,     1,     0,     1,     0,     2,     2,     1,     1,    -3,    -3,    -1,     0,     1,     1,     1,    -1,    -1,    -1,     0,     2,     0,    -1,    -3,    -4,    -3,    -3,    -1,     0,     1,    -1,    -1,     0,     0,     1,    -1,    -1,    -3,    -1,    -1,     0,     1,     0,     2,     1,     1,     2,    -1,     2,     0,    -1,     0,    -1,    -1,    -1,    -1,     1,    -1,    -1,     0,     0,     0,     0,    -2,    -1,    -2,    -1,    -1,     0,     0,    -2,     0,     1,     1,    -1,    -1,     1,     0,    -1,     1,     2,     1,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -2,    -1,     0,     0,    -1,     1,    -1,     0,     1,     0,     1,     1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -2,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     1,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     2,     1,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,    -1,     0,     0,     0,     0,     1,     3,     3,     1,     0,     1,     0,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,     1,    -1,    -1,    -1,     1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     2,     1,     0,    -1,    -1,    -3,    -1,    -1,    -1,     1,     0,     0,     1,     0,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0),
		    24 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -3,     0,     1,    -1,    -2,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -3,    -3,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -3,    -1,     0,    -2,    -2,    -2,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,    -1,    -2,    -2,    -3,     0,    -2,    -3,    -2,     0,     0,     1,     1,     1,     0,    -1,     0,     1,     1,     1,    -1,     0,     0,     0,     0,     0,    -1,     1,    -2,     0,    -1,    -1,     0,     0,     0,    -1,     1,    -1,     0,     1,     0,    -1,    -2,     1,     1,     2,     3,     1,     0,    -1,     0,     0,     0,    -1,     1,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,    -1,    -2,    -1,     1,     1,    -1,    -1,     0,    -1,    -1,    -5,    -6,    -2,     0,     1,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -3,    -5,    -5,    -1,     1,     1,     1,     3,     2,    -1,    -2,     1,    -1,    -1,    -1,     1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     1,    -1,    -3,    -5,    -4,    -1,     1,     0,     0,     1,     1,    -1,     0,     1,    -1,     0,    -1,     1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -4,    -5,    -3,    -1,     2,     1,     0,     1,     1,     0,     0,    -1,     0,     0,     0,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     1,     0,    -3,    -4,    -3,    -2,     2,     2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,    -1,    -1,    -3,    -2,     0,     0,     2,    -1,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1,    -3,    -2,    -2,     0,     2,     1,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     1,     1,     0,    -2,     0,    -1,     0,     0,     0,    -1,     2,     0,     2,     0,     1,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,     3,     2,     0,     1,    -1,     0,     0,     2,     1,     0,    -1,     0,    -1,    -1,    -1,     1,     0,     0,     0,    -1,     1,    -1,    -3,    -2,    -1,     0,     0,     0,     1,     0,    -2,     0,     1,     1,     2,     1,     3,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,    -2,    -2,    -1,     1,     2,     2,     1,     2,     1,    -1,     0,     0,     0,     0,     0,     2,     1,     1,     1,     1,     0,    -2,    -1,     1,    -1,     0,     0,     0,    -3,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     1,     1,     1,     1,     1,     1,     1,     1,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -2,     0,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     1,     1,     0,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -2,    -2,    -2,     0,    -1,     0,     0,    -1,     0,    -1,     1,     1,    -1,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,    -2,    -1,    -1,    -1,    -1,    -2,    -4,    -3,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,    -1,     1,     1,     0,    -2,    -1,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -2,    -3,    -2,    -3,     1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,    -2,    -1,    -2,     0,     1,     1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,    -1,    -1,     0,     0,    -2,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     0,    -3,    -2,    -1,    -1,    -2,     0,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -2,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0),
		    25 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,     1,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     1,     1,    -1,     1,     1,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -3,    -2,    -2,     0,     1,    -1,     1,     1,     0,    -1,     0,    -1,     1,     1,     1,     0,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     1,     2,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -4,     0,    -1,     1,     0,     0,    -1,     0,     1,     0,     0,     1,     1,     2,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -3,     0,    -3,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     1,     1,     1,     2,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     1,     1,     2,     2,     2,     0,     1,     0,     0,    -1,    -1,     0,     1,    -1,    -1,     0,     0,     1,     0,     1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     2,     3,     2,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,     1,    -1,     1,     1,     2,     0,    -1,    -1,     1,     1,     1,    -1,     0,     1,     2,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,     0,    -2,    -1,     0,     0,     0,     0,     2,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     1,    -1,    -2,    -4,    -4,    -4,    -4,    -4,    -4,    -3,    -1,    -1,     0,     1,    -2,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     1,    -1,     0,     0,     0,    -2,    -3,    -3,    -4,    -3,    -4,    -4,    -4,    -2,     0,     0,     1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     1,    -1,     0,     0,    -1,    -1,    -2,    -3,    -4,    -3,    -3,    -2,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,    -2,    -3,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     1,    -1,    -1,    -2,    -3,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,    -3,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,     0,    -2,     2,     1,    -1,    -2,    -2,    -1,    -2,    -2,     0,     1,     0,     0,     0,     1,     1,    -1,    -2,    -3,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     2,     2,     1,     0,     0,    -2,    -2,    -2,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -3,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     2,     1,     2,     2,     0,    -1,     0,    -1,    -1,     1,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     2,     1,     0,     0,     0,     0,     1,     0,     0,     1,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     1,     1,     0,     1,     1,     0,     1,     1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,     0,     1,     0,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     1,     0,     0,     2,     2,     2,     1,     2,     1,     0,     1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     0,     2,     1,     1,     1,     1,     0,    -1,    -1,     1,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     1,     0,    -1,    -1,     0,    -2,    -1,    -1,    -1,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     1,     1,     1,     1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0),
		    26 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     3,     2,     0,     1,    -1,     0,    -1,     0,     1,     1,     3,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     1,     2,     3,     2,     1,     1,    -2,    -1,     0,     0,     0,     1,     1,     0,     1,     1,     2,     1,     0,    -1,     0,     0,     0,     0,    -3,    -1,     0,     2,     2,     1,     0,     0,     0,    -2,    -2,     0,     1,     1,     0,     1,     1,     1,     0,    -1,     0,     2,     1,    -2,    -1,     0,     0,     0,    -2,     0,     0,     2,     0,    -1,     1,     2,    -1,    -1,    -4,    -1,     0,    -1,     1,     0,    -1,     0,    -1,     1,     1,     2,     0,    -2,     1,     2,     0,     0,    -2,    -2,     1,    -1,    -2,     1,     1,     0,    -1,    -3,    -1,    -1,     0,     0,    -2,     0,    -2,    -1,     0,     0,     0,     1,     0,    -1,     3,     2,     0,     0,     1,    -1,     0,    -1,    -2,     1,    -1,    -2,    -1,    -2,     0,    -2,    -2,     0,    -1,     0,     0,     0,     0,    -1,     1,     0,     1,    -1,     1,     1,     0,     0,     0,    -1,     1,     0,    -1,     0,    -1,    -2,    -2,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     0,     0,    -1,    -1,     1,    -1,    -2,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -3,     0,    -2,     0,    -1,    -1,     1,    -3,    -1,    -2,     0,     0,    -1,     1,     0,    -2,    -1,    -2,    -2,     0,     0,     0,    -1,    -1,     0,    -2,    -3,    -3,    -3,    -2,    -2,    -2,    -5,    -2,     0,     0,    -1,    -2,     0,     0,    -2,    -2,    -1,    -2,    -3,    -3,    -2,     1,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     1,     1,     2,    -1,    -3,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     1,     0,     2,     0,    -1,     0,    -1,    -2,    -2,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,    -2,     0,     1,     1,     2,     2,     1,     0,     0,     0,     0,     1,     0,    -1,    -3,    -2,    -1,     1,     2,     1,     0,    -3,     0,     0,     0,    -1,    -1,    -1,     0,     2,     1,     0,     1,     2,     1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     1,     2,     1,     1,    -1,     0,     0,     0,     0,    -2,    -2,     1,     1,     1,     2,     2,     1,     1,     0,    -1,     0,     0,     1,     0,    -1,     0,     0,     1,     2,     1,     0,     1,    -2,    -1,     0,     0,    -1,    -2,    -2,     2,     2,     2,     3,     3,     2,     1,     1,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     2,     1,    -2,    -1,    -3,    -1,     0,     0,     0,    -2,     0,     1,     1,     2,     3,     3,     2,     2,     2,     0,     0,     0,     1,     0,    -1,     2,     1,     0,     1,     2,    -1,    -2,    -2,    -1,     0,     0,     0,    -2,    -2,     1,     1,     1,     1,     1,     2,     1,     2,     3,     0,     0,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,    -2,    -3,    -2,     0,     0,     0,     0,    -1,    -1,     0,     1,    -1,     1,     1,     0,     2,     2,     1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -3,    -2,    -1,    -1,     0,     0,    -2,     0,     0,    -2,    -1,     0,    -1,     0,     0,     1,     1,     0,     0,     0,    -1,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,     0,    -2,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     1,     0,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     1,     2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     2,     2,     0,    -1,     0,     0,     0,     1,     0,     0,     1,     1,     1,     1,     0,    -1,     0,     0,     0,    -1,    -1,    -3,    -3,    -2,     1,    -1,     0,    -1,     1,     2,     0,     1,     1,     0,     0,     1,     0,     1,     0,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     1,    -1,     0,     1,     2,     0,    -1,    -2,    -2,    -2,    -2,    -3,     0,     0,     0,     0,     0,    -1,    -1,     0,    -2,    -2,    -3,    -3,    -2,    -1,    -1,     0,     1,     1,     1,     0,    -3,    -1,    -3,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    27 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     0,     0,    -2,    -1,    -2,    -3,    -3,    -2,    -3,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,     1,     1,    -1,    -1,    -2,    -2,    -1,    -2,    -2,    -5,    -6,    -4,    -3,    -1,     0,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     3,     2,     2,    -1,    -2,     2,     0,    -1,     0,     1,     1,     0,    -2,     0,     0,     1,     0,     1,     2,     0,    -3,    -3,    -2,    -2,     0,     0,     2,     0,     2,     2,    -1,     0,     0,     0,     1,     2,     1,     1,     0,     0,     0,     0,     1,     0,     1,     1,     1,     2,     2,     0,    -1,    -2,    -1,    -1,     2,     1,     2,     1,    -1,    -1,     0,     1,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     1,     0,     1,     1,     0,     1,    -1,    -3,    -1,     0,     1,    -1,     0,     1,     1,     0,     1,     1,     2,     1,     1,     2,     0,     0,     0,     0,     0,     0,     1,     0,     2,     0,     0,     0,    -1,    -2,     0,     0,     1,     0,    -1,     2,     1,     0,     1,     1,     1,     0,     2,     0,    -1,    -2,    -1,     0,     2,     0,     1,     1,     1,     0,    -1,    -1,    -2,    -2,     0,     0,    -1,     2,     0,     2,     1,     1,     1,     0,     0,     2,     3,     0,    -3,    -5,    -1,     1,     1,     0,     0,     1,    -1,     0,    -1,     0,    -2,    -1,     0,     0,     1,     0,     0,     0,     1,    -1,     1,     0,     0,     1,     0,    -3,    -7,    -5,     0,     1,     0,     0,    -2,     0,     0,     0,    -3,     0,    -1,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,     1,     1,     1,     1,     0,    -4,    -8,    -3,    -1,     0,     0,    -1,    -2,     0,     0,    -2,    -3,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,    -1,     1,     1,     1,     1,     2,    -2,    -6,    -6,     0,     0,     0,     0,    -2,     0,     0,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,     0,     0,    -4,    -7,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,    -1,     0,     0,    -2,    -2,    -4,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -3,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,    -2,    -3,    -1,     0,    -1,     0,     0,     2,    -2,    -2,     0,    -1,    -1,    -1,     0,     0,    -2,    -2,    -1,     0,    -1,     0,     1,     1,     0,     0,    -2,    -1,    -1,    -3,    -2,     0,    -1,     0,     1,     0,    -2,     0,     1,     0,    -2,     1,     1,    -1,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     2,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -3,    -2,    -2,    -2,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,     1,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -3,     0,     0,     0,     0,    -1,     0,     2,     1,     0,    -1,     1,     1,    -1,    -2,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,    -2,    -1,     0,     0,    -1,     0,     0,     0,     1,     2,     3,     2,     0,    -1,     0,    -1,     1,    -1,    -1,    -2,    -2,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -2,     1,     0,    -2,    -1,     0,     0,     0,    -2,    -1,     1,     0,     1,     0,     0,     0,     0,     0,     0,     2,     1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     1,     2,     0,    -2,    -1,    -1,     0,     0,     1,     1,    -1,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     2,     1,     0,     1,     1,     1,     0,     0,     2,     2,     0,     0,     2,     0,     1,     1,     0,     0,     2,     0,     0,     0,     0),
		    28 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -3,    -3,    -2,    -1,    -1,    -3,    -3,    -3,    -1,    -2,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -4,    -5,    -6,    -3,    -3,    -1,     2,    -1,     0,    -1,    -2,    -4,    -3,    -1,     1,     1,     2,     1,     0,    -1,     0,     0,    -1,    -1,    -2,    -3,    -4,    -2,    -2,    -1,    -1,     0,    -1,    -1,     1,     1,     0,     0,    -1,    -1,     1,     1,    -1,    -1,    -1,     1,    -1,     1,     0,     0,     0,    -2,    -2,    -1,    -3,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,    -1,     0,     0,    -2,     0,     0,     1,     1,     0,     2,     2,    -2,     0,     0,     0,    -1,    -3,    -1,    -1,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     1,    -1,     1,     1,     1,     2,     1,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,     1,     0,     1,     0,     0,     1,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,    -1,     1,     2,     1,    -1,    -1,    -2,     0,    -1,    -1,    -2,     0,     0,    -1,     1,     1,     0,     1,     0,    -1,    -1,     0,    -1,    -2,    -1,     0,     1,     0,     0,     0,     1,     1,     2,    -1,     1,     1,     0,    -1,    -2,     0,    -2,     0,     0,    -1,     1,     0,    -1,    -1,    -1,     0,    -1,    -2,    -1,     1,    -2,     1,    -1,    -1,     0,     1,     2,     0,     1,    -1,     0,     0,    -3,    -3,     1,     0,    -1,     1,     0,     1,    -1,     0,     0,    -1,     2,     0,    -1,    -1,     0,     0,     0,     0,     0,     3,     1,    -1,     1,     0,     0,     0,    -2,     2,     1,     1,     0,     0,     1,     0,     0,     0,     1,     1,     2,     2,     0,     0,     0,     0,     1,     1,     0,     1,     3,     3,     2,    -1,     0,     0,    -1,     2,     1,     1,    -1,     0,     0,    -1,    -1,     1,     2,     2,     1,     1,     1,     2,    -1,     2,     1,     0,    -2,     0,     1,     2,     1,    -1,     0,     0,    -1,     3,     0,     0,     0,     1,    -1,     0,     0,     2,     1,     2,     2,     2,     1,     1,     1,     2,    -1,    -2,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0,     2,     1,     0,     1,    -1,    -2,     0,     3,     2,     1,     2,     1,     0,     1,     1,     1,     1,    -2,    -3,    -1,    -1,    -2,     2,    -2,     0,     0,     0,    -1,     0,    -3,    -2,    -1,     1,     0,     2,     2,     1,     1,     2,     1,     1,     1,     1,     0,    -1,    -1,    -2,     0,     1,    -2,     2,    -4,    -2,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     2,     1,     2,     0,     1,     0,     2,    -1,    -1,     0,    -2,    -1,     0,     2,    -2,     1,    -4,    -2,     0,     0,     0,    -2,     2,     1,     3,     0,    -1,     1,     2,     2,     2,     2,     2,     0,     2,     0,    -2,    -1,    -1,    -1,     0,     3,     1,    -2,    -1,    -2,     0,     0,    -1,    -2,     2,     0,    -1,     0,     0,     0,     1,     2,     3,     4,     2,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,     1,     0,    -2,    -1,    -1,     0,     0,    -2,    -1,    -1,     0,     1,     0,     1,     0,     0,    -1,     0,     2,     0,    -1,    -2,    -1,     0,    -1,     0,    -1,     1,    -1,     0,    -3,    -4,    -1,     0,     0,    -1,     0,     0,     0,     1,     0,    -2,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     1,    -1,     1,    -1,    -1,    -2,    -2,     0,    -1,     0,    -1,     0,    -1,     0,     0,    -1,    -2,     0,    -2,    -2,    -2,    -1,    -1,    -2,    -2,     1,     1,    -1,     0,     0,     0,    -1,    -3,    -2,    -4,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,     0,    -1,    -2,     0,    -1,     0,     1,    -1,    -2,    -3,     0,    -2,     0,     0,     0,    -1,     1,     0,     0,    -2,     0,     0,     1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     2,    -1,     1,     1,    -1,     0,    -2,     0,     0,     0,    -1,    -1,    -3,    -3,    -2,    -3,    -2,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,     2,    -1,    -2,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,    -1,     0,     2,     0,    -2,    -1,     0,     1,     1,     0,     1,    -1,    -1,    -1,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -4,    -3,    -2,    -2,    -1,    -2,    -4,    -2,    -1,    -2,    -3,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0),
		    29 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -2,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -4,    -4,    -3,    -3,    -5,    -2,    -3,    -4,    -3,    -2,    -3,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -3,    -5,    -2,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,    -2,    -1,    -5,    -4,    -1,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     1,     0,     1,     1,     0,     0,     1,     1,     2,     1,    -2,    -2,    -2,    -1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,     0,     1,     1,    -1,    -1,     0,     0,     1,     1,     0,     2,     1,     1,     0,    -1,     1,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -2,     0,     0,     1,     2,     1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,    -1,     1,     0,    -1,    -1,     0,    -1,     1,     2,     2,     1,     1,     0,     1,     2,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,    -1,     0,    -1,    -2,    -3,    -1,    -2,    -3,    -1,     0,    -2,    -1,     1,     4,     2,     2,     1,     0,     0,    -1,    -1,     1,    -1,    -1,     1,     3,     2,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -1,    -1,     0,    -3,     0,     0,     2,     2,     2,     0,    -1,     0,     0,     0,     0,     1,     1,     1,     3,     2,     0,    -2,    -1,     0,     1,     1,     0,     2,     0,    -1,     0,    -1,     0,    -1,     2,     1,     2,     0,     0,     0,    -1,     0,     0,     1,     3,     2,     1,     0,     0,     0,     1,     0,     0,     1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     1,     2,     0,     0,    -1,    -1,     0,     0,     0,     2,     3,     3,     1,     0,     1,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     1,     3,     3,     2,     2,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     1,     0,    -1,    -1,     0,     0,     1,     3,     3,     2,     2,     1,     2,     1,     1,     1,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,    -2,    -2,    -1,    -1,     1,     0,     1,    -1,     1,     1,     1,     1,     3,     2,     0,     1,     2,     2,     2,     0,    -1,    -1,    -3,    -2,    -1,    -1,     0,     0,    -2,     0,    -1,    -2,     1,     2,     0,     1,     0,     2,     2,     1,     2,     1,     0,     1,     1,     1,     2,     0,     0,    -1,    -3,    -1,    -2,    -1,     1,     0,    -2,    -1,    -2,    -2,     2,     2,     2,     1,     1,     0,     0,     0,     0,     1,     0,     2,     1,     2,     1,    -1,     0,    -2,    -3,    -1,    -2,    -2,     0,     0,    -3,    -1,    -2,    -2,     1,     2,     1,     1,     1,     0,     0,     0,    -1,     0,     2,     2,     1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,    -2,    -1,    -2,    -1,    -1,     0,     1,     0,    -1,     0,     1,    -1,    -1,     0,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,    -2,    -1,    -2,     0,    -1,     0,    -1,     0,    -1,     0,     1,    -1,    -1,     1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     0,    -2,     0,     0,     0,    -2,     1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -2,     0,     0,    -1,    -2,    -2,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -2,    -2,    -2,    -1,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     1,    -1,    -1,    -2,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,    -2,    -2,    -1,     0,    -1,    -1,     0,    -1,    -1,    -2,     0,    -1,     0,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     2,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     1,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0),
		    30 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     1,     0,     0,    -1,     1,     2,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     2,     0,     0,     0,    -1,    -2,    -2,    -3,    -2,    -3,    -2,    -4,    -3,    -4,    -2,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -2,    -2,    -1,    -2,     0,     1,     1,    -1,    -3,    -1,    -1,    -2,    -3,    -1,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,     0,    -1,    -2,     0,    -3,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -2,     0,     0,     1,     0,     0,    -1,    -1,    -3,    -3,    -1,     0,     0,     0,    -1,    -2,     0,    -1,     1,     1,     0,    -1,     1,     0,    -2,    -2,    -1,    -1,    -1,     0,     1,     1,    -1,    -1,     0,    -2,     0,    -4,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,    -3,     0,    -1,    -2,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     1,     0,     1,    -3,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     2,     0,     1,     0,    -1,     0,     0,     1,     1,     0,     2,     1,     2,     0,     0,    -2,     0,     3,    -2,     1,     0,    -1,    -2,    -2,    -1,     0,     0,     1,     0,     1,     0,     0,     2,     2,     2,     0,     2,     2,     2,     2,     0,     0,    -2,    -3,    -1,     0,     0,     2,    -2,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     1,     1,     1,     1,    -1,     0,     2,     1,     0,     0,     1,    -2,    -1,     0,    -1,     0,     2,     1,    -2,    -1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,     2,     0,     0,     1,     1,     0,    -1,    -1,    -2,    -3,     0,     0,     2,    -2,     0,    -3,     0,     1,     0,     1,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     2,     0,    -2,    -3,    -2,    -2,     0,     0,     0,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,    -2,    -1,     0,    -2,    -1,     0,    -1,    -1,    -1,     0,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     1,     2,     1,     2,     1,     0,     1,     0,    -1,     0,    -2,    -1,    -2,    -1,     1,     0,     1,    -2,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     3,     3,     3,     1,     1,     1,     2,     1,     0,    -1,    -1,     0,    -2,     0,     0,     1,    -1,    -2,     0,    -1,     1,    -2,    -3,     0,     0,     0,    -1,    -1,     2,     3,     1,     2,     2,     3,     2,    -1,     2,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -3,    -1,     0,     0,    -1,    -2,     2,     2,     1,     1,     3,     3,     1,     2,     2,    -1,     0,     1,    -1,    -1,     0,    -1,    -1,    -2,    -2,     1,    -2,    -3,    -4,     2,     0,     0,    -1,    -3,     1,     1,    -1,     1,     1,     1,     2,     2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,     1,    -1,    -2,    -2,    -2,     3,     0,     0,     0,    -3,     0,     0,     0,     0,     1,     1,     1,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -1,     0,     1,    -1,    -2,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -3,    -2,    -1,     0,     1,    -1,    -3,    -1,     0,     0,    -1,    -2,    -2,    -1,     1,     0,     0,     1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -3,     0,     0,     0,     0,    -2,    -2,    -2,     0,     1,     0,    -1,    -1,    -1,     0,     1,     2,     1,     2,     1,     0,    -1,    -2,    -2,    -1,     0,    -1,    -1,    -1,     2,     1,     0,     0,    -3,    -1,    -3,    -1,     0,     1,     2,     0,     1,     1,     3,     1,     2,     2,     0,     0,    -1,    -1,     0,     1,     1,     1,    -1,    -1,     1,     1,     0,     0,    -1,    -3,    -3,    -1,     1,     0,     0,    -1,     0,     0,     1,     1,     1,     0,     1,    -1,    -1,    -1,    -1,     1,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     0,     1,    -1,    -1,    -2,    -3,    -3,    -2,     1,     2,     2,     2,     2,     0,    -1,    -3,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -5,    -4,    -1,     0,     0,    -3,    -3,    -2,     0,    -1,    -1,    -1,     0,     0,    -2,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -3,    -2,    -3,    -1,    -2,    -3,    -2,    -1,    -1,    -2,    -3,    -2,    -2,    -4,    -4,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0),
		    31 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,     1,     0,     0,     1,     0,     0,     2,     2,    -3,    -2,    -1,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,    -2,     1,     1,     1,     0,    -2,    -1,    -1,     0,     1,     0,     0,     0,     1,     1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     1,     2,     0,     0,     1,     0,     1,     0,     0,     1,     0,     0,     0,     2,     2,     2,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     1,     0,     2,     2,     1,     2,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     2,     1,    -1,    -1,     1,    -1,    -2,    -2,    -1,     0,     0,    -1,     0,     2,     2,     2,     1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     0,    -1,    -2,    -1,    -3,     0,     2,     2,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,    -1,     0,     1,     1,     0,     0,     1,     0,    -2,    -4,    -2,     0,    -2,    -2,    -3,    -3,    -1,     1,     0,    -1,    -1,     0,     0,     2,     1,     2,     0,     0,    -1,     1,     0,    -1,    -1,     1,     0,     0,    -2,    -6,    -1,     0,    -1,    -2,    -3,    -3,    -1,    -2,    -1,    -1,    -1,     0,     0,     2,     2,     1,     0,     0,    -1,     0,     0,    -1,    -2,     0,    -1,    -1,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -2,    -2,    -2,    -1,    -1,    -2,    -1,    -1,     2,     2,     1,     0,     0,     1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -2,    -2,    -2,    -2,    -1,     0,     2,     1,     1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,     2,     0,     0,    -3,    -1,     0,    -2,    -1,    -3,    -2,    -2,    -1,    -1,     0,     2,     0,     0,     1,     0,    -1,    -1,     1,    -2,    -2,    -1,    -2,     0,     0,     1,     0,     0,    -2,     1,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     2,     1,     0,    -1,    -1,    -3,    -2,    -2,    -2,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     1,     1,     0,     1,     1,     0,    -1,    -2,    -3,    -3,    -2,    -5,    -3,    -1,    -1,     0,     0,     1,    -2,    -2,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -2,     0,     0,     1,     1,    -1,    -1,     1,     1,     1,     0,     0,     0,    -1,     1,     1,     0,     1,    -1,    -1,    -1,     0,     0,     0,    -3,    -2,    -2,    -4,    -2,     0,     1,     1,    -1,    -1,    -1,     0,     2,     1,    -1,     0,    -2,    -1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,    -1,    -3,    -3,     0,     0,     0,     1,     1,     1,     0,    -1,     0,     1,     1,     1,    -1,    -1,    -2,    -2,     0,     1,     1,     2,     1,    -2,     0,     0,     0,    -1,    -3,    -1,     2,     2,     3,     0,     2,     2,     0,     1,     1,     1,     0,     0,    -1,     0,    -1,     1,     1,     2,     1,     2,     0,    -1,     0,     1,     1,     0,     0,    -1,     1,     1,     2,     2,     2,     1,     0,     1,     2,     0,    -1,     0,    -1,     0,     0,     1,     1,     1,     0,     0,     1,    -1,     0,     0,     1,    -1,     0,     0,     1,     2,     2,     1,     2,     1,     1,     1,     2,    -2,    -1,     0,     0,     0,     1,     2,     1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     1,     2,     1,     1,     1,     0,    -2,    -1,    -1,     1,    -1,     0,     1,     0,    -1,    -1,    -2,    -1,     2,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     1,    -2,     0,     0,    -2,    -2,    -2,     0,     0,    -2,    -1,     1,     0,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -3,     0,    -1,     0,    -1,     1,     0,    -2,    -2,    -2,    -3,    -4,    -3,    -5,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -2,    -3,    -5,    -5,    -4,    -3,     1,     0,    -2,    -2,    -2,    -2,    -1,    -3,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    32 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,     0,     0,     0,     0,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,     1,     1,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     2,     1,     2,     1,     0,     0,     1,    -1,    -1,     0,     0,    -2,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,     1,     1,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     1,     1,     1,     2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     2,     2,     1,     2,     1,     2,     0,    -1,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -3,    -2,    -1,    -1,     0,    -1,     0,     0,     1,     1,     1,     2,     1,     1,     1,     0,     0,     1,     0,     1,     0,    -2,    -1,    -1,     0,    -1,    -2,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -1,     0,     1,     0,    -1,    -2,    -1,    -3,    -3,    -1,     0,     0,     0,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -2,     0,    -1,    -3,    -2,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -2,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -2,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -2,    -1,     0,    -1,     0,    -1,    -1,     1,     0,     2,     1,     0,     0,     0,     0,     0,     0,     0,    -3,    -3,    -3,    -2,    -2,    -1,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     1,     0,     1,     2,     3,     1,     0,    -1,     0,    -1,    -1,     0,    -1,    -2,    -3,    -2,    -2,    -1,     1,     0,    -1,    -2,     0,    -1,    -1,    -2,     0,     1,     0,     0,     1,     1,     1,     0,     1,     1,     0,    -1,     1,     1,    -1,    -2,    -2,     0,     0,     0,     1,     0,     0,     1,     1,     0,    -1,     0,     0,     2,     2,     1,     0,     1,     2,     2,     1,     2,     0,     0,     1,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     1,     2,     0,     1,     1,     2,     0,     3,     1,     1,     0,     0,     2,     0,    -1,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,     1,     0,    -2,     1,     2,     0,     0,     1,     0,     0,    -2,     1,     0,     1,     0,     0,     0,     1,    -2,     0,     1,     1,     1,     0,    -1,    -1,     0,    -1,     0,    -1,     1,     2,     1,    -1,    -1,     0,    -1,    -1,     1,     2,     0,     3,     0,    -1,    -1,    -1,    -2,     0,     0,     1,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     1,     1,     0,    -1,    -2,    -2,     0,    -1,    -2,     0,     2,     2,     0,    -1,     0,     0,    -1,     0,     1,     1,     1,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     1,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,     0,     1,     1,     2,     1,     0,     0,     1,     1,    -1,    -1,    -1,     0,     0,     1,     0,     1,    -1,     0,     0,     0,    -2,    -1,    -2,    -2,    -2,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,     1,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -2,    -2,    -4,     0,     0,    -1,     0,    -1,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0),
		    33 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     1,     1,     1,     0,    -1,    -1,    -1,     0,    -2,     0,     0,     0,     0,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     1,     0,     1,     1,     1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -2,     0,     0,     0,     1,     1,     1,     0,     1,     1,     1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     3,     1,     1,     0,     1,     1,     0,     1,     1,    -1,    -1,     0,     1,     0,    -2,     0,     1,     0,     0,     1,    -1,     0,    -2,    -2,    -1,     0,     0,    -1,     2,     1,     0,    -1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,    -1,    -2,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,    -1,     0,     1,     2,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     1,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,    -2,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     0,     0,    -1,    -2,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     0,     1,     1,     1,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,     1,     0,     1,    -1,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -2,     0,    -2,    -1,     1,     2,     1,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     1,     0,    -1,     0,     0,     2,     3,     0,     1,    -1,     0,     0,     1,     0,    -1,    -3,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,     1,     2,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    34 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,     0,     1,     0,    -3,    -2,     0,    -1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     2,     0,    -4,    -5,    -1,     0,     2,     0,     1,    -1,     0,     0,     1,    -2,     0,    -2,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,    -1,     1,     1,     1,    -3,    -4,    -3,    -1,     1,     0,     0,     1,     1,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,     1,     0,    -1,    -2,     0,     1,     1,    -1,    -2,    -4,    -1,     0,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,     0,    -1,     1,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,     2,     0,     0,    -1,    -3,    -2,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     2,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -2,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,    -1,     0,     1,    -1,     0,     0,     1,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -2,     0,     0,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -1,    -2,    -2,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     2,     0,    -1,     0,     1,     1,     1,     0,    -1,     1,     1,     0,    -1,    -2,    -1,    -2,    -2,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     1,     1,    -1,     0,     1,     2,     1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     2,    -1,     0,    -1,     1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     1,     1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,     0,     1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,    -1,    -2,    -1,    -2,    -1,    -2,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -2,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -2,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,    -1,     1,     0,     1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,     0,     0,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     1,     1,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,    -1,     2,     1,     1,     1,     1,     1,     0,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,     1,     1,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,    -2,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0),
		    35 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -4,    -2,    -1,    -1,    -1,     0,     0,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -2,    -3,    -2,    -1,    -1,     0,    -1,    -1,    -1,     1,     2,     1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,     0,    -1,     0,     1,    -1,    -2,    -1,     1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,    -1,     0,    -2,    -1,    -1,    -1,    -1,    -3,    -3,     0,     1,    -1,    -1,     0,    -1,    -2,     1,     0,     0,     0,     1,    -1,    -2,     1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,     0,     0,     0,     0,     1,    -1,    -2,     1,    -2,    -1,     0,     0,     2,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -3,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,     1,    -1,    -1,     1,     1,     1,     1,     0,     1,     1,     1,     2,     2,     1,     1,    -1,     1,     0,     0,    -1,    -1,    -1,    -2,     0,     1,     0,     0,     0,    -1,    -1,     0,     1,     1,     2,     3,     2,     2,     2,     2,     2,     1,     3,     2,    -2,     0,     0,     0,     0,    -1,     0,     0,     1,     1,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,     1,     2,     2,     2,     2,     2,     1,     3,     2,     1,     2,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -1,     0,     0,     1,     0,     2,     2,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,     1,     1,     0,    -1,    -1,    -2,    -2,    -4,    -7,    -4,    -3,    -3,    -2,    -1,     1,     2,    -1,     0,     0,     0,     0,     0,    -1,    -2,     1,     0,     0,     2,     1,     1,     0,     0,     0,    -1,     0,    -2,    -3,    -4,    -2,    -3,    -3,    -1,     0,     1,    -1,     1,     0,     0,     0,     1,     0,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -2,    -3,    -2,    -2,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     1,     2,     1,     0,     2,     1,     1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     1,     0,    -1,    -1,    -2,    -1,    -1,     1,     0,    -1,     0,     0,    -1,     0,     1,     2,     0,     1,     0,     1,     0,    -1,    -1,     0,    -2,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,    -1,     0,     0,    -2,     0,     1,     1,     0,    -1,     0,     1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,    -2,    -2,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -1,     0,    -1,    -1,    -1,    -2,     1,     1,    -1,    -1,     0,    -1,     0,    -1,     0,     1,    -1,     0,     1,     0,    -1,    -2,    -1,     0,     0,     0,    -2,     1,     1,     0,    -1,     0,    -2,    -2,    -2,     0,     1,    -1,    -1,     0,     0,     0,     1,     0,    -1,     1,     2,     2,     2,    -2,    -2,     0,     0,     0,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     1,    -3,    -1,     0,     0,     0,     1,     1,    -1,     0,     0,     2,     3,    -2,     0,     0,     0,     0,    -1,     0,     1,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     2,     3,     1,     0,     0,     0,    -1,     0,     0,     1,     1,    -1,    -2,     0,     0,     0,     1,     0,     0,     1,     0,     1,     0,    -1,     0,     0,    -1,     2,     3,     3,     3,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     1,     1,    -1,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     3,     3,     3,     4,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -1,    -1,    -1,     0,     1,     1,     0,     1,     0,     0,     0,    -1,    -1,     0,     1,     2,     1,     1,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -2,    -2,    -1,    -1,     0,     2,     1,     0,    -1,    -1,    -1,     0,     0,    -1,     1,     1,     2,     2,     0,     0,     0,     0,     0,     0,     0,    -1,    -3,    -4,    -3,    -3,    -3,    -3,    -2,    -2,    -3,    -5,    -1,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,     0),
		    36 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,     0,     0,     1,    -1,     0,     0,     1,     1,     1,     3,     1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     1,     1,     2,     1,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     2,     1,     1,     0,     2,     2,     2,     1,     2,     0,     0,     0,     0,    -2,     0,    -1,     1,     2,     2,     0,    -1,    -1,    -2,    -3,     0,     1,     1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -2,    -1,    -1,     0,     0,     0,    -3,     0,     1,     2,     1,    -1,    -2,    -1,    -2,    -3,    -4,    -2,    -2,    -1,     0,    -1,     0,     3,     2,     0,    -2,    -2,    -4,    -3,    -1,     1,     0,     0,    -1,    -1,     1,     2,     1,    -1,    -1,    -1,    -1,    -3,    -2,     0,     0,    -1,    -1,     0,     1,     1,     1,     1,    -1,     0,    -2,    -3,     0,     0,     0,     0,     1,     0,     0,     1,     1,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,     1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -2,    -4,    -3,    -1,    -1,     1,     1,    -1,    -1,     0,    -2,     0,     0,     1,    -1,    -3,    -3,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     1,    -1,    -2,    -3,    -3,    -1,     0,     0,     0,     0,     0,    -1,    -3,     0,    -1,    -1,    -1,    -3,    -3,    -1,    -1,    -2,     0,     0,    -1,    -1,     2,    -1,     0,     0,    -2,    -2,    -1,     0,    -1,     0,     1,     0,    -1,    -2,    -3,    -4,    -5,    -4,    -4,    -4,    -3,    -2,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -3,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -3,    -3,    -3,    -3,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -2,    -2,    -1,    -1,     0,    -1,    -1,     0,    -3,    -3,    -3,    -2,    -2,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     1,     1,     0,     2,    -1,     0,    -1,     1,     0,     0,    -1,    -1,     1,     0,    -1,    -3,    -3,    -2,     0,     0,     0,    -2,    -1,    -1,    -1,    -2,     0,     0,     1,     2,     0,     1,     0,     0,     0,     1,     2,     0,     0,     0,     2,     2,    -2,    -3,    -2,     0,     0,     0,     0,    -2,    -1,     0,    -2,     0,    -1,     1,     1,     0,     0,    -1,    -1,     0,     0,    -3,     1,     1,     0,     2,     1,     0,     0,    -1,    -2,     0,     0,     0,     0,    -2,     0,     0,    -1,     0,     1,     1,     1,    -1,    -1,    -1,     0,    -2,    -1,    -2,     0,     1,     1,     2,     1,     0,    -2,    -2,    -3,    -2,     0,     0,     0,    -1,    -1,     1,     0,     1,     0,     1,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     1,     2,     1,     0,    -2,    -2,    -3,    -2,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     1,     1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     1,     2,    -1,     0,    -2,    -2,     0,    -2,     0,     0,     0,     0,     2,     0,    -1,     0,     0,     2,     1,    -1,     0,    -1,     0,     2,     0,     1,     1,     1,     0,     0,    -3,    -2,    -2,    -2,     0,    -1,     0,    -1,    -1,     0,     1,    -1,     0,     0,    -1,     0,     1,     1,     0,    -2,    -1,     1,     0,     0,     1,    -1,    -1,    -1,    -3,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,     1,     1,     0,     0,     0,    -1,     0,     1,     1,    -1,     0,     0,    -2,    -1,    -2,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -2,     0,     1,     1,     0,     1,     1,    -1,    -2,     1,     2,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,     1,     2,     0,     0,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    37 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -3,    -3,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -2,    -3,     0,    -1,     1,     3,     1,    -2,    -2,    -1,     1,    -1,     0,    -3,    -3,    -2,    -3,    -3,    -2,    -2,    -2,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -1,    -2,    -1,    -1,    -3,     0,     1,     0,     0,     2,     0,    -1,    -2,     0,    -2,    -1,     0,     0,     0,     1,     1,     0,     1,     1,     0,     0,     0,    -2,    -1,     0,    -1,    -2,    -2,     0,     0,    -3,    -2,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     2,     1,     0,     2,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     1,    -1,    -1,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     1,     0,     0,     3,     0,     0,     0,     0,     0,    -1,     1,     2,     1,     1,     1,    -1,    -1,     0,    -1,     0,     1,     1,     2,     0,    -1,    -1,     1,     0,     2,     1,     1,     3,     1,     1,    -1,     0,     1,     0,     1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     2,     1,    -2,     0,    -1,     1,     0,     1,     2,     2,     2,     0,    -1,     0,    -1,     0,     0,     1,     0,     0,     0,     1,    -1,    -1,    -1,     0,    -1,     1,     1,    -1,    -3,    -2,    -1,     2,     0,     0,     0,     3,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     1,     0,    -1,     1,     0,     0,     1,     1,    -2,    -1,     1,    -1,     1,     0,     1,     1,     3,     1,     1,    -1,    -1,    -1,    -1,     1,     1,     0,    -2,     1,    -1,     0,     0,    -1,    -1,     2,     1,     1,     0,     0,     2,    -1,    -1,     0,     1,     3,     3,     0,     1,    -1,    -1,    -1,     0,     1,     1,    -1,    -3,    -1,    -1,     0,     1,     0,     1,     1,     1,     1,     2,     2,    -1,    -1,     0,     0,     0,     2,     1,    -1,     0,     0,     0,    -1,     0,     1,     0,    -2,    -2,     0,    -1,    -1,     0,     0,     2,     1,     0,     1,     1,     1,    -2,    -1,    -1,     0,     0,     1,     0,     2,     1,    -1,     1,     1,     2,     0,     0,    -3,    -1,    -1,     0,     0,     0,     0,     1,     0,     2,     3,     2,     1,    -4,    -2,     0,     0,     0,    -1,     0,     1,     0,    -1,     0,     1,     1,    -1,    -2,    -3,    -2,     1,     1,     0,     0,     0,     0,     1,     1,     3,     1,     0,    -4,    -1,    -2,     1,     0,     1,    -3,     0,     0,    -1,     1,     1,     0,    -1,    -2,    -5,    -2,     1,     1,     0,     0,     0,    -1,     0,     1,     1,     0,    -2,    -1,     0,    -1,     0,     1,     0,    -2,    -1,     0,     1,     0,     0,     0,    -3,    -5,    -5,    -1,     2,     0,    -1,     0,    -1,    -1,    -1,    -2,    -4,    -2,    -1,    -2,     0,     0,     0,     1,     0,    -1,     1,     2,     1,     1,     0,    -3,    -4,    -6,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -3,    -2,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,     0,    -2,    -3,    -3,    -3,     0,    -1,     0,     1,     1,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,    -2,    -2,    -3,    -2,     0,     0,     1,     1,     0,     0,     2,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     1,     0,     1,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -1,    -1,    -1,     1,     0,     1,     1,     1,     1,     0,     0,     1,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -3,    -2,    -1,    -2,    -1,     1,     1,     1,     2,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     1,     1,     0,     0,    -2,    -2,    -1,     1,     1,     0,    -1,     0,     1,     1,     1,     0,     0,     0,     0),
		    38 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -2,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,     1,     1,    -1,     0,    -2,    -1,     0,    -1,     0,     0,     0,    -2,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     1,     0,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     2,     2,     0,     0,    -1,     0,    -1,     0,    -1,     0,     1,     2,     2,     1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     1,     1,     0,    -1,    -1,     0,    -1,     0,     0,     1,     1,     1,     1,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     1,     1,     1,     0,    -2,    -1,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     1,     0,     0,    -1,     0,     0,    -1,     0,     1,     0,    -1,    -1,     1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     1,     1,     0,     0,     0,    -2,    -1,    -2,     0,     0,    -1,    -2,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -2,    -1,    -1,     1,     1,    -1,    -3,    -2,     0,     0,     1,     1,     0,     1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     2,     1,    -1,    -1,     0,     1,     1,     1,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,     1,     1,     1,     1,     0,    -1,    -2,    -1,     0,    -2,    -3,    -2,    -1,     0,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,     0,     0,     0,     1,     2,     3,     2,     1,     1,     0,    -1,    -1,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     1,     1,    -1,    -1,    -2,     0,     1,    -1,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     2,     1,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     2,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,    -1,     0,     0,    -1,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     2,     1,     2,     1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     1,     0,     0,     0,     1,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    39 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,     0,    -1,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     1,     0,     0,     1,    -1,    -2,    -1,    -2,    -3,    -1,    -1,    -2,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,    -1,     1,     1,     1,     0,     0,     2,     0,    -1,    -2,    -1,    -3,    -1,    -2,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     2,     1,     0,     0,     1,    -1,    -2,    -1,    -2,    -1,    -2,    -3,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     1,     1,    -1,    -2,    -1,    -2,    -1,    -1,    -2,     0,     0,    -1,    -1,     0,     0,     0,     0,    -2,     0,     0,    -1,     0,     1,     1,    -1,    -1,     1,     0,     1,     1,     0,    -1,     0,    -1,    -2,    -1,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     2,    -1,     1,     0,     1,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -2,    -1,     0,    -3,    -3,    -2,    -1,     0,    -1,     0,    -2,    -1,     1,     0,     0,     2,     1,    -1,    -2,    -1,    -1,    -1,     0,     1,     1,     0,     1,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -3,     0,    -1,     0,    -2,    -1,     1,     0,     1,     1,    -1,    -1,     0,    -1,    -2,    -1,     0,     1,     1,     0,     1,     0,    -1,     0,     1,    -1,    -1,     0,    -2,    -1,    -1,     0,    -2,    -1,     0,    -1,     1,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,    -1,     0,     1,     0,     1,     1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     2,     0,     1,     0,     0,     0,     1,     1,     1,     0,     1,    -1,    -2,    -1,     0,     1,     0,    -1,     1,     0,     0,     1,    -2,    -1,     0,     0,     0,     0,     1,     1,     1,     1,    -1,     0,     0,     0,     1,     1,    -1,     0,    -2,    -2,    -1,     1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,     0,     0,    -1,     0,     2,    -1,     1,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     2,     1,     0,     0,    -1,     0,     1,     0,    -1,    -2,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     1,     1,    -1,    -1,     0,     1,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     1,     1,     0,    -1,     0,     1,     1,     0,     0,     1,     1,     1,    -1,     0,     1,     1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     1,     0,     1,     1,     1,     2,     1,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -1,     0,     0,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -2,    -2,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,     2,     0,     0,    -1,     0,     2,     0,    -2,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,    -3,    -3,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -2,    -1,     1,     0,     0,    -1,     0,     1,    -1,    -3,     0,     0,     0,    -1,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,     1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     1,    -2,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,     2,     2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,     2,     0,     2,     3,     1,     1,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -2,    -2,    -2,     0,     1,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,     1,     1,    -1,    -2,    -1,    -2,    -1,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,    -1,    -1,     1,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0),
		    40 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -2,    -2,    -1,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -3,    -1,    -1,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -1,    -1,     1,     0,    -1,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,     1,    -1,     0,    -1,    -1,     1,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     1,     0,     0,    -2,    -2,     0,    -1,    -1,     1,    -1,    -1,     0,     0,    -1,     1,     0,     1,     0,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     1,     1,     0,    -1,    -2,     0,     0,    -1,     0,    -1,     0,     0,     0,     1,     2,     2,     0,     0,     0,     1,    -1,    -1,    -2,     1,     2,    -1,     1,     0,     1,     1,    -1,     0,     0,     0,     0,    -1,     2,     0,     1,     0,     1,     1,     1,    -1,     0,     1,     0,     1,    -2,    -3,    -2,     0,     0,     0,     1,     0,    -2,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     1,     0,    -1,     0,     1,     0,     2,    -1,     0,     0,     0,    -3,    -2,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,    -1,    -2,     0,     0,     1,     0,     0,     0,     0,    -1,     1,     1,     2,     0,     0,    -2,    -2,     0,     0,     3,    -1,     0,    -1,    -2,     1,     2,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     1,     1,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -1,     2,     1,     1,     1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     1,     1,     0,     0,     0,     0,    -2,     0,     0,     1,     1,     1,    -1,     1,     1,     1,     2,     1,     0,     0,    -2,    -1,    -1,    -3,    -2,    -2,     1,     0,     0,     1,     1,     1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     2,     2,     3,     2,     1,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,     0,     1,     1,     0,     0,     2,     0,     0,    -2,     0,     0,     0,    -1,    -1,     0,     1,     0,     1,     2,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -2,     0,     0,     1,     2,     1,     2,     2,     0,    -2,    -1,     0,     0,    -1,    -1,     1,     0,     1,     2,     1,     0,     1,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,    -1,    -1,     1,     1,     0,     1,    -1,    -3,     2,     0,     0,    -1,    -2,     0,    -1,     0,     0,     1,     1,     0,    -1,    -2,    -2,    -1,     1,     0,     0,    -1,    -1,     0,    -1,     2,    -1,     0,    -1,    -2,     2,     0,     0,    -1,    -2,    -1,    -2,     0,     1,     3,     1,     0,    -1,    -2,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,    -1,     0,     2,     1,     1,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     2,     0,     1,     0,     0,    -2,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     1,     1,     3,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -1,     1,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,    -2,    -1,    -1,    -1,     1,    -1,    -1,    -1,     1,     0,     0,     0,    -2,     0,    -2,     0,     0,     0,     1,     1,     1,    -1,     0,     0,    -1,     0,    -1,    -2,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     1,     1,     0,     0,     0,    -2,    -2,    -1,     0,     0,     0,     1,     1,     1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     1,     1,     1,     1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -2,    -2,    -2,    -2,    -3,    -1,    -1,    -3,    -3,    -3,    -3,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -2,    -2,    -3,    -2,    -2,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0),
		    41 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     2,     2,     3,     2,     1,     1,     3,     2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     1,     2,     0,    -1,    -1,     1,     1,     0,    -3,    -3,     0,     0,     0,     1,     2,     1,     1,     1,     2,     2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,    -1,     0,    -1,    -2,    -2,     0,     2,     2,     1,     1,     0,     0,     1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     1,     1,     0,     1,     1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     1,     2,     0,     0,    -1,    -1,     1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -2,     0,    -1,    -2,    -2,     0,     1,     1,    -1,     0,     0,    -1,     1,     0,     0,     0,    -3,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,     0,    -1,    -2,    -1,    -1,     0,     3,     0,    -1,    -1,     0,     1,     1,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -2,     0,    -1,    -1,     0,     0,     1,     1,     0,    -1,    -1,     0,     1,     1,     1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,    -2,     0,    -1,    -2,    -1,     1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     0,     1,    -1,    -2,     0,     0,     0,    -2,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -4,     0,     1,     0,    -1,    -3,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     1,     1,     0,    -2,    -4,    -2,     1,     0,    -1,    -2,    -3,    -2,    -2,    -2,    -1,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     2,     1,    -1,    -2,    -3,     0,     0,     0,     0,    -2,    -3,    -3,    -2,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -4,    -3,    -4,     0,    -1,    -1,    -2,    -3,    -4,    -2,    -2,    -1,    -1,    -2,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     2,     0,    -1,    -1,     0,    -2,    -3,    -1,     0,    -1,    -1,    -2,     0,     1,     1,     0,     0,    -2,     0,    -3,    -1,    -1,     0,     0,     0,     0,    -1,     2,     0,     0,     1,    -1,     0,    -3,    -3,    -1,     0,     0,     1,     0,     0,     1,     2,     0,    -1,     0,     0,    -1,    -2,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,    -1,    -2,     0,     0,     0,     2,     0,    -1,     1,     1,     0,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     1,     1,    -3,     0,    -1,     0,     3,     1,     0,     0,     1,     1,     1,     1,     1,     2,     1,     1,     1,     2,     1,     0,    -1,    -1,     0,     1,     1,     0,     2,     2,     1,     0,     1,     1,     1,     2,    -1,     0,     1,     0,     0,     0,     0,     1,     0,     1,     1,     0,    -1,     0,     1,    -1,     0,     1,     1,    -1,     1,     1,     3,     2,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     2,    -1,    -2,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -4,    -4,    -3,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -2,    -1,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -2,     0,     1,    -1,    -4,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -2,    -2,     0,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    42 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     2,     0,     0,     1,     1,     1,     2,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     1,     1,     2,     0,     0,     0,    -1,     0,     0,     2,    -1,     0,     0,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     1,     3,     1,     0,     1,     0,    -1,     0,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     2,     1,     1,     1,     1,     1,     0,     0,     1,     1,     0,    -1,    -1,    -1,     0,    -3,    -1,     0,     0,     0,    -1,     0,     1,     1,     2,     1,     0,     1,     0,     0,    -1,     0,     1,     1,     1,     1,     0,     1,     1,    -1,    -3,    -3,     0,    -2,     0,     0,     0,     1,    -1,     0,     1,     1,     1,     1,     0,    -1,     0,     1,     1,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,    -2,     0,     1,    -3,    -1,    -1,     1,     1,     0,     0,     0,     1,     0,    -1,     0,    -1,     1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     2,     1,     0,    -2,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,     0,    -1,     1,     0,    -2,    -1,    -1,     0,    -1,     2,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,     0,     1,     0,     0,    -2,     0,     0,     0,    -1,     0,    -1,     1,    -1,    -2,     0,    -1,    -2,    -1,     0,     0,     0,    -1,     1,     2,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     1,    -1,     1,     2,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,     1,     1,     0,    -1,     0,     0,     0,    -1,     0,     1,     1,     2,     1,     1,     1,     1,    -1,    -1,     2,     0,     0,    -1,     0,     0,    -1,    -2,     0,     2,     2,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     2,     2,     1,     2,     2,     2,     2,     0,     1,     1,     0,    -1,     1,     0,    -1,    -1,     0,     0,     2,     1,    -1,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     2,     2,     1,     1,     1,     0,     0,     0,     1,     0,     0,     1,    -1,    -1,    -1,     0,     1,     1,     1,     0,     1,    -1,    -2,    -1,     1,     0,     1,     2,     2,     2,     3,     1,     3,     1,     1,     2,     1,     0,     0,     1,     0,    -1,    -1,    -1,     0,     1,     2,     2,     1,     1,     0,     0,     1,    -1,     0,     2,     3,     2,     1,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,     2,     1,     0,     0,    -1,     0,     0,     1,     2,     3,     2,     1,     0,     1,     1,    -1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     2,     1,     1,     1,    -2,     0,     0,     0,     4,     4,     4,     1,     1,     1,     0,     0,    -1,     0,     1,     0,    -1,     0,     0,     0,    -1,    -2,     0,     1,     0,     1,     1,     1,     0,    -1,     1,     3,     3,     3,     2,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     1,     0,    -2,     0,     0,    -1,    -1,     0,     0,     0,     0,     2,     3,     3,     2,     2,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     0,     0,     2,     4,     3,     4,     1,     1,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,    -1,    -2,    -2,     0,     0,     2,     3,     5,     4,     3,     1,     0,     1,    -1,     0,     1,     1,    -1,     0,     0,     0,    -1,    -1,    -3,    -3,    -1,    -1,     0,    -2,    -2,    -1,    -1,     1,     2,     2,     3,     3,     2,     1,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,     1,     0,     0,    -1,     0,     2,     3,     3,     3,     3,     2,     1,     1,     1,     0,    -1,    -2,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -3,    -1,    -2,    -2,    -2,    -2,    -2,    -2,    -1,    -2,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,     0,     0,     0,     0),
		    43 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,    -3,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     2,     0,     0,     2,     2,     1,     1,    -1,     0,    -1,    -1,    -3,    -3,    -1,     0,     0,     0,     1,    -2,     1,     1,    -1,    -1,    -2,     1,     1,     2,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -1,     0,     2,    -2,    -3,    -3,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     1,     1,    -1,    -2,     0,     1,    -1,    -1,     2,     0,    -3,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,     0,    -1,    -2,     0,     1,     1,     1,     2,     1,     1,     1,     1,     1,     1,     2,    -3,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,     1,     1,     0,    -1,     0,     0,     3,     1,    -4,    -2,    -1,    -1,     0,     1,     1,     0,     0,    -1,     0,     0,    -1,     1,     0,     1,     1,    -1,    -1,     0,     0,     1,     2,     0,    -1,     1,     1,     0,    -5,    -3,     0,     0,    -2,     0,    -1,     1,     0,    -1,    -2,    -2,     0,    -2,     0,     3,     2,     1,     0,     1,     0,     0,     0,     1,     0,     2,     1,    -2,    -4,    -3,    -1,     0,    -2,     0,     1,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -1,     2,     3,     3,     1,    -1,    -1,    -1,    -1,     0,     1,     0,     1,    -2,    -2,    -2,    -1,     0,    -1,     0,     1,     0,    -1,    -3,    -3,    -1,    -2,    -4,    -1,     0,     3,     2,     1,     1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -6,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -3,    -1,    -1,     1,     1,     4,     2,     0,     1,     1,    -1,     0,    -1,    -4,    -4,    -4,    -2,    -2,     0,     0,     0,    -4,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,     0,     1,     3,     1,     2,     1,     1,     1,     0,    -1,    -2,    -1,    -3,    -3,    -2,     0,     0,     1,     0,    -2,    -2,    -2,    -1,    -1,    -1,     0,    -2,    -1,     0,     1,     1,     2,     1,     0,    -1,    -1,    -1,    -2,    -1,     0,    -2,    -2,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,    -2,    -2,     1,     2,     2,     2,     2,    -1,    -2,    -2,    -1,    -1,     0,     1,     1,     1,    -2,     0,    -1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,     2,    -1,    -2,    -1,    -1,     0,    -1,    -1,     1,     0,     1,    -3,    -2,    -1,     0,     0,     1,     1,     1,    -1,    -1,     0,    -2,    -1,     0,     1,     0,     1,     0,    -2,    -2,    -1,    -1,     0,    -2,     0,     0,     0,     0,    -3,    -1,    -1,    -1,     0,     1,     1,     0,     0,     0,     1,    -1,     0,     1,     2,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     1,    -1,    -1,    -1,    -2,     0,    -1,     0,    -1,     1,     2,     1,     2,    -1,     1,     0,     1,     1,     0,    -1,    -1,    -2,     0,     0,     1,     1,     0,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -1,    -2,     1,     0,    -1,    -1,     1,     1,     0,     1,     0,    -2,    -1,    -1,     1,     1,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,     1,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -2,    -1,     0,     0,     0,     0,     1,    -1,    -1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -2,    -2,    -3,     0,     0,     0,     0,     1,     2,     0,     0,     2,     0,     1,     0,     1,     1,    -1,     1,    -1,     0,     1,     0,     1,     0,    -1,    -1,    -1,    -2,     2,     0,    -1,     0,     0,     0,     1,     2,     0,     0,     1,     0,    -1,    -1,     0,     3,    -1,     0,     2,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     2,     2,     3,     1,     0,    -1,     1,     0,     0,     1,    -1,    -3,    -3,    -4,    -2,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,     1,     1,     1,     0,    -2,    -1,     0,     0,     1,    -1,    -1,    -2,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0),
		    44 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -2,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -1,    -1,    -1,    -1,     0,    -2,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -2,    -2,    -2,    -1,     1,    -1,    -2,    -4,    -2,     0,    -1,     0,    -2,    -2,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,    -2,    -3,     0,     0,    -3,    -3,    -4,    -3,    -2,    -1,     0,     0,     1,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -2,     0,     2,    -1,    -1,     0,    -1,    -6,    -3,     0,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     1,     3,     0,    -2,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,    -4,    -5,    -2,     1,     1,     0,     0,     1,     1,    -3,     1,    -2,     0,    -2,     0,    -1,     0,     3,    -1,    -1,    -1,     0,     0,     1,     0,     1,     0,    -2,    -5,    -5,     0,     2,     1,     0,     0,     1,    -1,    -1,     1,    -3,    -1,    -2,     0,    -1,     0,     1,    -1,     1,    -1,     0,    -1,     0,     1,     1,     0,    -2,    -6,    -2,     1,     1,     0,     0,     1,    -1,     0,     2,     1,    -2,     0,    -2,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,     2,     1,    -3,    -3,     1,     2,     1,     1,     0,     1,     1,     2,    -2,    -2,    -1,     0,    -1,    -1,     0,     1,     2,     0,    -1,     0,     0,    -1,     0,     0,     2,    -1,    -3,    -2,     1,     2,     1,     0,     0,     1,     1,     1,    -3,    -1,     0,     0,    -1,    -1,    -2,    -1,     1,     2,     0,     1,    -1,     0,     0,     1,    -1,    -2,    -3,    -2,    -1,     0,     0,    -1,     1,     0,     0,     1,    -1,    -1,    -1,     0,     0,    -1,    -2,    -3,    -1,     0,     1,     1,    -1,     0,     1,     1,     1,    -3,    -2,     0,     0,     0,     1,     0,     1,     0,     1,    -2,    -1,    -3,    -2,     0,     0,    -2,    -2,    -2,    -1,     0,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     1,    -1,     1,     1,     1,     0,    -1,    -3,    -2,    -2,     0,     0,     0,     0,    -2,    -2,     0,     0,     0,     0,     1,     0,     1,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,    -2,    -2,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     1,     1,     0,     0,     1,     0,    -1,     0,     0,     2,    -3,    -1,    -1,     0,    -1,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,    -1,     0,     1,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,     0,     0,     0,    -2,     0,     0,    -1,    -1,     0,    -1,     2,     3,    -1,    -1,    -2,    -1,    -1,    -3,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,     1,     1,     0,     1,     0,     0,     0,    -1,    -1,     2,     1,    -1,    -2,    -1,    -1,    -2,    -2,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,     1,     0,    -1,     0,     0,     0,    -2,    -2,    -2,    -2,    -1,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -2,    -3,    -1,     0,     0,     0,    -1,    -1,    -2,     3,     0,     0,     2,     2,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -2,     0,     0,     0,     0,     1,    -1,    -4,    -1,     0,     0,     0,     0,    -1,    -2,     1,     2,     1,     1,     0,     1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     1,    -1,    -1,     1,     0,     0,     0,     0,    -1,    -2,    -4,     1,     1,     1,     1,     1,     0,     1,     0,     0,     0,     1,    -1,    -1,     0,     0,     1,     0,     1,    -1,     0,     1,     0,     0,     0,     0,     0,    -3,    -3,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     1,     1,    -1,    -3,    -1,    -1,     1,     0,     1,    -1,     1,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -2,     0,     0,    -1,     0,     0,     1,     1,     0,    -1,    -1,    -3,    -2,    -1,     0,    -1,     1,     2,     0,    -1,     0,     0,     0,     0,     0,    -2,     0,    -2,    -2,    -3,    -1,    -2,    -2,    -1,    -2,    -3,    -4,    -5,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,     0,    -1,    -2,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0),
		    45 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -2,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -2,     0,     0,     0,     0,     0,     0,     1,     3,    -1,    -1,    -1,     0,     1,     0,    -2,    -2,    -3,    -2,    -1,     1,     0,     0,     0,     0,     1,    -2,    -2,     0,     2,     2,     0,     0,     0,    -1,     2,     0,     0,    -1,    -1,    -1,     0,     0,    -2,    -2,    -2,    -1,    -1,    -2,    -2,     0,     2,     0,     0,    -1,     0,     2,     2,     0,    -1,     0,     0,    -2,     3,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -2,    -1,    -1,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     1,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     2,     2,     1,     2,     2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     1,     0,     1,     1,     0,    -1,     0,     1,     1,     1,     1,     0,     3,     1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     2,     3,     1,     2,     1,     1,     0,     1,     1,     0,    -1,    -3,    -2,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,    -1,     1,     0,     1,     1,     3,     3,     1,     1,     0,     0,    -1,    -1,    -1,     1,    -1,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     1,    -1,    -5,    -5,    -3,    -3,    -3,    -1,     0,     1,     0,     1,     0,     0,     0,     1,     1,     1,    -1,    -1,    -1,    -2,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -3,    -3,    -5,    -4,    -4,    -3,    -3,    -1,     0,    -1,     0,     0,     0,     1,     1,     0,    -2,    -2,    -2,    -1,     0,    -1,    -2,     0,     1,     0,    -1,     1,     0,    -1,    -2,    -4,    -3,    -6,    -4,    -2,     0,    -1,     0,     0,     0,     2,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     1,     0,     1,     1,     0,     0,     1,     2,     1,     1,     0,    -2,    -3,    -1,     0,    -1,     0,     0,     0,     1,    -1,    -2,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,     1,     1,    -1,     0,     1,     1,     0,     0,     1,     1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     1,     0,    -1,    -2,     0,    -1,    -1,     1,     0,    -1,    -1,     0,    -1,     0,     2,     0,     0,     1,     2,     0,     0,     0,     0,    -1,    -2,     0,     0,    -2,     2,     0,     0,    -2,    -2,    -2,    -1,     0,     0,    -1,     1,     1,     0,     0,     2,     1,     0,    -1,     0,     1,     0,     0,     0,    -1,    -3,    -1,     1,     0,     1,     3,     1,     0,     0,    -1,    -3,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     0,    -2,    -2,     0,     0,    -1,    -1,     0,     0,    -2,     0,     0,     0,     1,     2,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -2,     0,     0,     2,    -2,    -1,     0,     1,     2,     1,     2,     1,     1,     1,     1,     0,     0,     0,    -1,     0,     1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     1,    -3,    -2,     0,     0,    -1,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     1,    -1,     0,    -2,    -1,    -1,     1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     1,     1,     0,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,     0,    -1,     0,     1,     1,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -3,    -2,    -1,    -3,    -3,    -1,     0,    -1,    -1,    -2,    -1,     0,     1,     1,     0,     1,     0,     0,    -2,    -1,     0,     0,     0,     0,     1,    -1,    -1,     0,    -1,    -2,     0,    -3,    -3,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     1,     2,     2,     2,     1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0),
		    46 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     2,     2,     1,     1,     0,     1,     1,     0,     0,     0,     0,     0,     2,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,     1,     1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     1,     1,     0,     2,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     0,     1,     1,     1,     1,     1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     1,    -1,    -1,    -1,     0,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,    -1,    -1,    -2,    -1,    -1,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,     0,     0,     1,     0,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     1,     1,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     1,     1,     0,    -1,     0,     0,     1,     1,     1,     0,    -1,     0,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,     0,     1,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -2,    -2,     0,     1,     0,     0,     0,     0,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     1,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    47 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,    -2,     0,     0,     0,    -1,    -3,    -3,    -2,    -2,    -3,    -3,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -2,    -4,    -3,    -1,     1,     1,     0,    -1,    -2,     1,     1,     0,     1,     2,     1,     1,    -1,    -1,    -1,     0,     0,     1,     1,     1,     1,     0,     1,     0,    -1,    -3,    -3,    -3,    -2,    -1,     0,    -2,     0,     0,     1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     2,    -1,     0,     0,     0,     1,     1,    -1,    -2,    -2,    -2,    -1,    -2,    -2,    -2,    -1,    -1,     0,    -1,    -1,    -2,    -1,     1,     1,     0,    -2,    -1,    -1,     1,    -1,    -1,     0,     0,     2,     0,     0,    -1,    -2,    -1,    -1,    -2,     0,     0,     0,     0,     0,    -1,    -1,     2,     1,     2,     2,     0,    -2,     0,     0,     1,     0,     0,    -2,    -1,     1,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     1,     1,     1,     0,     1,     1,     0,    -1,     0,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     2,     1,     1,     1,     0,    -1,    -1,     0,     1,     0,     1,     0,     1,     0,    -1,     0,     2,     0,     0,     1,     1,     1,     1,    -1,     1,     1,     0,     0,     1,     2,     0,    -1,    -1,     1,     1,     0,     0,     0,     0,     1,     0,     2,     1,     2,     2,     0,     0,     1,     1,     1,     0,     0,    -2,     0,     0,     1,     0,     0,    -1,    -1,    -1,     1,     0,     0,     0,     1,     1,     1,    -2,     2,     2,     1,     0,     0,     1,     2,     1,     0,     2,     0,    -2,     1,     1,     1,     0,    -2,    -3,    -1,    -1,     0,    -1,     1,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     2,    -1,     1,     0,     1,     0,     1,     1,    -1,    -4,    -3,    -2,     0,     0,     1,     0,     1,     1,     0,     0,    -2,    -2,     0,     0,     0,     0,     0,     0,     1,     2,     0,     0,     1,     0,     0,    -1,    -5,    -6,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,    -1,    -2,    -3,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     0,     0,    -1,    -3,    -4,    -3,     0,    -1,     0,    -1,     0,    -1,    -1,     1,     1,     0,    -1,    -2,    -2,     0,    -2,     1,     0,     1,    -2,     0,     0,     0,     1,     0,    -3,    -4,    -2,    -1,     0,     0,     0,    -2,     0,    -1,    -1,     1,     1,     0,    -2,    -2,     0,     0,     0,     0,     1,     0,    -2,     0,     0,     1,     0,    -1,    -3,    -3,    -1,    -1,     1,     0,     0,     0,     1,    -1,     1,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,    -1,    -1,     1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -3,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,    -1,     2,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     1,     0,     1,    -1,    -1,     1,    -1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,     0,    -1,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,     1,     1,    -2,     1,     0,     0,     0,    -1,    -2,     1,     0,     0,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     1,     1,     1,     0,     2,     1,     1,     0,     0,     0,     0,     0,     0,    -2,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     2,     1,     0,    -1,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     1,     0,     0,     0,     1,     0,    -1,     0,     1,    -2,     0,     0,     2,     2,     2,     0,     0,     0,     0),
		    48 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     2,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,    -1,     1,     2,     3,     1,    -2,    -2,    -1,     1,     0,     0,     0,    -1,     0,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -2,    -2,    -1,    -2,     0,     1,     2,     1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     0,     2,     0,     0,     1,     0,    -1,    -1,     0,     1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,     0,     0,    -1,     1,     0,    -1,     0,     2,     1,     0,    -1,     0,     1,     1,     0,    -1,    -1,    -1,     1,     0,     0,     1,     0,     0,     0,    -1,    -2,    -3,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     1,     0,    -1,    -2,    -2,    -1,     0,     1,     1,     0,     1,     1,     0,     0,     0,     0,    -2,     0,    -1,     0,     0,    -1,     1,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -2,     0,     1,     0,     0,     1,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,     1,     2,     0,    -1,    -2,    -2,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     2,     1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,     1,     0,     1,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,     1,     0,     0,    -2,    -1,    -1,    -1,    -2,     0,     0,     1,     1,     1,     1,     0,    -2,    -2,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     1,    -1,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,    -2,    -3,     0,     0,     1,     1,    -1,    -1,    -2,     0,     0,    -1,     1,     1,     1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,     2,    -1,     0,     1,    -1,     1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,     2,    -1,     0,     1,    -1,     1,     1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -1,     0,     1,     1,     1,    -1,    -1,     0,    -2,     1,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -2,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -3,    -2,    -2,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,    -1,    -1,    -2,    -1,    -1,     1,    -1,     0,     0,     2,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     1,     2,     1,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    49 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -2,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -3,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -2,    -4,    -2,    -3,    -3,    -3,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -2,    -3,    -4,    -1,    -2,    -2,    -1,     0,     1,    -4,    -2,    -3,    -2,     0,     0,    -2,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,    -2,    -1,     0,    -1,     1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -3,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,    -3,    -6,    -3,     0,     0,     2,     0,     1,     0,     2,     0,     0,     0,     1,     1,     0,     1,     1,    -2,    -2,    -3,    -2,    -2,    -1,     0,    -1,    -2,    -2,    -4,    -5,     0,    -2,    -1,     0,     1,     1,     2,     0,     0,     1,     0,     1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -3,     0,     0,    -2,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,    -1,     0,     1,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -1,     0,    -1,    -3,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -2,    -2,    -1,     0,    -2,    -3,     0,     1,     0,    -1,    -1,    -1,     1,     0,     1,     0,    -1,    -1,    -1,     0,     1,     0,     1,     1,     0,     1,     0,    -1,     3,    -2,    -2,     0,    -4,     1,     0,     1,     0,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,    -1,     0,     2,     0,     0,     1,     1,     2,    -1,     0,     3,    -2,    -2,     0,    -1,     1,     1,     2,     1,     0,     1,     0,     2,     0,     1,    -2,    -2,     0,     0,     1,     2,     2,     2,     1,     1,     2,     2,    -2,    -5,    -3,    -1,     0,    -2,    -1,     0,     3,     2,     1,     2,     2,     1,     1,     0,     0,     0,     1,     1,     2,     0,     1,     1,     2,     1,     3,     1,    -4,    -2,    -2,     0,    -1,    -1,    -1,     1,     2,     2,     1,     1,     2,     1,     1,    -1,    -1,     1,     0,     0,     1,     0,     1,     2,     0,     1,     4,     0,    -6,    -4,     0,     0,     0,     0,    -3,     1,     2,     0,    -1,     1,     2,     1,     0,    -1,    -1,     0,    -1,     1,     1,     2,     1,     1,    -1,    -1,     0,    -1,    -5,    -3,     1,    -1,     0,     0,    -3,    -2,     0,    -1,     0,     0,     0,    -1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -1,    -1,    -4,    -2,     0,    -2,     0,     0,    -3,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,     1,     0,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -3,     0,    -1,    -1,     1,     0,    -3,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,     0,     0,     1,     0,    -2,     0,     0,    -3,    -6,    -1,    -2,    -1,     0,     0,    -2,     2,    -1,    -2,    -2,    -2,    -1,    -2,    -1,    -1,    -2,    -4,    -1,     0,    -1,    -1,     0,     1,     0,    -1,     1,    -1,    -3,     0,    -1,     0,     0,     0,    -3,     2,    -1,     2,    -1,    -4,    -3,    -2,    -2,     0,    -2,    -2,     0,    -1,     0,     0,    -1,     1,    -2,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,    -3,     2,     1,     2,    -1,    -2,    -2,    -2,    -2,    -2,    -2,     0,    -2,    -1,     0,    -1,    -2,    -1,    -2,    -1,    -1,    -2,    -1,     1,    -5,     0,     0,     0,    -3,     2,    -1,    -1,     0,     1,     1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,    -2,     0,    -1,    -3,    -1,     0,     0,    -2,     1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,     1,    -1,     1,    -1,     0,     0,     1,     0,    -1,    -2,     0,     0,    -1,     0,     1,    -1,     0,     1,     2,     0,    -1,    -1,     0,     0,     0,     1,    -1,     2,     1,    -2,    -3,    -1,    -1,    -2,    -1,     0,     0,     2,     0,     1,     1,     1,     1,     2,     3,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     2,     0,     1,     2,     3,     1,     2,     2,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     1,     0,     1,     1,     0,     1,     0,    -1,     1,     1,     1,    -2,    -1,     1,     0,    -2,     1,    -1,     0,     0,     0,     0),
		    50 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -1,     0,     0,     1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     1,     0,     1,     1,     1,     1,     0,     0,     0,    -1,     0,     1,     1,     0,    -1,    -2,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,    -2,     0,     0,     1,     0,     1,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,    -1,    -1,     2,     1,    -2,    -2,     0,     0,     0,    -1,     0,    -1,     1,     1,     0,     0,     1,     1,     0,     0,     0,     1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     1,     1,    -1,    -1,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,     0,     0,     2,     1,     1,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     1,     1,     2,     1,     1,     0,     2,    -2,    -2,     0,     0,     0,     0,    -1,    -2,     0,     0,     0,     1,     0,     1,     0,    -2,    -1,     0,     0,    -1,     1,     1,     0,    -1,    -1,     2,     0,     2,    -1,    -1,     0,     0,     1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     1,    -2,    -2,    -2,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,     0,    -1,    -1,    -1,     0,     1,     0,     0,     1,     0,     0,     0,     2,     0,    -1,    -3,    -3,    -4,    -3,    -2,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     2,     1,     1,     1,     0,    -1,    -4,    -3,    -3,    -1,    -2,    -3,    -2,    -1,     0,    -1,     0,    -1,     1,     2,     0,    -1,     0,     0,     0,     0,    -2,     1,     1,     2,     0,     0,     1,     1,    -2,    -4,    -2,    -1,    -1,    -2,    -2,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -2,     1,     1,     0,     2,    -1,     0,     0,    -1,    -1,    -2,     0,    -1,    -3,    -2,    -2,    -2,     1,     2,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,     1,     2,     1,     1,    -1,    -3,    -4,    -2,    -3,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,     1,    -1,     1,     2,     1,     0,     0,    -1,     0,     0,    -1,    -2,    -3,    -3,    -1,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,    -1,     0,     1,    -1,     0,     1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     2,     2,    -1,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     1,     0,     0,     1,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     2,     0,     1,     0,    -1,     0,    -1,     0,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,     1,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     1,     2,     0,     1,     1,    -1,     1,     0,     1,     1,     1,    -1,    -2,    -2,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -3,    -3,    -4,    -2,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -2,    -1,    -2,    -2,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0),
		    51 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,    -1,     0,     2,     0,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     3,     2,     0,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -1,     0,     2,     2,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     2,     3,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     1,     1,     0,    -1,    -2,     1,     0,     1,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     2,     1,     0,     0,     0,    -1,    -3,    -3,    -1,     0,    -1,     1,     0,     0,     1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,    -3,    -3,    -2,     0,     0,     2,     1,    -1,     0,    -2,    -1,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -1,    -4,    -2,     0,     1,     1,     2,     0,     0,    -1,    -2,    -1,    -3,    -2,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -4,    -2,     0,     0,     0,     1,     2,     1,    -2,    -1,    -1,    -3,    -1,    -1,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,     1,     0,    -2,     0,     2,     2,    -1,    -2,     0,     0,    -1,     0,     1,     0,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,    -1,     0,    -2,    -1,    -1,    -2,     1,     0,    -1,     1,     1,     0,    -1,    -2,    -1,     0,    -1,    -2,     0,     1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,     0,     1,    -1,     0,     2,     0,     0,    -1,    -2,    -1,     1,     0,     1,     1,    -1,    -1,    -1,     2,     0,     0,    -2,     1,     0,     0,    -1,    -1,    -1,     1,     0,     0,     0,     0,     1,    -1,     0,    -2,    -2,    -1,     2,     0,     0,     1,    -1,     0,     0,     2,     0,     0,    -2,     0,     0,     0,     0,     0,     2,     1,    -2,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,     1,     2,    -1,    -1,    -2,    -2,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,    -1,    -1,    -2,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,    -2,     0,     0,     0,     2,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,    -1,    -1,     2,     1,     2,     1,    -2,     0,     0,     1,    -1,     1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,     1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -1,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -3,    -1,    -1,     2,     1,     0,     0,     0,     1,    -2,     1,     0,    -2,    -2,    -2,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,    -2,    -2,    -1,     0,     1,     2,     1,     0,    -1,    -1,    -3,    -1,    -1,    -2,    -1,    -1,     1,     1,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,     1,     0,     1,     1,     0,     0,    -1,    -1,     0,    -2,    -3,    -1,     0,     0,     1,     0,     1,     0,     0,    -1,    -1,     0,    -1,    -3,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,     1,     0,     1,    -1,    -2,    -2,    -1,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     1,     0,     1,     0,    -2,    -1,    -2,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,     0,     2,     0,     1,     0,     0,     0,     0,     0,     2,     1,     0,     1,    -1,     0,    -1,    -1,     0,     2,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     2,     0,    -2,    -1,    -2,    -3,    -1,    -2,    -1,    -1,    -1,    -2,     0,    -1,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -4,    -3,    -2,    -2,    -1,    -2,    -2,    -3,    -2,    -2,    -4,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    52 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     2,     2,     1,     1,    -1,     0,    -1,    -2,    -2,     0,     1,     0,     1,    -1,     0,     1,     1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,    -1,     1,     1,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,     1,    -1,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     1,    -1,     1,    -1,     0,     1,    -1,    -1,    -2,    -2,     1,    -2,    -1,     0,     0,     0,    -1,     0,    -2,    -2,    -3,    -1,     0,     1,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -2,     2,    -1,     0,     0,     0,     0,     2,     1,    -2,    -1,    -1,     1,     1,     1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     2,     2,     1,     0,     0,     0,     0,     0,     1,     0,     1,     0,     1,     1,     1,     0,     1,    -1,    -1,     2,     0,    -1,    -1,    -1,    -1,    -1,     2,     0,     2,     1,     1,    -1,     0,    -1,     1,     0,     0,     0,    -1,     0,     0,     1,     1,     0,     1,    -1,     0,     1,     1,    -3,    -2,    -1,    -1,     0,    -1,     1,     0,    -1,     0,    -1,    -1,     0,     1,    -1,     0,     1,    -2,     0,     0,     1,     0,     0,     1,     0,    -1,    -1,     1,    -3,    -2,    -1,     0,     0,     0,     0,     1,    -2,     2,     1,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,     1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,     1,     0,    -1,    -1,    -3,     0,    -1,    -2,    -2,    -2,     0,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,    -2,     0,     0,    -2,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -2,    -3,    -1,     0,     0,    -2,     0,    -1,     0,     0,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -3,    -2,    -4,    -2,    -2,    -2,    -3,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     1,     1,    -1,     0,    -1,    -1,     0,    -2,    -3,    -3,    -3,    -5,    -3,    -2,    -2,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -2,     0,    -2,     0,     0,     2,     1,     0,    -1,     0,    -1,    -3,    -2,    -1,    -2,     0,     0,    -1,     1,     0,     1,     0,    -2,     0,     0,    -2,    -2,    -2,    -1,    -2,    -1,     1,    -1,     2,     3,     0,     0,    -1,    -2,    -3,    -1,    -1,    -1,    -1,     1,     1,     1,    -1,     0,     1,    -1,    -1,     0,    -1,    -2,    -1,    -1,     1,    -1,     1,     2,     2,     2,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,     2,     1,     0,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,     3,     2,     1,     0,     0,     0,    -3,    -1,    -1,     1,     1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     1,    -1,    -1,    -2,     1,     1,     1,     2,     4,     0,     2,     0,    -1,     1,    -1,    -2,    -1,     1,     1,    -1,    -1,     1,     0,     0,     2,     2,     1,     1,     0,     0,    -1,     0,     1,     1,     1,     0,     1,     1,     2,     0,     0,     1,     0,     0,    -1,     3,     1,     1,     1,     2,     2,     1,     3,     1,     1,     2,     0,     0,     0,     2,     2,     1,     1,     0,     1,     1,     0,     0,     1,     1,     2,     0,     0,     1,     1,     0,     1,     1,     1,     0,     2,     2,     1,     1,     1,     1,     1,     1,     1,     1,     3,     1,     1,     1,     0,     0,     0,     0,     0,     0,     2,     2,     1,     0,     1,     0,     0,     0,     0,     1,     1,    -1,    -1,     0,    -1,     0,     1,     2,     3,     2,     0,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     2,     1,     1,     1,     1,     2,     2,     1,     0,     0,    -1,    -1,    -1,     0,     1,     2,     3,     2,     2,     0,    -1,     0,     0,     0,    -2,    -1,     0,    -1,     0,     1,     2,    -1,     0,     0,     1,    -1,     1,     0,    -2,     0,     0,     0,    -2,    -1,     0,     2,     3,     2,     1,     0,     0,     0,    -1,     0,    -1,    -3,     1,     0,    -2,    -3,    -4,    -1,    -1,     0,     1,     1,    -1,     0,    -2,    -3,     0,     0,    -2,    -1,     1,     2,     1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -2,    -4,    -3,    -2,    -2,    -2,    -1,    -3,    -3,    -2,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0),
		    53 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     1,     1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     1,     1,     1,     1,     0,    -1,     0,     1,     1,    -1,     0,    -1,     0,    -2,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -2,     0,    -1,    -1,    -2,    -1,     0,    -1,    -1,     1,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     2,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -2,    -1,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     1,     1,    -1,    -3,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     1,    -2,    -2,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,     1,     2,     1,    -2,    -4,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -1,     1,     1,     2,     1,     1,    -1,    -1,    -1,    -1,    -1,     1,     1,     1,    -2,    -4,    -2,    -2,     0,     0,    -2,    -1,     1,     0,     0,     2,     0,     3,     1,     1,     1,     0,     0,     0,    -1,    -2,     0,     1,     1,     1,     0,     1,    -1,    -4,     0,    -1,     0,     0,    -2,    -1,     2,     2,     2,     0,     1,     1,     2,     1,    -1,    -3,    -3,    -2,     1,     1,     1,     1,     1,     2,     0,     0,     0,    -2,    -2,     0,     0,     0,    -2,    -1,     2,     1,     1,     0,     1,    -2,    -1,    -2,    -4,    -3,    -1,     1,     2,     1,     0,     1,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,    -1,    -3,     1,    -2,    -1,    -1,    -1,    -2,    -4,    -4,    -3,    -1,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,    -2,    -2,     1,    -1,    -1,     0,    -1,     0,     0,    -1,    -2,    -2,    -3,    -3,    -3,    -2,    -1,    -1,     1,     1,     1,     0,     0,     0,    -2,    -1,    -1,    -1,    -2,     0,     2,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -3,    -3,    -3,     0,     1,    -1,     1,     2,     3,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,     2,    -1,     1,     0,     0,     0,     1,     2,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -3,     0,     0,    -1,    -1,     1,     1,    -1,     0,     0,     2,     0,    -1,     1,    -2,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -4,    -5,    -6,    -5,    -3,    -2,     1,     0,    -1,     1,     1,     2,     1,    -1,     0,    -2,     0,     0,    -1,     0,     2,     0,     2,     0,    -1,     0,     0,    -2,    -2,    -3,    -4,    -3,    -2,    -2,     0,     1,     1,     1,     0,     0,     1,     0,    -3,    -1,     0,    -1,     0,    -1,    -1,    -1,     1,     1,     0,     0,    -1,     1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,    -1,     1,     0,    -1,     0,     0,    -1,     0,     1,     1,     1,     1,     0,     1,     1,     2,     1,     0,    -1,    -2,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,    -1,     0,     0,     1,     0,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     1,     1,     1,     1,     0,    -1,     0,     0,    -2,    -1,    -1,     0,    -1,     1,     0,     1,     1,     0,     0,     1,    -2,    -1,     1,     1,     0,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,     0,     1,     0,     0,     1,     0,     0,    -1,     1,     1,    -1,    -2,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -2,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -2,    -3,    -3,    -2,    -1,    -1,    -1,    -1,    -3,    -3,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0),
		    54 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     1,     2,     1,    -1,    -2,    -3,    -2,    -2,    -1,    -2,    -3,    -3,    -2,    -1,    -1,     0,     3,     2,     1,    -2,     0,     0,     0,    -1,     0,    -1,     0,    -1,     1,     3,     1,    -2,    -3,    -2,    -1,     3,     2,     1,    -1,    -3,    -4,    -1,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,     0,    -1,     1,     2,    -1,     1,     1,    -1,    -3,    -4,    -1,     0,     0,     1,     1,     0,    -3,    -5,    -5,    -1,     2,     2,     1,    -3,     1,    -2,     0,    -1,     0,    -1,     1,     1,     1,     1,     0,    -1,    -2,    -1,    -2,     0,     1,     1,     1,     1,    -4,    -6,    -3,     1,     2,     3,     0,    -3,     0,    -2,    -1,    -1,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,    -2,    -2,     0,     1,     2,    -1,    -3,    -5,    -3,     0,     1,     1,     0,     0,    -1,     1,    -2,     0,     0,     0,    -2,     0,     0,     1,     2,     0,    -1,    -1,    -2,    -1,     0,     2,     1,     0,    -3,    -3,    -1,     1,     1,     0,     0,     0,    -1,     1,    -1,     0,    -1,    -1,    -2,    -1,     0,     0,     0,    -2,     1,     0,    -2,     1,     0,     2,     0,     0,    -2,    -2,     0,     1,     0,     0,    -1,     0,     1,     0,    -1,     0,     0,    -1,    -1,    -1,     1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,    -1,    -3,    -1,     1,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     1,     0,     0,    -1,     0,    -1,    -2,    -2,     0,     0,    -1,    -2,    -1,     0,     0,     1,     0,     1,     2,     0,    -1,     1,    -1,    -1,     1,     0,     0,     1,     0,     0,     0,     0,    -1,    -2,    -2,     0,     0,     0,    -1,    -2,    -1,     0,     1,     0,     0,     1,     1,     0,     0,     1,     1,    -1,     0,     1,    -1,     0,     0,     1,     1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -2,     0,     0,     1,     2,     1,     1,     1,     1,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -2,    -1,     1,     1,     2,     1,     0,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     1,    -1,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     1,     1,     0,    -1,    -1,    -1,     0,    -2,    -2,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,     2,     1,    -3,    -2,    -1,    -1,     0,    -3,    -2,    -1,    -2,     0,     0,    -1,    -1,     1,    -1,    -2,    -2,    -2,    -2,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,    -1,     1,     0,    -1,     0,     1,    -1,    -3,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -2,     0,     1,     0,     0,     0,    -2,     0,    -1,     0,    -1,     0,     0,    -2,     0,    -1,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     1,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     1,     0,     2,     1,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,     1,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -2,    -2,     1,     1,     0,     0,     0,     2,     1,    -1,     0,     0,    -2,     0,     0,     1,     1,     0,     1,     1,     0,     2,     0,     0,     0,     0,     0,     0,    -1,    -3,     0,     0,     0,     0,     1,     1,    -2,    -3,    -1,     0,    -2,     0,    -1,    -2,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -1,    -2,    -2,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,     0,    -1,    -2,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0),
		    55 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -3,    -4,    -2,     1,     1,     1,     1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -4,     1,     1,     0,     0,     0,    -1,    -2,    -1,     0,     1,     2,     0,     1,     0,    -1,    -1,     1,     2,     0,     0,    -1,    -1,     0,    -2,     0,     0,     0,     0,     0,     1,     0,     1,    -1,     0,    -1,    -2,    -1,     1,    -1,    -1,     0,    -1,    -1,     2,     2,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     0,     2,     2,    -1,     1,     1,     0,    -1,    -3,    -1,     0,     0,     0,     1,     0,     2,     1,     0,     0,     0,     0,    -2,    -2,    -1,     0,     1,     1,     0,     0,     2,     2,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     1,     2,     2,     2,     0,     0,     0,    -1,     0,    -3,    -3,    -1,     1,     2,     2,     1,     2,     1,     0,     0,     1,     0,     1,     0,    -2,     0,     0,     0,     0,     0,     1,     1,    -1,     1,     0,    -1,    -2,    -4,    -2,     1,     0,    -1,     0,     1,     1,     0,     0,     0,     1,     1,     0,     1,    -1,    -3,    -1,    -1,     0,     0,     3,     1,    -2,     1,     0,     0,    -2,    -3,    -1,     1,     1,    -2,     0,    -1,     0,     2,     1,     2,     3,     2,     0,    -1,    -3,    -3,    -3,    -1,     1,     0,     2,     2,    -1,    -1,     0,     0,    -2,    -5,     2,     2,     1,     1,    -1,    -1,     1,     2,     3,     2,     2,     2,     0,    -3,    -1,    -2,    -2,    -1,    -4,    -3,     1,     2,     2,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,    -1,    -1,     0,     1,     1,     1,     1,     2,     1,     0,    -1,    -2,    -1,    -1,    -4,    -4,     0,     0,     1,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,     0,    -3,    -2,    -4,    -2,     2,    -2,     0,     0,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,    -1,    -2,    -4,    -3,     0,    -1,     0,     0,     0,     0,    -2,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     1,     0,    -1,     0,     1,     0,     0,     2,     0,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     2,     1,    -2,    -2,    -2,     0,    -1,    -2,     2,     0,     1,    -3,    -4,    -2,    -2,    -1,     2,     0,     0,     0,    -1,     0,    -1,     0,     1,    -1,    -1,     0,     1,    -1,    -4,    -2,    -2,     0,     0,    -3,     3,     1,     0,    -1,    -3,    -2,    -2,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     1,     0,     0,     0,     1,    -2,    -4,    -3,    -3,     0,     0,    -2,     3,     3,     2,     0,    -2,    -3,    -4,    -1,    -2,    -1,    -2,     0,     0,     1,     1,     0,    -1,     1,     1,     1,     2,     0,    -1,    -3,    -1,     0,    -1,     2,     0,     3,     2,     1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     1,    -1,     1,     2,     0,     2,     0,     1,     2,     2,     1,    -2,    -2,     0,    -1,     1,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,     1,     1,     0,    -1,     1,     0,     2,     1,     1,     2,    -2,     0,     0,     0,    -2,    -3,     0,     1,    -1,    -1,     1,     1,     0,    -1,    -1,     0,     1,     2,     1,     1,     1,     1,     0,     1,     0,     2,     1,     3,     1,     0,     0,     0,    -2,    -1,    -2,    -2,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     3,     3,     3,     2,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -2,     0,     0,     0,    -1,     1,     1,     0,     0,     0,     1,     1,     0,     1,    -1,     2,     2,     2,     2,     0,     0,     0,    -2,     0,    -1,    -1,    -1,     1,     1,     2,     2,     1,     0,    -1,    -2,     0,     0,     2,     1,     2,     1,    -1,     0,     0,     2,    -1,    -1,     0,     0,     0,     0,     1,    -2,    -3,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,     0,     2,     2,     2,     1,     0,     2,     3,     2,     2,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -3,    -1,     0,     1,     0,     0,    -1,    -2,     1,     0,     1,     1,     2,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -3,    -2,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0),
		    56 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,     1,     0,     1,     0,     0,     0,     0,     0,     0,     2,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     2,     1,     1,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     1,     1,     2,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,    -1,    -3,    -1,    -1,     0,    -1,     1,     2,     1,     1,     0,     2,     1,     0,     0,     0,     0,     0,    -2,    -2,     1,     2,     1,     0,    -1,     1,     0,    -2,    -2,    -3,    -2,     0,     0,    -1,    -2,     0,     0,    -1,    -1,     0,     1,     1,     2,     2,     0,     0,    -1,    -2,     3,     1,     1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     2,     1,     0,     0,     0,     0,     2,     1,     1,     0,     2,     1,    -1,    -2,    -2,    -2,    -1,    -1,    -2,    -1,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,     2,     0,     0,     0,    -1,     2,     1,     0,     1,     1,     1,    -1,    -2,    -2,    -1,     0,    -2,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,     2,     0,     0,     0,    -1,     2,     0,     0,     1,     0,     0,    -1,    -2,    -3,     0,     0,    -2,     0,     1,     0,     1,     1,     0,    -1,     0,     0,    -1,     1,    -1,     0,     0,     0,    -1,     1,     0,    -1,     1,     0,    -1,    -3,    -3,    -3,    -1,     0,    -1,     1,     1,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     1,     1,     1,     2,     0,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,     1,     2,     0,     0,     0,    -1,    -2,    -2,    -1,     2,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     1,     1,     1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,    -1,    -2,     0,     1,     0,    -1,     0,     0,    -1,    -1,    -1,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     1,     1,     0,     0,     0,    -2,     0,     0,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     2,     0,     0,     1,    -1,    -1,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     1,     0,     0,     2,     0,     1,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     0,    -1,     1,     0,     0,     1,     0,     0,    -1,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,     1,     1,     1,     1,    -1,     0,    -1,    -2,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     1,    -1,     0,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    57 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -2,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -3,    -3,    -2,    -3,    -4,    -4,    -3,    -3,    -3,    -2,    -1,    -1,    -2,    -1,    -2,    -5,    -3,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -4,    -5,    -6,    -6,    -1,     0,     0,    -1,    -1,    -3,    -5,    -4,    -3,    -2,    -2,    -3,    -4,    -4,    -2,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -2,    -1,     0,     1,    -1,     1,     1,     1,     0,     0,    -1,    -2,    -3,    -4,    -4,    -3,    -3,    -6,    -4,    -4,     0,     0,     0,     0,    -1,    -1,    -1,     1,     1,     1,     0,     1,     2,     2,     0,     0,    -1,    -1,     1,    -1,     0,    -2,    -2,    -1,    -2,    -2,    -3,    -3,    -2,    -1,     0,     1,    -1,     0,     0,     2,     1,     1,     1,     1,     2,     0,     1,     1,     1,     0,     1,     1,     1,     1,    -1,     0,     0,    -1,    -2,    -4,    -3,    -2,    -1,     1,     0,     1,     0,     2,     0,     1,     0,    -1,     1,     1,    -1,    -2,    -1,     1,     1,     1,     1,     1,     1,     1,     0,     0,    -2,    -2,    -2,    -1,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     1,     1,     0,     0,     1,     0,     1,    -2,     0,     2,     3,     0,     1,     0,    -1,     1,    -2,     0,    -1,     0,     0,     0,     1,    -1,    -1,     0,     0,     1,     1,     2,     1,     1,     0,     1,     0,     0,     1,     2,     3,     0,     0,     0,    -1,     1,     1,    -1,    -1,     0,     1,     0,    -1,     0,     1,     0,     0,     1,     1,     1,     1,    -1,     0,     1,     1,     0,    -2,     0,     2,     0,     1,     1,     0,     1,     2,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,     1,     1,     1,     1,     0,     0,     0,     0,     1,     0,     1,     2,     3,     0,     0,     2,     0,     1,     2,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     1,     2,     0,    -1,     0,     1,     1,     0,     0,     1,    -1,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,     1,     0,     1,     0,    -1,     0,    -1,     0,    -3,    -3,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     1,     1,    -1,     0,     1,     1,     0,     0,    -1,    -2,    -3,    -3,     0,    -2,     0,     0,     0,    -1,     0,     1,    -1,    -1,    -1,     1,     1,     0,     1,     2,     1,     2,     1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -3,    -2,    -2,     0,     0,    -1,    -2,     1,     0,     0,    -1,    -1,    -2,    -1,    -1,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,    -2,    -1,    -2,     0,     0,     1,    -4,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     1,    -1,    -2,     0,     0,    -1,     1,     1,     0,     1,     0,    -3,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -2,     0,    -1,    -1,     0,     1,     1,     0,    -2,     0,     0,     0,     0,     0,     2,    -1,    -1,     1,    -3,    -2,    -1,     0,     0,    -1,    -1,    -3,    -2,    -2,    -1,    -2,    -1,    -2,    -2,    -1,     1,     0,    -1,     0,     0,    -2,     0,     0,     0,    -1,    -3,    -1,    -2,    -2,     0,     0,     0,    -1,    -2,    -3,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -2,    -1,    -1,     1,    -1,    -2,    -3,    -1,    -1,     0,     0,     0,    -1,    -2,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     1,     0,    -1,    -6,    -3,     0,    -1,     0,     0,     0,    -1,    -2,     0,     1,     0,     0,     1,     1,     0,     1,     2,     1,     2,     0,     1,     1,     0,     0,     1,     0,    -1,    -5,    -3,    -1,    -2,     0,     0,     0,     1,    -1,     2,     2,     2,     2,     2,     0,     1,     1,     2,     3,     3,     0,     2,     1,     0,     1,     1,     1,     0,    -4,    -2,    -2,    -2,     0,     0,     0,     0,     1,     1,     1,     1,     1,     1,     1,     2,     2,     2,     1,     1,    -1,     3,     1,     1,     1,     0,     1,     2,    -1,     0,    -2,    -1,     0,     0,     0,     0,    -1,    -1,    -2,     0,     1,     1,     2,     2,     2,     2,    -1,    -3,     0,     1,     0,     0,     2,     1,     1,     2,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     1,     1,     0,     0,    -2,     0,     1,    -1,     1,     1,     1,     0,     1,     1,     2,     0,     0,     0,     0),
		    58 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -3,    -1,     0,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -4,     0,     1,     1,     0,    -1,    -1,    -1,     1,    -1,    -2,     0,    -1,    -1,    -1,     1,     2,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -2,    -1,     1,     3,     2,     2,     1,     0,     0,     1,     1,     1,     2,     0,    -1,    -2,    -2,    -1,    -2,    -2,     0,     1,     0,     0,     0,    -2,    -2,    -2,    -2,     0,     3,     1,     1,     1,     2,     2,     1,     0,     0,     1,     2,     0,     2,     0,     0,     1,    -1,    -1,    -1,    -2,    -1,     0,     0,    -3,    -2,    -2,    -1,    -1,     1,    -1,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,     0,     0,     1,    -1,    -1,    -1,     0,     0,    -2,    -2,    -2,    -2,    -2,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     1,     0,     0,     0,     0,    -1,     0,    -1,     2,     1,    -2,    -2,     1,     1,    -1,    -2,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,    -1,     2,     1,     2,     2,    -1,     2,     2,     0,    -1,    -2,     1,     1,    -1,     0,     1,     1,     0,    -1,     0,     0,     0,     1,     0,     0,     1,     0,     0,     1,     1,     1,     1,     0,    -1,     2,    -3,     0,     0,    -3,    -2,     3,     1,    -1,     1,     1,     0,     1,     0,     0,     0,     1,    -2,    -2,     0,     0,     0,     0,     2,     1,     1,     1,    -2,     1,    -1,     0,     0,    -1,     0,     2,     2,     0,     1,     0,     0,     1,     0,    -1,    -1,     0,    -2,    -2,    -1,     0,     0,     1,     1,     1,     1,     2,     1,     2,    -1,     0,     0,    -2,     0,     2,     4,     0,     0,     1,     1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,     1,     1,     2,     0,     1,    -1,     1,    -2,     0,     0,    -1,     0,     1,     2,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,    -1,    -1,     1,     0,     2,     0,    -1,    -1,     1,     0,     0,    -1,     0,    -1,    -2,     0,     1,    -2,     1,    -3,    -2,     0,    -1,    -1,     0,     0,    -1,    -2,     0,    -1,    -2,     1,     0,    -1,    -2,     0,    -1,    -1,     0,     0,    -1,     1,    -4,    -1,    -1,    -1,     1,    -1,    -1,     0,    -2,     0,     1,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -2,    -3,    -1,    -3,    -2,     0,     0,    -1,     1,    -3,    -1,    -2,    -3,    -2,     0,    -2,    -1,     0,     1,     0,    -1,    -1,    -2,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -3,    -2,     0,     0,    -1,    -2,    -1,    -2,    -2,    -2,     0,    -1,    -1,    -2,     0,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -3,    -1,    -2,     0,     0,    -1,    -3,     0,    -2,     0,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -3,     0,     0,     0,     1,     0,    -1,     0,     0,     0,    -3,    -1,    -2,     0,     0,    -2,    -3,    -1,    -2,    -1,     1,     2,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,     1,     1,    -1,     0,     1,     2,    -4,    -3,    -2,     0,     0,    -1,    -2,    -2,     0,     1,     0,     2,    -1,     2,     0,     1,     0,    -1,     0,     1,     1,     0,     0,     1,     1,     1,     3,     1,    -5,    -3,     0,    -1,    -1,    -1,    -1,    -2,     0,     2,     0,     1,     2,     1,     1,     0,     1,     1,     2,     0,     2,    -2,     1,     0,     0,     2,     2,    -1,    -3,    -2,     0,    -1,    -1,    -1,    -1,     1,     2,     1,     2,     2,     2,     2,     2,     1,     2,     3,     3,     0,     0,     1,    -1,     0,     0,     2,     1,    -1,     0,    -2,     0,     0,     0,     0,    -1,     2,     0,     1,     0,     1,     1,     0,     0,     2,     2,     2,     2,     2,     2,     2,     3,     1,    -1,     3,     1,    -1,     0,    -2,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     1,     1,     1,     0,     2,     1,     1,     1,     3,     0,     0,     0,     0,    -1,     0,     0,    -1,    -3,    -2,     0,     0,     0,    -1,     0,    -4,    -3,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,     1,     1,     0,    -1,     1,     0,    -2,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -3,    -1,     0,     0,    -1,    -1,     1,     0,    -2,    -5,    -2,    -1,    -1,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0),
		    59 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     1,     0,     1,     1,     1,     0,    -1,     1,     0,    -3,    -3,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,    -1,     0,     1,     0,     1,    -1,    -2,    -1,    -2,    -3,    -4,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     1,     0,    -2,     1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -2,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     1,     1,     0,     1,     1,    -1,    -1,     0,     0,    -1,    -2,     1,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -2,     1,     1,     1,     0,     0,    -3,    -2,     0,     2,     0,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,    -2,    -1,     1,    -1,    -2,     1,     1,     1,     0,    -1,     0,     1,     3,     0,     0,     0,     1,     0,     0,    -2,    -3,    -2,    -2,    -1,    -1,     0,    -1,     0,    -1,    -1,     1,    -1,     1,     1,     0,     0,     1,     1,     0,     1,     2,    -1,    -2,     0,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     3,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     2,     0,    -1,    -1,     1,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     1,    -1,    -1,     0,     0,    -1,     1,     0,    -1,    -2,    -1,     0,     1,     0,     0,     0,    -3,    -3,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -3,     0,     0,    -1,     0,     3,     1,     0,     0,    -1,    -1,    -1,     0,    -1,    -4,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -3,     0,    -2,    -1,     1,     1,     1,     0,     0,    -1,    -2,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -1,     1,    -1,     0,    -1,     0,     0,    -1,     0,    -1,    -2,     0,    -1,    -2,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -2,    -2,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,    -1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -3,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,     1,     0,     0,     1,     1,     1,     1,     0,     0,     1,     0,     0,     1,     0,     1,     0,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     1,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     1,    -1,    -2,    -2,     0,     0,     1,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -2,    -1,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,    -1,    -1,     1,     0,     1,     1,     0,     3,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     0,     0,    -1,    -1,     2,     2,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     0),
		    60 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -2,     2,     2,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     2,    -1,    -1,     0,     0,    -1,    -2,    -2,    -2,    -4,    -2,    -1,     0,    -2,    -1,    -1,    -1,    -1,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     2,     1,    -2,    -2,    -2,    -2,    -1,    -1,    -2,    -3,    -2,    -2,    -2,     1,     1,     0,    -1,    -2,    -2,    -3,    -2,    -1,    -1,    -2,     0,     0,     0,     0,    -1,    -1,    -4,    -1,    -2,     0,     2,     0,     0,    -2,     0,    -1,     1,     2,     1,     0,     0,    -1,    -1,    -1,    -1,    -3,    -4,    -2,     0,     0,     0,    -1,    -1,    -1,    -2,     1,     0,     0,     2,     2,     1,     0,     0,     1,     1,     1,     1,     1,     0,     0,     0,    -1,    -1,    -2,    -4,    -1,     0,     0,     0,    -1,     0,    -3,     1,     2,     1,     1,     1,     2,     1,     0,     0,     1,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -3,    -2,    -4,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,    -1,     1,     0,     0,     0,     1,    -1,    -2,    -1,     0,    -1,    -1,     0,    -1,     0,     0,    -2,    -1,    -2,     0,     3,    -2,     0,    -2,    -2,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -2,     0,     0,     1,     0,    -1,    -1,     0,     0,     1,    -2,    -4,    -2,     0,     0,    -1,     1,     0,     0,     0,    -1,    -1,     0,     1,    -1,     1,     1,     0,     0,     1,     1,     1,     0,     1,     1,     0,     0,     1,     0,    -3,    -1,     0,     0,     0,     1,     1,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     1,     3,     2,     2,     2,     0,     1,     1,    -1,     0,     1,     0,    -1,    -2,     0,     0,     3,    -2,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     1,     3,     1,     2,     4,     3,     3,     2,     1,     1,     1,     1,     2,    -2,    -2,     0,     0,     0,    -2,    -1,     1,    -2,    -2,    -2,    -2,     0,    -1,     0,     2,     3,     2,     2,     1,     1,     1,     1,    -1,     0,     0,     0,     1,    -1,    -2,    -1,     0,     0,     0,    -1,     1,     0,     0,    -1,     0,    -1,    -1,     1,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     1,     1,    -3,    -1,     0,     0,     0,    -2,    -1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -2,    -3,    -3,    -1,     1,     0,     1,     2,     2,     1,     2,     2,    -2,     0,     0,     0,    -2,    -2,     0,    -1,    -1,     1,     0,    -2,    -1,    -1,    -2,    -2,    -4,    -2,    -1,     0,    -1,     0,     1,     1,     0,     1,     2,     2,    -2,    -2,     0,     0,    -1,    -1,     1,    -1,    -2,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,     0,    -2,    -2,    -1,     1,     1,     0,    -1,    -1,     0,    -1,    -3,    -1,     0,     0,    -1,     0,     0,     0,    -1,     1,     0,     0,     1,     1,     0,     1,    -1,    -1,    -1,     0,     0,     1,     0,    -2,     0,    -1,     0,    -2,    -2,     1,     0,     0,    -1,    -1,     1,     1,     1,     0,     0,     1,     1,     1,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,     1,    -2,    -2,    -2,    -1,     0,     0,     0,    -1,     0,     2,     1,     2,     1,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,     2,    -1,    -1,     0,     1,     0,    -3,     0,     0,     0,     1,    -1,    -1,     2,     1,     1,     1,     1,     2,     0,     1,     2,     1,     0,     1,     0,     1,     0,     0,    -1,    -2,    -1,     0,    -1,    -4,     0,     0,     0,     0,    -2,    -1,     0,     0,     2,     2,     2,     1,     1,     0,     1,     0,     0,     1,     1,     0,     1,     0,    -1,    -1,     0,     0,    -2,    -2,     4,     0,     0,     0,    -1,    -1,    -3,    -1,     0,     2,     2,     0,     2,     1,     0,    -1,     1,     1,     1,     1,    -1,     0,    -2,    -2,    -1,     0,    -1,    -1,     2,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,     0,     2,     1,     1,    -1,     1,     0,     0,     1,     1,     2,     0,    -2,    -3,    -2,    -2,    -1,    -2,    -2,    -2,     0,     0,     0,    -1,    -1,     1,     1,    -2,    -1,    -1,     0,    -1,    -3,    -2,    -2,    -2,     1,     0,     0,    -1,    -2,    -1,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -4,    -2,    -2,    -3,    -2,    -2,    -1,    -2,    -2,    -5,    -4,    -4,    -4,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -2,    -1,    -2,    -2,    -2,    -1,    -1,    -2,    -3,    -3,    -2,    -2,    -3,    -2,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0),
		    61 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     3,     2,     0,     0,     0,     1,     0,     0,     0,     0,    -2,    -5,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,     3,     1,     0,    -1,     0,     0,     0,     0,     2,     2,     1,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -3,    -3,     2,     1,     1,     1,     1,     1,     0,     1,     1,    -1,    -2,    -2,    -2,    -1,     0,     0,     2,     2,     1,     0,    -1,    -1,    -4,    -2,    -3,    -3,    -3,    -2,     0,     1,     0,    -1,    -2,    -1,     0,     1,     1,     0,    -1,    -2,    -2,    -2,     0,     0,    -1,     1,     2,    -1,     2,     2,    -1,    -3,    -4,    -4,    -2,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,     0,     0,    -2,    -2,    -1,    -1,     0,    -2,    -2,     0,    -1,     2,     2,     2,    -3,    -3,    -6,    -3,    -2,    -1,     0,     0,     1,     1,     0,     1,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -2,    -2,     1,    -1,     1,     1,     0,    -2,    -2,    -2,    -3,    -3,    -2,     0,     1,     1,     1,     0,     1,     1,     0,    -1,    -1,    -3,    -1,    -2,     0,     0,     0,    -2,     0,    -1,    -1,     1,     2,     1,     0,    -1,    -3,    -1,    -2,     0,     1,     2,     1,     1,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,     1,    -2,    -1,    -1,    -2,     0,     2,    -1,     0,     1,     0,    -1,    -2,     0,     1,     1,     1,     0,    -1,    -2,    -3,     0,     0,    -1,     0,     0,     2,     0,     0,     0,     1,     0,     1,     1,    -2,    -3,    -1,     1,    -1,    -3,     0,     0,     1,     1,     0,    -1,    -3,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,     1,     0,     2,     2,    -1,    -1,     0,     0,    -1,    -1,     1,     1,     0,     1,     1,    -2,    -2,    -1,     2,     0,    -1,    -1,     1,     0,     1,     0,     0,     0,     1,     1,     1,     1,     0,     1,     1,    -1,    -1,    -1,     0,     1,     0,     0,     1,    -3,    -4,    -2,     1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     2,    -1,    -1,    -3,     1,     0,     0,    -1,    -1,     1,     1,    -1,     1,    -1,     0,    -2,    -1,     2,     1,     0,    -1,     2,     2,     0,     0,     0,     0,     2,     1,    -2,     0,     0,     1,     0,     0,     1,     0,     0,    -1,    -1,     1,     1,    -3,    -3,    -1,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,     1,     0,     0,     0,     0,    -2,     0,     0,    -2,     0,    -1,     1,     0,     0,     1,     0,    -2,    -3,    -2,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -2,     1,     0,     0,    -1,    -1,    -1,    -1,     1,     0,     1,     0,    -1,     0,    -2,    -2,    -2,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,     1,     0,    -1,    -2,    -2,    -1,    -2,    -2,     0,     0,     1,     0,     1,     0,     1,     0,     0,     1,     1,     0,    -2,    -1,    -1,     0,     1,     0,     1,     0,     1,     0,     0,    -2,    -1,    -1,    -2,    -1,     0,    -1,     1,     1,     2,     0,     1,     0,     0,     1,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,     0,    -2,     0,    -1,     1,    -1,     0,     1,     2,     2,     0,     0,     1,     1,     1,     1,     0,     1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -2,     0,     1,     2,     1,     0,     1,     2,     1,     0,     0,     1,     1,     1,     1,     0,     1,     0,    -2,    -1,     0,    -1,    -1,     0,     0,     1,     2,     1,     0,     2,     1,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     2,     0,    -1,     0,     0,     1,     2,     1,     2,     1,     0,    -2,    -2,     0,    -1,     1,     2,     2,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     0,     0,     2,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -3,     0,     1,    -4,    -3,     0,     0,     1,    -1,    -2,    -3,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -3,    -3,    -1,    -1,    -3,    -3,    -1,    -1,     1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    62 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     3,     1,     0,    -1,    -1,    -2,    -4,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     2,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     1,     0,    -2,    -2,    -2,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     1,     3,     3,    -1,     0,     1,     2,     1,     2,     2,     1,     0,     0,     0,    -1,     0,     1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     2,     0,    -1,     1,     0,     1,     1,     0,     1,     1,     0,     0,     0,    -1,     1,     2,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     0,    -2,     1,     1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     1,     3,     1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,    -2,     0,     1,     0,     1,     0,     0,     1,     2,     1,     0,    -1,    -1,    -2,     0,     0,     1,    -2,    -2,    -2,     0,    -1,    -1,     1,     1,     0,     1,    -1,    -1,    -1,     0,     0,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     2,    -1,     1,     1,    -2,     0,     0,     0,     0,    -1,     0,    -3,    -5,     0,     1,     1,     0,     0,     0,     0,     0,     1,    -2,    -1,     1,    -1,     0,     0,     1,     1,     0,     0,    -1,     2,     1,    -1,    -1,    -1,    -2,    -4,    -2,    -1,     0,     0,    -1,     0,    -1,     0,    -2,     1,    -1,    -1,     1,     0,     0,     0,    -1,     1,     1,     0,     0,     0,     0,    -3,    -2,    -3,    -4,    -4,    -1,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,     2,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -3,    -3,    -3,    -3,    -2,    -3,    -1,     0,    -1,     1,     0,    -1,    -1,     0,     0,    -1,     1,     0,     1,     1,    -1,     0,     0,     1,     0,    -1,    -2,    -3,    -4,    -5,    -5,    -2,    -2,    -1,     1,    -1,    -1,     1,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -3,    -4,    -2,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     0,    -2,    -2,    -1,    -1,     0,     1,     1,     1,    -1,     1,     0,    -1,     0,    -1,    -2,    -1,    -2,     0,     0,    -1,     0,     1,     1,     2,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -1,     1,     0,     1,     0,     0,     0,    -2,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,    -1,     2,     1,     1,     0,     0,     0,     0,    -1,     0,    -2,    -1,     0,     0,     0,     1,     1,     1,     0,    -1,    -1,    -2,    -3,    -2,     0,     0,    -2,    -2,    -1,     1,     0,     1,     0,     0,    -1,     1,     1,     0,     0,     0,     1,     1,     0,     0,     2,     0,     0,    -2,    -2,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     3,    -1,     2,     0,     0,     0,     1,     1,     0,     0,     1,     2,     0,     1,     1,     2,     1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,    -2,     1,     1,     2,     2,     0,     0,     1,     2,     2,     2,    -1,     1,     0,     0,     0,     1,     1,     1,     0,     1,     0,     1,    -2,     0,     0,     1,     0,     0,     1,     1,     2,     0,     0,     1,     2,     1,     1,     1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     1,    -1,     0,     2,     0,     1,     1,     1,     3,     3,     1,     0,     0,     0,     2,     1,     0,     0,     0,     0,     1,    -1,     1,     0,     0,     0,     1,     1,     0,    -2,    -1,     1,     1,     0,     1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     1,     0,     0,     2,     0,     0,     1,     0,    -1,     1,     2,     0,    -2,     1,     1,     0,     1,     1,     1,     1,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -4,    -3,    -1,     0,     0,     1,     1,     2,     0,    -1,     0,     1,     1,    -1,     1,     3,     2,     2,     1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -3,    -1,     0,    -1,     0,     2,     2,     1,     3,     0,    -3,     0,     1,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,    -2,    -1,    -3,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    63 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,     1,     1,    -1,    -2,    -2,     0,    -1,    -1,     0,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     2,     1,     0,    -1,     1,     1,     1,     2,     1,    -1,     0,    -1,    -1,     0,     0,    -3,    -4,    -2,    -1,     0,     0,     0,     0,    -1,     1,    -2,     0,     2,     1,     0,    -1,    -1,    -1,     0,     1,     2,     0,     0,    -2,    -1,     0,    -1,     1,     0,    -5,    -4,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,    -1,    -2,     0,     1,     1,     0,     1,     0,     1,     0,     0,     1,     1,     2,     1,     2,     1,    -4,    -1,     0,     0,     0,     1,     0,     1,     0,     1,     1,    -2,     0,     1,     2,     1,     1,    -1,    -1,    -1,     0,     1,     0,     2,     2,     0,     0,     1,    -3,    -2,    -1,     0,     0,     0,     1,     3,     1,     2,     1,     0,     0,     1,     1,     1,     0,     1,     1,    -2,     0,     0,     1,     0,     0,    -2,     0,     1,    -3,    -3,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,     1,     1,     1,    -1,     1,     2,     1,     1,    -1,    -1,    -1,    -4,    -3,    -1,     0,    -1,     0,    -1,     1,     1,     0,    -1,     0,    -1,    -1,     0,     0,     1,     1,     1,     1,     1,     1,     1,    -1,    -1,    -1,    -1,    -4,    -4,    -4,    -1,     0,    -2,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     1,     1,    -1,     0,     1,     2,     1,    -2,     0,    -3,    -2,     0,    -3,    -2,    -3,    -1,     0,    -1,    -2,     0,    -1,    -1,     0,     1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     3,     1,     0,     0,    -2,    -1,    -1,    -4,    -5,    -3,     0,     0,    -1,    -2,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,     1,     0,    -1,     0,     1,     2,     1,     2,     1,     0,     0,    -1,    -5,    -3,    -1,     0,     0,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     1,     0,     0,    -1,     2,     2,     0,     1,     1,     0,    -1,    -1,     0,    -3,    -2,    -1,     0,     1,     0,    -1,    -2,     0,     0,     0,     0,    -1,     0,     1,     0,     0,    -1,    -1,     0,     2,     1,     2,     1,     1,     0,     0,     1,    -3,    -2,     0,     0,     1,     0,     0,    -1,     2,     2,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     1,     1,     1,     1,     1,     0,     1,     0,     2,    -2,    -1,    -1,     0,     0,     0,     1,     0,     1,     2,     1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     1,     2,     1,     0,     2,     1,     0,    -1,     0,    -3,    -3,    -1,     0,     0,     0,     2,     0,     0,     2,     2,    -1,    -1,     0,     0,     1,     0,    -2,     0,     1,     1,     0,    -1,     0,     0,     0,    -1,    -3,    -3,    -1,     0,    -1,     0,     0,     2,     0,     0,     2,     1,     0,     0,     1,     0,     0,    -2,    -1,     1,     1,     0,    -1,     0,     0,     0,    -1,    -1,    -3,    -3,    -1,    -1,     0,    -1,     0,     0,     1,     1,     1,     2,     1,     1,     1,     0,    -2,    -2,    -1,     0,    -2,    -2,    -1,     0,     0,    -1,     1,     0,    -2,    -3,    -3,    -1,     0,    -1,    -1,     0,     0,     2,     1,     1,     0,     0,     1,     1,    -2,    -2,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -2,     2,     0,     0,    -2,    -1,     0,     0,     0,     1,     0,     0,     1,     1,     0,     0,     0,     1,     2,     0,    -2,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,    -2,    -1,     0,    -1,    -1,     1,     0,     0,     1,     1,    -1,     0,     0,     2,     2,     1,    -1,    -1,     1,     0,     0,     1,     0,     0,     0,     1,    -1,    -3,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,     1,     2,     1,     2,     1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,    -1,     2,     0,     0,     0,     1,     2,     2,     2,     0,     0,     1,     1,     1,     2,     1,    -1,    -1,     0,     0,     0,     0,    -3,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     1,     1,     1,     1,     2,     1,     0,     1,     0,     1,     1,     1,     1,     1,     1,     1,     0,    -1,    -4,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -2,     1,     1,     1,    -2,    -2,     0,     0,    -1,    -2,    -1,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    64 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -3,    -2,     0,    -1,    -2,    -1,     0,     0,     0,     1,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,    -1,    -1,     0,     2,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     1,     0,     1,    -2,    -3,    -4,    -4,    -1,     1,     1,    -2,    -2,    -1,    -1,     0,     1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,     1,     1,    -1,    -3,    -4,    -6,    -4,    -1,     0,     1,    -1,    -3,    -1,     0,     1,     2,    -1,    -2,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     1,     2,     1,    -2,    -5,    -7,    -2,     1,     1,     1,    -2,     0,     1,     2,     3,     1,    -2,    -2,    -1,    -2,    -1,    -1,     0,    -2,    -1,    -1,     1,     0,     0,     2,     1,    -1,    -6,    -4,    -1,     0,     2,     0,    -2,    -1,     0,     1,     0,     1,    -2,     0,    -2,    -2,     0,    -1,     0,    -2,    -1,     0,    -1,     1,     1,     1,     1,    -1,    -2,    -2,    -1,     0,     1,    -1,    -1,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,     0,     0,     0,     1,     1,     2,     1,     0,    -2,    -3,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,     1,     2,     1,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     1,    -1,    -2,     0,     0,     0,    -2,    -1,     0,     1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -2,    -2,     0,    -1,    -2,     0,     0,    -1,    -1,    -2,    -1,     1,     1,     0,     1,     1,     0,     0,     1,     0,     1,     0,     0,     1,     2,     0,     0,     0,    -2,    -2,     0,    -1,     0,     0,     0,    -2,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,     0,     1,    -1,    -3,    -2,     0,     2,     0,     0,     0,     1,     0,     2,     0,     1,     0,     1,    -1,    -1,    -1,    -1,     0,    -1,     1,     0,     0,     0,     0,    -2,     0,     0,     1,    -2,     1,     3,     0,     0,     0,    -1,     1,     0,    -1,    -1,     1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -3,     0,     0,     0,     2,     2,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     1,     0,     0,     1,     2,     2,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,     1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     1,    -1,    -1,    -1,    -2,    -2,     0,     0,     1,     0,    -1,     1,     0,    -2,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,    -2,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -3,    -2,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     1,     2,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -2,     0,     1,     0,     0,    -1,    -2,     1,     1,    -1,     2,     0,    -1,    -2,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     1,     1,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,    -1,    -1,     0,     1,    -2,    -1,    -1,     1,     1,     0,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -3,    -4,    -4,    -2,     0,    -1,    -2,    -3,    -3,    -3,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0),
		    65 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,     1,     0,     1,     2,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     1,     1,     1,     2,     2,     1,    -1,    -1,     1,     2,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,    -2,     1,     1,     0,     0,    -2,    -1,    -1,    -2,    -1,     1,    -1,    -1,     1,     0,    -1,     0,     1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -1,     1,     0,     0,     1,     2,     0,    -3,    -1,    -1,    -1,    -1,     1,     1,     1,    -1,    -1,     1,     1,     0,     0,     0,     1,    -1,    -1,    -2,    -3,    -3,    -2,     0,     1,     0,     2,     2,     0,    -1,    -1,     0,     0,     1,     2,     1,     1,     0,     0,     3,     3,     1,     0,     0,     1,    -1,    -1,    -1,    -3,    -3,    -2,     1,     0,     0,     1,     1,    -1,     1,     1,     1,     2,     2,     2,     0,     1,     0,    -1,     1,     3,     0,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     1,     1,     2,     3,     2,     2,     0,     0,     1,     0,     0,     2,     1,     0,     0,    -2,    -2,    -2,    -2,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,     2,     1,     0,    -1,    -1,     0,     0,    -1,     1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,     1,    -1,     0,     0,    -1,    -2,    -5,    -5,    -4,    -3,    -4,    -4,    -1,    -2,    -4,    -2,     0,     2,     2,     0,     0,     0,     0,     2,     0,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -3,    -4,    -5,    -5,    -5,    -5,    -3,    -2,    -3,    -2,    -1,     0,     2,     0,     0,     0,     1,     1,    -1,    -2,    -1,    -1,     0,     1,     0,     0,     2,     0,     0,    -1,    -2,    -1,    -2,    -2,    -3,    -3,    -3,    -2,    -1,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     1,     1,     1,    -1,    -1,    -1,    -1,     0,    -3,    -4,    -3,    -2,    -1,     0,    -1,     0,    -1,     0,     1,     0,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -2,    -1,     1,     0,     1,    -1,    -1,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     1,     2,    -1,     0,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     0,     1,     1,     0,     1,     0,    -1,     0,     0,    -2,     0,     0,    -1,    -2,    -2,     0,    -1,    -2,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,     0,     1,    -1,     0,     0,     0,    -1,     0,     1,    -1,    -1,    -2,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,    -2,    -3,    -2,    -2,    -1,     1,     0,     0,    -2,    -1,     1,     0,     0,     0,     1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     2,     0,     0,    -1,    -2,    -3,    -3,    -4,    -1,     0,    -1,    -2,     0,     1,     0,     0,     1,    -1,    -1,     1,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,    -2,     0,    -1,    -2,     0,     0,     0,    -1,     0,     0,     1,     1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,     0,     2,     1,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,    -1,    -1,     0,     1,     0,    -1,     1,     1,    -1,     0,    -1,     0,     0,     0,    -2,     2,     1,    -1,     0,    -1,     0,     2,     2,     1,     0,    -1,     1,    -1,     0,     1,     0,     0,     0,     0,     0,     2,     0,    -1,     0,     0,     0,     0,     1,     2,     2,     1,     1,     0,     0,    -1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     2,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     1,     0,    -1,     0,     3,     1,     1,    -1,    -1,     0,     0,     0,     0,     2,    -2,    -2,    -1,    -1,    -2,     0,    -1,    -1,     0,     1,     0,     0,    -3,     0,     1,     0,     1,     2,     3,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     1,     1,    -3,    -3,    -3,    -3,    -1,     1,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0),
		    66 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     1,     0,     1,     1,    -1,    -1,     0,     0,     1,     1,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     1,     1,     1,     1,     1,     1,     0,     1,     1,     1,     2,     2,     1,     3,     2,     1,     1,     0,     0,     0,     0,    -2,     1,     0,     2,     2,     2,     2,     3,     3,     3,     4,     2,     3,     2,     1,     0,     0,     0,    -1,    -1,    -1,     0,     1,    -2,    -2,     0,     0,     0,    -1,     0,     1,     2,     2,     2,     1,     3,     2,     1,     2,     0,     3,     2,     1,     1,     0,     1,     2,     1,     0,    -1,    -1,    -2,    -1,     2,     0,     0,    -1,    -1,     2,     1,     1,     2,     1,     1,     2,     0,    -1,     1,     2,     1,     0,     2,     0,    -1,     0,    -1,     0,     0,     2,     1,     2,     1,     0,     0,     0,     0,     2,     1,     2,     1,     0,     1,     0,    -1,     1,     0,     1,     0,     0,     0,    -2,     0,     0,    -1,    -1,    -1,     0,     1,     2,     2,     0,     0,     0,    -1,     2,     1,     1,     1,     0,    -1,    -1,     0,    -1,    -2,     1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     1,     1,     0,    -1,    -1,    -3,     2,     1,     0,    -1,     0,     1,    -1,    -1,    -1,    -1,     0,    -1,    -3,    -1,    -1,     0,     1,     1,    -1,    -1,    -1,    -3,     0,    -2,     0,     0,    -1,    -2,     2,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,    -1,    -3,     0,     0,     0,     1,     0,     0,    -2,    -3,    -2,    -2,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,    -2,    -1,    -2,    -2,    -2,    -2,     0,     0,     0,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,    -2,    -2,    -1,     0,     0,    -1,    -2,     0,     1,     1,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,    -2,    -1,    -2,    -1,     1,     1,    -1,     1,     1,     0,    -3,    -1,     0,     0,    -1,    -2,    -1,     1,     0,    -1,    -1,     1,     2,     1,     1,     1,     1,     0,     0,    -2,    -1,     1,     1,     1,    -1,     1,     1,    -1,    -3,     0,     0,     0,     0,    -2,    -2,     1,    -1,    -2,     0,     1,     2,     2,     2,     1,     0,    -1,     0,    -1,     0,     1,     0,     1,     1,    -1,     0,     2,    -2,    -1,     0,     0,    -1,    -1,    -3,    -1,    -1,     0,    -1,     0,     0,     1,     0,     2,     1,    -1,    -1,    -2,     0,     1,     0,     0,    -1,     0,     0,     1,    -1,    -3,     0,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,     2,    -1,     0,     0,     0,     0,     1,    -2,    -2,     0,     0,    -2,    -2,    -1,     1,     0,     1,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     1,     1,     1,     1,     1,     0,     0,    -1,     0,     1,    -1,    -3,     0,     0,    -2,    -3,     0,     0,    -1,     0,     0,     0,     1,    -2,     0,     0,     0,    -1,     0,     1,     3,     2,     0,    -1,     0,     0,     0,     2,     0,    -1,     0,     0,    -2,    -2,     0,     1,     1,     0,     0,     0,     2,     2,     1,     0,     0,     1,     0,     1,     0,     2,     0,     0,     0,    -1,    -2,     1,    -1,     0,     0,     0,    -2,    -3,     0,     0,     0,     1,     0,     0,     2,     2,     2,    -1,     0,     0,     0,     1,     1,     1,     1,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     0,    -2,    -2,    -2,    -2,    -1,     1,     2,     0,     1,     0,     3,     1,     0,     0,     2,     1,     1,     1,     0,    -1,     0,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -2,    -3,    -4,    -6,     0,     0,     1,     1,     0,     0,     0,     0,     1,     2,     2,     2,     0,     0,     0,    -2,    -1,    -4,    -1,     0,     0,     0,     0,     0,    -2,    -3,    -3,    -3,     0,    -1,     0,    -1,     0,     1,     0,     1,     1,     0,    -1,     0,     0,     0,     1,    -2,    -3,    -2,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -3,    -4,    -5,    -3,    -4,    -2,    -2,    -1,     0,     1,     1,     2,    -3,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -2,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    67 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -3,     0,     0,     0,     0,    -2,    -4,    -3,    -2,    -2,    -2,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -2,     0,     2,     0,     0,     0,     1,     0,     1,     0,     0,     0,     2,     0,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,    -2,     1,     1,     2,     1,     0,     0,     0,    -1,     1,     0,     0,     1,     0,    -2,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     0,     1,     0,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     2,     2,     0,    -1,    -1,    -2,    -1,    -1,     0,    -1,     0,     2,     0,     1,     1,     0,     2,     1,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,     1,     1,     1,     1,     0,    -2,    -1,     0,    -1,     0,     0,     1,     1,     1,     1,    -2,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     2,     0,     0,     0,    -1,     1,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     1,     0,    -1,     0,     0,    -2,    -1,     0,     2,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,    -1,     1,     0,    -1,    -1,    -2,    -2,    -2,    -1,     1,    -1,    -2,    -1,    -2,    -1,    -1,    -2,    -2,    -3,    -1,    -1,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -4,    -3,    -2,     0,    -1,     0,    -1,    -2,    -2,    -2,    -2,    -3,    -2,     0,    -1,    -1,     0,     1,     0,     1,     0,     1,    -2,    -1,    -2,    -3,    -5,    -4,    -2,    -2,    -1,     0,    -1,     0,     1,     0,    -1,     0,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,    -3,    -2,    -2,    -2,     0,     0,     0,    -1,     0,     0,     1,     1,     0,     1,     1,     0,     0,     0,     1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -2,    -1,     2,    -1,    -1,     2,     1,     0,     0,     1,     1,     0,     1,    -1,     0,    -1,    -1,     0,     0,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     1,     1,     0,    -2,    -2,    -2,    -2,    -1,    -3,    -2,    -2,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,     1,     0,     2,     0,     2,    -1,     1,     1,     0,    -2,    -2,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,    -2,    -1,    -1,     1,    -1,    -1,    -1,    -1,    -1,     2,     2,    -1,    -1,    -1,     1,     1,     1,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,    -2,    -1,     0,     0,     1,     0,    -3,    -1,     0,     1,     1,    -1,    -2,    -1,     0,     1,     0,    -1,    -3,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,     0,    -1,    -1,    -2,     0,     0,     1,     0,     1,    -2,    -1,    -1,    -1,     0,    -1,    -3,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -2,    -1,     1,     0,     1,     0,     1,    -1,    -1,    -1,    -3,    -4,    -3,    -2,    -1,    -2,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -3,    -3,    -4,    -2,    -2,    -1,    -1,    -1,     0,     0,    -2,    -3,    -2,    -2,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -3,    -4,    -4,    -3,    -2,     0,     0,     0,     1,     0,     0,    -2,    -2,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -3,    -2,     1,    -1,    -1,     0,     2,     0,     0,     0,     1,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     1,     1,    -1,    -1,     1,     1,     1,     0,     0,     0,     4,     3,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     1,     2,     1,     1,     1,     0,     1,     1,     2,     3,     2,     1,     0,    -1,     0,     0,     0,     0,     0),
		    68 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,    -1,     0,    -2,    -1,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     2,     2,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     1,     2,     2,     1,    -1,    -2,    -1,     1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     1,     1,     1,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     1,     0,     1,     1,     1,    -1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,    -1,     1,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -2,    -1,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,    -1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     1,     0,     0,    -1,    -1,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,     0,     1,     1,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     1,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    69 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,    -4,    -2,    -2,    -1,    -2,    -1,    -3,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -2,    -4,    -5,    -7,    -6,    -4,    -5,    -5,    -5,    -7,    -6,    -2,    -3,    -4,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -4,    -3,    -3,    -3,    -2,    -1,     0,     0,    -1,    -1,    -1,    -2,    -4,    -7,    -4,    -4,    -4,    -2,    -2,    -3,    -2,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -2,     0,     0,     0,     1,     2,     1,     1,     2,     2,     0,    -1,    -2,    -1,    -4,    -2,    -3,    -3,    -2,     0,     0,     0,    -1,    -3,    -2,    -2,    -1,    -1,     0,     1,     1,    -1,    -1,     2,     1,     2,     3,     2,     0,     1,     0,     0,    -1,     0,     0,    -1,    -2,    -2,     0,    -1,    -2,    -2,    -1,    -3,     0,     0,     0,     1,     0,     0,     1,     2,     2,     2,     4,     2,     0,     1,     1,     0,     1,     1,     0,     0,    -2,    -2,    -2,    -2,    -2,    -2,    -2,     0,     1,     0,     0,     1,     0,     0,     1,     1,     2,     3,     2,     2,     2,     2,     0,     1,     0,     1,     1,     0,    -2,    -1,     0,    -1,    -2,    -2,     1,     1,     1,     1,     1,     1,     0,     0,     1,     2,     2,     1,     1,     1,     0,     0,     1,     0,     0,    -1,    -1,    -2,    -3,    -2,     0,    -1,    -3,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,     1,    -3,    -1,     0,    -5,     0,    -1,     0,     2,     1,    -1,    -1,     0,     0,    -1,     0,    -2,    -1,    -2,     0,     0,    -1,    -1,     1,    -1,    -2,    -1,    -2,     0,    -2,    -1,     0,     0,     0,    -1,     1,     1,     0,    -1,    -2,    -2,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,    -2,    -3,    -2,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     1,    -1,    -1,     1,     0,     0,     1,     1,     0,    -1,    -1,    -3,    -1,    -3,    -2,     0,     0,     0,    -2,    -1,     0,     0,     1,     0,     1,     1,    -1,    -1,    -1,     0,     1,     1,     1,     1,     1,     2,     2,     1,     0,    -2,    -1,    -3,    -1,    -2,     0,     0,    -1,    -1,     0,     1,     1,     0,     1,     0,     0,    -2,    -2,     0,     1,     1,     0,     1,     0,     1,     1,     0,     0,    -1,    -1,    -4,    -2,    -2,     0,     0,    -2,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,     0,    -1,     0,     0,    -1,    -3,    -3,    -1,    -4,    -2,    -1,     1,     0,    -2,     2,    -1,    -1,     0,     0,    -2,    -1,    -1,    -1,    -2,     0,    -1,    -1,     1,     0,    -2,     0,     0,    -1,    -1,    -1,    -1,    -3,    -2,    -1,     0,    -1,    -2,     1,     0,    -1,    -2,    -1,    -2,    -1,     0,    -1,     0,    -1,     0,    -1,     1,    -1,     0,     0,     0,    -1,     0,     1,    -1,    -2,    -2,    -1,     0,    -1,    -4,     0,    -1,     0,     0,    -3,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -2,     0,     2,     2,     1,    -1,     0,     0,     0,    -3,     0,    -1,     1,     1,    -1,    -1,    -2,     0,     0,    -1,    -1,     0,    -1,     1,     1,     0,    -1,    -2,     0,     0,     2,     1,     0,    -3,     0,     0,     0,    -3,     1,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,     1,    -1,     1,     0,     2,     1,     0,    -1,    -1,     0,     2,     2,     2,    -2,    -2,     0,     0,     0,     0,     1,    -1,     0,     0,     2,     1,     0,    -1,     0,     0,     1,     2,     1,     1,     1,     1,     0,    -1,     0,     1,     2,     2,    -1,    -2,     0,     0,     0,    -1,    -2,    -1,     1,     2,     3,     2,     1,     0,     1,     0,     1,    -1,    -1,    -1,     1,     3,     1,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,     0,     1,     2,     2,     2,     2,     0,     1,     0,    -1,     1,     0,     0,     2,     1,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     1,     2,    -1,     1,     0,    -1,     1,    -1,     2,     2,     1,     0,     1,     0,     2,     1,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     1,     1,     1,     0,     1,    -1,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0),
		    70 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,    -1,     0,     0,     1,     2,     2,     1,     1,    -2,    -2,    -1,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     2,     1,     1,     1,     0,    -2,    -1,     1,    -1,    -2,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     1,     1,     0,     0,     2,     0,     0,     0,     0,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     0,     1,     0,     1,     0,     0,     1,     1,     2,     1,     0,     1,     1,     1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,    -1,     1,     0,     1,    -1,     0,     1,     1,     0,    -1,     1,     1,     0,    -1,    -1,     1,     0,     0,     1,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     2,     0,     0,    -1,    -1,    -1,     1,     1,     1,     0,     0,     1,     0,     0,    -1,     0,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,    -1,     0,    -1,    -1,     1,     1,     0,     0,     0,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,     0,    -1,    -1,     0,     0,     2,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     1,    -1,    -2,    -4,    -3,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -3,    -3,    -4,    -2,     1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -2,    -3,    -2,    -1,     0,     1,     0,    -1,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,    -1,     1,     2,     0,    -2,    -2,    -1,    -1,    -2,     0,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -2,    -1,     0,     1,     2,     0,    -1,    -2,    -1,    -1,    -3,     0,     0,     0,     1,     1,     1,    -1,    -1,     1,    -1,    -1,     0,     0,     0,     1,     1,    -1,    -1,    -1,     0,     1,     1,     1,    -1,    -1,    -1,    -1,    -4,     0,    -1,     0,     1,     0,     1,    -1,    -2,    -1,    -3,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,     1,     0,     0,    -2,    -3,    -5,    -2,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     1,     1,     0,    -1,    -2,    -4,    -4,    -3,    -1,     1,     0,     1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     2,     1,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,     1,     1,    -2,    -1,    -1,     0,     1,     1,    -1,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,    -2,     1,     0,     0,     0,     0,     0,     0,     0,    -2,     0,    -1,    -1,     0,     1,     1,     1,     1,     1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     1,     0,     1,     1,     0,     0,    -1,     0,     1,     1,     0,     0,     1,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     1,     0,    -1,     0,     1,     1,     1,     2,     2,     1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -2,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,     0,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0),
		    71 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,     2,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,     0,     0,    -2,    -1,     1,     1,     1,     1,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     1,     0,     0,     1,     0,     0,     0,     0,     1,    -1,    -2,     0,     0,     1,     1,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,     1,     0,     1,     1,     0,    -1,     0,     1,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -3,    -4,    -2,     0,     0,    -1,    -1,     0,     0,    -2,     1,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     1,     1,    -1,    -3,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,     1,     0,     1,     2,     1,     0,    -1,     0,    -1,     0,     0,     0,    -2,    -1,    -2,     0,     2,     0,    -2,    -1,     0,     0,     1,     1,     0,     0,    -1,    -1,    -1,    -2,     0,     1,     1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     1,     0,    -1,    -1,    -1,     1,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,     1,     0,     2,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -1,    -2,     0,     0,     1,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,     1,     1,    -1,     1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     1,     1,    -1,     1,     1,     2,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     1,     0,     0,     0,     1,    -2,    -2,    -1,    -1,    -1,     0,     0,     2,     2,     2,     0,     0,     0,     0,     0,     1,     0,     0,     1,     1,    -1,     0,     0,    -2,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,    -2,    -1,     2,     2,     0,     0,     0,     0,     0,     0,     1,     1,     0,     2,     2,     1,    -1,    -2,    -2,     0,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     1,     2,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,    -1,    -1,    -2,    -1,    -1,    -2,     0,     0,    -1,     0,     0,     0,    -1,     0,     1,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,    -2,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -1,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,     1,    -1,    -2,     0,    -1,    -2,    -3,     0,     1,     0,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     0,    -1,    -1,    -2,     1,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -4,    -3,    -3,    -1,     0,     1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -3,    -1,    -2,    -1,    -2,    -2,    -3,    -2,    -1,     1,     1,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,     1,     1,     0,     0,    -2,     2,     1,     1,     1,     2,     0,     1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     1,     1,     1,     1,     1,     0,    -1,     0,     0,    -1,    -1,     1,     1,     2,     0,     2,     1,     1,     0,    -2,    -1,    -1,     0,    -1,     0,     1,     0,    -2,    -1,     2,     3,     2,     1,     0,    -1,    -1,    -1,     0,    -1,     0,     3,     1,    -1,     0,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,    -2,    -1,    -2,    -2,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,    -1,    -2,    -2,     0,     0,     1,    -1,    -3,    -1,    -1,    -2,    -1,    -2,     2,     2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,    -3,    -1,    -2,    -2,    -3,    -2,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -2,    -2,     1,     0,     1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    72 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -2,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,     1,     1,     0,     0,    -3,    -2,    -3,    -2,    -1,     0,    -1,    -3,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     1,     1,     0,    -1,    -3,    -2,    -3,    -3,    -2,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     1,     1,     0,     0,     1,     0,    -1,    -3,    -2,    -2,    -2,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     1,    -1,     1,     1,     1,     0,     1,    -1,     1,     0,    -1,     0,    -3,    -3,    -2,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     2,     1,     0,     1,     1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,     2,     0,     0,    -2,     0,     0,     0,     0,    -1,     1,    -1,    -1,     1,     1,     0,    -1,     0,    -1,    -1,    -3,    -3,    -2,    -2,    -2,    -1,    -1,    -1,     0,    -1,    -1,     1,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     3,     1,     0,    -1,    -2,    -1,    -2,    -2,    -3,    -1,     2,    -2,    -1,    -1,     0,    -1,    -1,     0,    -2,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     2,     1,    -1,    -1,    -1,    -1,    -2,    -2,     0,     1,    -1,    -1,    -1,     0,     0,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     2,    -1,    -2,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,    -1,    -2,     0,     0,     0,    -2,     0,     0,     1,    -1,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     1,     0,     0,    -2,    -1,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,    -2,     0,     0,     0,    -2,    -3,    -1,    -1,    -2,    -1,    -1,     0,    -1,     1,     0,     0,    -1,    -1,     0,     1,     2,     0,    -1,     0,     1,     1,     0,     0,     0,    -1,    -1,     0,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     1,     2,     1,     0,     0,     0,     3,     1,     0,     0,     1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     2,     1,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     1,     2,     0,     0,     1,     0,     1,    -1,     0,     0,    -2,     0,     0,     1,     0,     1,     1,     1,     1,     1,     0,     1,     0,     1,     1,     1,     0,     1,     0,     1,     0,     0,     2,     0,     1,    -1,     1,     0,    -1,     0,     1,     1,     0,     0,     1,     1,     1,     1,     1,     2,     1,     1,     0,     0,     0,    -1,    -2,     1,     0,     0,     1,     1,     1,     1,     2,     0,    -1,     0,     1,     1,    -1,     0,     0,     1,     0,     0,     1,     1,     0,     1,     1,     1,     2,     1,    -1,     1,     0,    -1,     0,     2,     0,     1,     1,     0,     0,     1,     0,     0,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -1,     0,     1,     2,     1,     1,     1,     2,     0,    -1,     0,     1,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -2,     0,    -1,     0,     0,    -2,     1,     0,     0,     0,     0,     1,     1,     0,     2,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -1,    -3,    -4,    -1,    -1,    -1,    -2,    -2,    -3,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -3,    -4,    -4,    -1,    -1,    -2,    -2,    -3,    -2,    -2,    -2,    -3,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -2,    -2,    -4,    -3,    -4,    -3,    -4,    -4,    -3,    -3,    -3,    -3,    -2,    -3,    -3,    -1,    -3,     0,     0,     0,    -1,     0,    -3,    -1,    -2,    -1,     0,    -1,     0,    -1,    -6,    -4,    -4,    -3,    -3,    -4,    -3,    -3,    -3,    -3,    -2,    -2,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,    -3,    -3,    -2,    -3,    -3,    -2,    -3,    -3,    -2,    -2,    -3,    -3,    -2,    -1,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -3,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0),
		    73 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -3,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -1,     1,     1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,    -3,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     1,     2,     0,     0,     1,     0,     0,     1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -3,    -2,    -1,     0,     0,     0,    -1,     0,     2,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -4,    -1,    -3,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     1,     1,     1,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,    -3,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,     2,     1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,    -3,    -2,    -2,    -1,     0,    -1,     0,     1,     1,     1,     0,     0,     1,     0,    -1,    -2,    -6,    -2,    -1,    -1,    -1,     0,    -1,     0,     1,     2,     0,     1,    -2,    -2,    -1,     0,     0,    -1,     2,     0,     2,     1,     0,    -2,    -2,    -3,    -3,    -4,    -3,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     1,    -2,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -4,    -4,    -3,    -2,    -1,     0,     2,     1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     1,    -1,    -1,    -3,    -3,    -4,     0,     1,     1,    -1,     0,     1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -3,    -5,     2,     2,     0,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -1,    -1,    -1,     1,     0,     0,     0,     1,    -1,    -1,    -1,     0,    -1,     1,     1,     1,     1,     1,     1,     1,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,    -2,    -2,    -1,    -1,     0,     1,     2,     1,     2,     2,     0,    -2,    -1,     0,     0,     0,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -3,    -3,    -1,    -1,     0,     1,     1,     2,     0,     0,    -1,    -1,    -1,     1,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -3,    -2,    -3,    -2,    -3,    -1,    -2,    -1,    -1,    -1,     1,     1,     1,     0,    -1,     0,    -1,    -2,    -2,     0,    -1,     0,     0,    -1,     0,     2,    -1,     0,    -2,    -4,    -4,    -6,    -8,    -6,    -5,    -2,     0,    -1,     0,     1,     1,     1,     0,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,     0,     1,     3,     2,     0,     0,    -2,     0,    -1,    -1,    -2,    -1,    -1,     0,     1,     0,     0,     1,     0,     1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     1,     3,     2,     2,     1,     1,     1,     1,     1,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     2,     2,     2,     1,     0,     0,     1,     0,     1,     2,     0,     1,    -2,     0,     0,    -1,     1,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,     1,     2,     0,     1,     1,     0,     0,     1,     1,     1,     1,     0,     0,    -1,     0,    -3,    -1,     1,     1,     1,     1,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     3,     2,     2,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -1,    -1,    -2,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -2,     0,     0,     0,     0,    -2,     0,     0,    -1,     0,     0,    -2,     0,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0),
		    74 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -1,     1,    -3,    -3,    -2,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -3,    -4,    -3,    -1,     0,    -1,    -2,    -1,    -2,    -3,    -3,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -4,    -1,    -2,     0,    -3,    -3,    -2,    -3,    -4,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -2,    -3,    -1,     0,     0,     0,     0,     0,    -3,     0,     0,     0,     1,     0,    -2,    -1,    -1,     0,     1,     1,     1,     0,     1,     1,     0,    -1,     0,     3,     0,     0,    -1,    -2,    -1,     0,     0,    -1,    -2,     0,     1,     0,     2,     1,     1,     1,     0,     1,     1,     2,     0,     0,     1,     1,     2,     0,     1,     1,     2,     2,     1,    -2,     0,     0,     0,    -1,     0,     1,     1,     0,     2,     2,     2,     1,     1,     0,     2,     2,     3,     2,     0,    -1,     0,     1,     0,     0,     2,     2,     1,     1,    -1,     0,    -1,    -1,     1,     1,     1,     1,     2,     1,     5,     3,     4,     2,     3,     2,     2,     1,     1,     0,     2,     1,    -1,     0,     0,     1,    -1,     3,    -2,    -1,    -2,     2,     1,     1,     0,     2,     1,     0,     4,     2,     3,     0,    -1,     0,     1,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,     0,     1,     1,    -2,     0,    -1,     1,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,    -2,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,     0,    -2,     0,     0,    -1,    -1,    -1,     0,    -1,     1,    -1,    -1,    -1,    -3,    -1,    -1,     0,    -1,    -2,     0,    -2,    -1,    -1,    -1,     0,    -2,     0,    -2,    -1,     0,    -1,    -3,    -1,     0,    -2,     0,    -1,     1,    -1,    -1,    -1,     1,    -2,     0,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     1,    -1,    -1,    -3,    -1,    -1,    -2,    -3,    -1,    -1,    -3,     0,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     0,    -1,     1,     2,     1,    -2,     0,     0,     1,     0,    -1,     0,     1,     0,    -1,     0,     2,    -1,    -2,     0,    -1,    -2,    -2,    -2,     0,     0,     2,     1,    -1,     1,     2,     2,     0,     1,     0,     0,     1,     1,     0,     0,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     1,    -3,    -2,     0,     0,     0,     3,     2,     1,     2,     1,     1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,     0,     1,    -2,     0,     0,     0,     1,     0,     2,     0,     1,     1,     2,     1,     0,     0,     1,     1,     0,     0,     1,     2,     0,    -1,     0,     0,     1,     1,    -1,     0,    -1,    -2,     0,     0,    -2,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     1,     0,     1,     2,     1,     1,     0,     1,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     0,    -1,     1,     0,     0,    -2,    -1,     0,    -1,     0,    -1,     1,     0,    -1,     0,     0,     1,     0,     2,     1,    -2,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,    -2,    -1,     1,    -1,     0,    -1,    -1,    -2,    -1,     2,     3,     2,     1,     2,     1,    -1,    -1,    -2,     0,    -1,    -2,     3,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -2,     0,     0,     1,     1,     0,    -2,     0,     1,     1,     1,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,     1,    -1,    -2,    -2,    -2,    -1,     1,     0,     0,     0,     0,     0,     1,     1,     0,     1,     1,     2,     1,     0,     0,    -2,    -2,    -1,     0,    -1,     0,    -1,     1,     1,    -1,    -1,    -1,     0,     0,     0,     1,    -1,    -1,     0,     1,     1,     1,     0,     2,     3,     3,     3,     1,    -1,    -3,    -2,     0,     0,     0,    -1,    -2,    -4,    -2,     0,     1,     2,    -1,     2,     0,     0,     0,    -1,    -1,     1,     1,     0,     3,     3,     3,     2,     2,     0,     0,    -1,     0,     0,     0,     0,    -2,    -3,    -6,     1,     2,     2,     2,     3,     2,     1,     0,     0,    -1,     0,     0,     1,     3,     3,     1,    -1,     1,     0,     2,    -1,     0,     0,     0,     0,    -1,    -3,    -1,     2,     3,     1,     2,     0,     2,    -1,     0,     0,    -2,    -1,    -1,     1,     3,     0,    -1,     0,     0,    -2,     2,    -1,     0,     0,     0,    -1,     0,     3,     4,     1,    -1,    -1,     0,     1,     1,    -1,     1,    -2,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -2,     4,     3,     2,    -1,    -1,    -2,    -4,    -1,    -1,    -1,    -1,    -3,    -3,    -2,    -1,     0,    -2,    -5,    -4,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,    -2,    -4,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0),
		    75 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -2,    -2,    -1,    -1,    -3,     0,     0,     0,     0,     1,     2,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     1,     1,     1,     0,    -1,    -1,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     1,     0,     1,     0,    -2,    -1,     0,     1,     1,     1,     0,     0,    -1,     0,     0,     1,     1,     1,     1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     2,     1,     0,     1,     1,     1,     1,    -1,    -1,     0,     0,    -1,    -1,     1,     1,     2,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     2,     2,     1,     1,     1,     1,     1,     1,     0,     0,     0,     0,    -1,     0,     2,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     1,     1,     2,     1,     1,     1,     0,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     0,     0,     1,     1,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     2,     1,     1,     1,     0,     0,     0,    -2,    -2,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     1,     1,     2,     2,     1,     0,     1,     0,     0,     0,     0,    -2,     0,     0,     0,     1,    -1,     0,     0,     1,     2,     0,     1,     0,    -1,    -1,     0,     1,     2,     3,     2,     2,     2,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,    -1,     1,     1,     0,     1,    -1,    -1,    -2,     2,     1,     2,     1,     1,     1,     2,     1,     0,    -1,     0,     0,     0,    -2,     1,     1,     1,     1,     2,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     2,     1,     0,     0,     1,     1,     1,     1,    -1,     0,     0,     0,    -2,     0,     1,     1,     1,     1,     1,     2,     1,     1,    -1,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,    -1,    -1,     0,     1,    -1,     0,     0,     0,    -3,     0,     0,     1,     1,     1,     1,     2,     0,     0,     0,     0,    -1,     0,     0,     2,     1,     1,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     1,     2,     2,     0,     0,     0,     1,     0,     0,     1,     1,     1,     1,     1,     0,     0,     0,    -1,    -1,    -2,     0,     0,    -1,     0,     1,     2,     1,     0,     1,     1,     1,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,     1,     2,     1,     0,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,     1,     2,     1,     1,     2,     1,     0,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     1,     1,     1,     0,     0,    -1,    -2,    -2,     0,     0,    -1,     0,     0,     2,     1,     1,     2,     1,     0,    -1,    -2,     1,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,     1,    -1,    -3,    -1,     0,     0,     1,     0,     0,     1,     1,     2,     1,     0,    -1,    -1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -3,    -1,     0,     0,     1,     1,     1,     0,     1,     1,     2,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     0,     1,     1,    -1,     0,    -2,     0,     0,     0,     0,     0,     0,     1,     1,     2,     1,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     1,     0,     1,     1,     2,     1,     0,     2,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     0,     0,     1,     1,     1,     0,     0,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     1,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,     0,     0,     1,    -2,    -2,     0,     0,    -1,    -1,     1,     1,     1,     0,     0,     0,     1,     1,     1,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,    -1,     0,     1,     0,     0,     1,     1,     1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,     0,     0,     0,     0,     0),
		    76 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     2,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     2,     3,     2,     2,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -1,    -1,    -2,     0,     2,     2,     1,     1,     2,     2,     0,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -3,    -2,    -1,    -1,    -1,     0,     0,     2,     0,     2,     1,     0,     1,     1,     0,     0,    -1,    -1,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     2,     2,     2,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     1,     2,     1,     1,     2,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     1,     2,     0,     0,     0,     0,     1,     0,    -2,    -1,     0,     0,    -2,    -2,    -2,    -2,    -2,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,    -2,    -1,     2,    -1,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,    -2,    -2,    -2,    -2,    -1,     1,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,    -2,    -3,    -2,    -2,     0,     0,     1,    -1,    -1,    -2,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -1,    -3,    -2,    -2,    -1,     0,     1,     0,    -1,    -3,    -3,    -2,    -2,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -2,    -2,     0,    -1,     1,     0,     0,    -1,    -2,    -3,    -2,    -2,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     1,     1,     0,     0,    -1,     1,     1,     0,     0,    -1,     0,     1,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     1,     2,     1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -1,     0,    -1,     1,     0,    -1,     0,    -2,     0,     1,     0,     1,     2,     1,     1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     1,     0,     1,     1,     0,     0,     0,    -1,    -1,     0,     2,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,    -1,     1,     1,     1,     1,     1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     1,     0,     0,     1,     2,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     1,     1,     0,     1,     1,     1,     0,     0,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    77 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,    -2,    -3,    -4,    -3,    -2,    -3,    -3,    -3,    -3,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     2,     1,     1,     2,     2,     0,     1,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,    -3,    -3,    -2,    -2,    -2,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,     2,     2,     0,     0,     1,     2,     2,     2,     0,     2,     1,     1,     1,     1,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     1,     0,     0,     0,     1,     2,     2,     1,     1,     1,     2,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -3,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -3,    -3,    -3,    -1,    -1,     0,     0,    -1,     0,    -2,    -1,    -2,    -1,    -1,    -1,     1,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -3,    -2,    -4,    -2,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,     1,     1,    -1,    -2,    -1,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -3,    -2,    -3,    -2,    -3,    -2,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,    -1,     0,     0,     1,     1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     1,     1,     0,     0,     0,     1,     1,     1,     1,     1,     1,     0,     1,     2,     0,     0,     1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,     0,     1,     0,    -1,     0,     0,     1,     1,     1,     0,     0,    -1,     0,    -1,    -2,    -3,    -2,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -2,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     1,     1,    -2,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     1,     0,    -1,     0,     0,    -2,    -2,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     2,    -2,     0,     0,     0,     0,     1,    -1,     0,    -2,    -2,     0,    -1,     0,    -1,    -1,     0,    -1,    -3,    -1,     0,     0,    -3,    -3,    -2,    -2,    -1,     1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,    -1,    -1,    -1,    -2,    -1,    -3,    -3,    -1,    -1,    -2,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     0,     0,     0,     0,     1,    -2,     0,     1,     0,    -1,    -2,    -2,    -2,     0,     0,    -2,     0,    -1,     0,     0,     0,     0,    -2,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -2,    -2,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,    -1,     0,     1,     1,     0,     1,    -2,    -2,     0,     0,    -2,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     0,    -1,     0,     1,    -2,     0,     1,     1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,     1,     1,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    78 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,     1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -1,     1,     1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     1,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     0,     0,     1,     0,     0,    -1,    -1,     1,     0,     0,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,     1,     0,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -2,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,    -2,    -2,    -1,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -2,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -3,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -3,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,     0,     1,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     1,     0,    -1,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,     2,     1,     0,     0,     2,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,     1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    79 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     1,     1,     1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     2,     0,     0,     0,     1,     2,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,    -2,    -1,    -1,    -1,    -1,     1,     1,     1,     1,     0,     1,    -1,    -2,    -2,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -4,     1,    -2,     1,     1,     1,     1,     1,    -1,    -1,    -2,    -4,    -2,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -2,    -3,     2,    -1,     1,     1,     1,    -1,    -2,     0,    -2,     0,    -1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,    -1,    -1,     0,    -2,    -1,    -4,    -1,     2,     0,     1,     0,    -2,    -2,    -1,     0,     0,     1,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     2,     1,    -1,     0,    -1,     1,     2,     1,     0,     1,     2,     1,    -1,    -2,    -1,    -2,    -1,    -1,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,     1,     2,     2,     1,     1,     2,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     1,     0,     2,     1,     0,    -2,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,     0,    -1,    -1,     0,     1,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -3,    -3,     0,     1,     1,     1,     0,     0,    -1,     1,     1,    -2,    -2,    -2,     0,     1,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -4,    -3,    -2,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,    -3,    -2,     0,     1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -2,    -3,    -5,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -3,    -1,     0,    -1,    -1,     1,     0,     0,     0,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -4,    -2,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -3,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -2,    -2,     1,    -1,    -2,    -2,    -3,    -1,    -1,     0,    -1,    -1,    -2,    -1,     0,    -2,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -2,     0,     1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     1,    -2,     0,     1,     2,     1,     0,     0,     0,    -2,    -1,    -2,     0,     0,     0,    -1,    -1,     0,     1,     1,     1,    -1,     0,     0,     0,    -2,    -1,     0,    -1,    -2,    -1,     1,     1,     0,     1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,     1,     2,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     1,     1,     1,     1,     1,     1,     0,     0,     1,     0,     0,    -1,     1,     0,     1,     0,     0,     0,     0,     0,     0,    -2,     0,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,    -1,    -2,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,    -2,     0,     1,     1,     0,     0,     2,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,     0,     1,     2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    80 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     2,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     2,     1,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,    -2,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     1,     0,     1,     1,     2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -3,    -2,     0,     0,     0,    -1,     1,     1,     1,     1,     1,     2,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -2,    -3,    -2,    -3,     0,     1,     0,     0,    -2,    -1,     0,     0,     0,     2,     1,    -1,    -2,    -3,    -1,     0,     0,     0,     0,    -1,     1,     2,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,     1,     1,     0,    -1,    -2,     1,     1,    -1,     1,    -1,     0,     1,     1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     1,    -1,     0,     0,     1,     0,     0,     1,     1,     1,    -1,    -2,    -2,     0,     0,     0,     1,     0,    -1,     1,    -1,    -1,    -1,    -3,    -1,    -2,    -1,     0,     1,     1,    -1,     0,     0,     0,     1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,    -1,     0,    -1,     0,     1,     0,     0,     1,     0,    -1,    -2,    -1,     2,     1,     1,     1,     1,     0,    -2,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,     1,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -3,    -3,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,     1,     1,     1,     1,    -1,    -4,    -4,    -1,     1,    -1,     0,     1,     2,     0,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     1,     1,     1,     0,    -1,    -5,    -2,     1,     0,    -1,    -1,     0,     4,     1,     1,    -1,     0,     0,     0,     0,    -3,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -4,    -3,    -4,    -2,    -1,    -1,    -1,     0,     0,     2,     1,     0,    -2,     0,     0,     0,    -1,    -3,     0,    -1,     0,     1,     0,     1,    -2,    -1,     1,     0,    -3,    -2,    -1,     0,    -1,    -1,    -2,     0,     0,     1,     2,    -1,    -2,    -1,     0,     0,     0,    -2,     1,     0,     0,     1,     1,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     1,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     1,     1,     1,    -1,     0,     0,    -1,    -3,    -2,    -1,     0,    -1,     0,     0,     1,     1,    -1,    -1,     0,     1,    -2,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,     1,     2,     1,    -1,    -3,    -2,    -1,     0,     0,     0,     0,     1,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,    -2,    -1,     2,     0,     0,     1,     0,     1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     1,     0,     1,    -1,     0,     0,     0,     0,    -2,     1,     2,     0,     1,     0,     1,     1,     0,     0,    -1,    -1,     0,    -2,     0,     0,     0,    -2,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,     1,     0,     0,     1,     1,     0,     1,     0,     0,    -1,    -1,     0,     1,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,     1,    -1,     0,     0,     0,     0,    -3,     0,     0,     1,     1,     1,     1,     0,     1,    -1,    -1,     0,     1,     0,    -2,    -2,    -1,    -1,    -3,    -2,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,     0,     0,     0,     1,     1,     1,     0,     1,     1,    -1,    -2,    -1,    -2,    -2,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     2,     2,     0,    -1,     0,     1,     2,     1,     2,    -2,    -2,    -2,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -2,    -3,    -2,    -1,    -2,    -2,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    81 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     2,     4,     3,     2,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,    -2,    -1,     1,     0,    -1,    -2,    -1,     0,     1,     2,     3,     0,     0,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     1,     1,     0,    -1,     2,     2,     1,     0,     0,    -1,     0,     1,     1,     0,     0,    -1,     1,     1,     1,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     2,     3,     1,     1,     1,     0,     0,    -2,    -2,     0,     1,     0,    -1,     0,     0,     1,     1,     1,     1,     0,     0,     0,    -1,    -1,     0,     0,    -2,     0,     0,     1,     1,     0,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,     1,     0,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,     0,     1,     1,    -2,     0,     1,    -1,     0,    -1,     0,     1,     0,     0,     1,     2,     0,     0,     1,     0,    -1,     0,    -1,    -1,     0,     0,    -3,    -2,    -2,     0,     0,     0,     0,     1,     0,     0,     1,    -1,    -1,     0,     1,     0,     1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,    -3,    -1,    -1,    -1,     0,     1,     1,     0,     0,     2,     2,    -1,    -2,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,     0,    -2,    -1,    -2,     0,     1,     1,     1,     2,     1,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,     0,    -1,     1,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     0,    -2,     1,     1,     1,     2,    -1,    -1,     0,     0,    -1,    -1,     1,     0,    -1,    -1,    -4,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,     1,     1,     0,     0,    -2,    -3,    -2,    -1,    -1,     0,     1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -3,     0,     1,     0,     0,    -1,    -1,    -3,    -2,    -2,    -1,    -2,    -4,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -3,    -2,     0,     2,     1,     0,    -1,    -1,    -2,    -2,    -3,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -4,    -2,    -2,     1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,    -2,    -2,     0,    -1,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -3,    -2,    -2,    -6,    -5,    -3,     0,    -1,     0,     0,     0,     0,     1,     1,     2,    -1,    -4,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -3,    -2,     0,     0,    -1,    -2,    -3,    -2,    -1,    -1,     1,     1,     0,    -1,     0,     1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,     1,     0,    -2,    -1,     0,     0,     1,     2,     0,     0,     0,     1,     1,     2,     1,     2,     2,     2,     0,     1,     1,     0,     0,    -1,     0,     1,     0,    -1,     1,     1,     0,     1,     1,     2,     2,     1,     1,     0,     1,     1,     1,     0,     1,     2,     1,     1,     0,    -1,    -1,     0,     1,    -1,     0,     1,     0,    -3,    -2,     1,     2,     1,     0,     0,     1,     1,     0,     0,     1,     0,     0,    -1,     1,     0,     1,     1,     1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     1,    -1,    -2,    -2,    -2,    -1,     0,     1,     1,    -1,    -1,    -1,    -2,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -2,    -1,    -3,    -2,    -2,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    82 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,     0,     0,     0,     2,     2,     1,     0,     1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,     0,     1,    -1,     1,     0,     0,    -1,     1,     1,     1,     1,     0,    -1,    -1,    -1,     0,    -1,    -3,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,    -2,     1,     2,     0,     0,     1,     1,     0,     1,     0,     2,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,     0,    -2,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,    -1,     1,     0,     0,    -1,     0,     1,     0,     0,    -2,     0,     1,     1,     0,    -2,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,    -1,     0,     1,     1,     1,     1,    -1,    -1,    -2,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -1,     0,    -1,    -2,     0,     0,    -1,     0,     0,     1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,    -4,    -6,    -6,    -4,    -4,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -4,    -5,    -4,    -4,    -2,    -1,    -2,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     1,    -1,    -2,     0,    -1,    -1,     0,    -1,    -2,    -2,    -3,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,     0,     1,     1,    -2,    -2,     2,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     2,     1,     0,    -1,     0,     2,     2,     1,     0,     0,     0,    -1,    -1,     0,     1,     2,     0,     0,     1,     0,     0,     0,    -1,    -1,     2,     1,     0,     2,     2,     2,     1,     2,     1,     1,     2,     2,     0,     1,    -2,    -1,     0,     1,     0,     0,     0,     0,     1,     1,     1,     0,    -1,     0,     4,     2,     2,     1,     1,     1,     1,     2,     1,     1,     1,    -1,     1,     0,     0,    -1,     0,    -1,    -1,     0,     1,     0,     1,     3,     2,     0,     0,     0,     1,    -1,     2,     3,     1,     1,     1,     1,     0,    -1,     1,     1,     1,     0,     1,     0,     0,    -1,    -1,    -1,     0,    -1,     2,     3,     1,     0,     0,     0,    -1,     1,     1,     2,    -1,     1,    -1,    -1,     0,     0,     0,     1,     1,     1,     0,     0,    -1,     0,    -2,    -1,    -2,    -2,     0,     1,     2,     0,     0,    -1,     0,     0,     1,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,     1,     1,     1,    -1,    -1,    -1,     0,     1,     1,     2,     0,    -1,    -1,     0,     1,     1,     1,     1,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     1,     1,     0,     2,     2,     1,     1,     0,    -1,     0,     0,     1,     2,     1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     2,     0,     1,     0,     0,     1,     0,     0,     1,     1,     1,     0,     1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     1,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -2,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     2,     1,     0,    -2,     0,    -1,    -2,    -1,    -1,     0,    -2,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     0,     1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -2,    -2,    -3,    -2,    -2,    -2,    -1,    -1,    -2,    -3,    -2,    -3,    -2,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -2,    -1,     0,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0),
		    83 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,     1,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     4,     3,     1,     1,     1,     1,     0,     0,     2,     2,     1,     1,     3,     5,     1,    -3,    -3,    -2,    -1,     0,     0,     0,     0,    -2,     0,     1,     1,     0,     2,     3,     0,     2,     1,     1,     0,     1,     0,     1,     2,     1,     1,     1,    -2,    -2,    -7,    -5,    -2,    -1,     0,     0,     0,     0,     0,     0,     1,     2,     3,     0,     1,     1,    -1,    -1,     0,    -1,     0,     1,    -1,     0,     1,     0,     0,     0,     0,     1,    -2,    -1,     0,     0,     0,     1,     0,     0,     2,     3,     3,     1,     1,     1,     0,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,    -3,    -1,     0,     0,     0,     0,     1,     0,     0,     3,     4,     2,     0,     0,     2,     0,    -1,     0,     0,     1,    -1,    -1,     1,    -1,    -1,    -1,     0,     1,    -3,    -2,    -1,    -1,     0,    -1,     0,     1,     2,     0,     1,     0,     0,     0,    -1,    -2,    -1,     0,     2,     1,     1,    -1,     1,     0,    -1,     1,     0,    -1,    -2,    -2,     0,     0,    -1,    -3,    -1,     3,     3,     1,     1,     2,    -1,     1,    -1,    -1,     0,    -1,    -1,     0,     2,     1,     0,     1,    -1,     2,     1,    -4,    -2,    -1,     0,     0,     0,    -3,     0,     1,     2,     2,     2,     0,    -1,    -2,    -2,    -1,    -2,     0,    -1,     0,     1,     1,     0,    -1,    -1,     1,     2,    -2,    -2,    -1,     0,     0,    -1,    -2,     2,     3,     3,     2,     1,     1,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -2,    -1,     0,    -1,    -4,    -3,    -1,     0,     0,     0,    -2,     1,     2,     3,     2,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,    -1,    -2,    -1,     0,    -3,    -2,    -1,     0,     0,     0,    -1,     0,     3,     2,     1,     1,     2,     0,     1,    -1,    -1,     0,    -1,     1,    -3,    -1,     1,     1,    -1,    -1,    -1,     1,     0,    -3,    -1,     0,     0,     1,     0,     1,     1,     2,     2,     0,     1,     0,    -1,     0,     0,    -1,     1,    -1,    -1,     0,     1,     1,     1,     0,    -1,     1,     0,    -4,    -2,     0,     0,     1,    -1,     0,     1,     3,     2,    -1,    -1,    -2,     0,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,     2,     0,     0,     1,     2,     2,    -4,     1,    -1,     0,     0,     0,     3,     2,     2,     0,     1,    -2,     0,     0,    -2,    -2,     0,     0,    -1,    -2,    -1,     1,     2,     0,    -1,     1,     0,     1,    -5,    -2,    -1,     0,     0,    -1,     1,     2,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     1,     2,     0,     0,    -1,    -1,    -1,    -4,    -1,    -1,    -1,     0,     0,     1,     2,     1,     0,     0,    -1,    -1,     0,     0,    -1,     1,     0,     1,     0,     1,     2,    -1,     1,    -1,     0,    -2,    -1,    -4,     0,    -1,     0,    -1,     1,     0,     1,     1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     1,     1,     0,     1,     1,    -1,     1,     0,    -1,    -1,     1,    -2,    -1,    -1,     0,     1,    -2,     0,     1,     1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     1,     1,     2,     2,     0,     0,     1,     1,     1,     1,     0,    -3,    -1,     0,     0,     0,     1,     0,     0,    -1,     1,     2,     0,     0,    -1,     0,     1,     1,     2,     2,     1,     1,     1,     2,     0,     1,     1,     0,    -2,    -3,    -1,     0,     0,     0,     1,     1,    -1,     1,     2,     2,     0,     0,     1,     0,    -1,     0,     1,     1,    -1,     1,     0,     1,     0,     1,     3,     1,    -2,    -2,    -1,     0,     0,     0,     1,     0,    -1,     0,     1,     2,     1,     1,     0,     1,     0,    -1,    -1,     1,     1,     0,    -1,    -1,     0,     3,     3,     1,     2,     1,    -1,     0,     0,     0,     2,     3,     2,     0,     2,     2,     1,     2,     1,    -1,    -1,     0,     1,    -1,     0,     0,    -1,     1,     3,     2,     1,     1,    -2,    -1,     0,     0,     0,     0,     0,    -1,     0,     2,     2,     0,     1,     1,    -1,     0,     1,     2,     0,     0,     0,     0,     1,     1,    -1,    -3,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -3,     1,     1,     0,     1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     3,     3,     3,     1,    -1,    -1,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -2,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0),
		    84 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -2,    -3,    -4,     0,     1,     0,    -2,    -2,    -2,    -3,    -2,    -4,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -3,    -2,    -2,    -1,    -2,    -2,    -3,    -3,    -3,    -2,    -4,     0,     0,    -2,    -1,    -1,     0,     1,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -3,     0,     0,     1,     0,    -2,     0,     0,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     1,     1,    -1,    -2,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     1,     0,     1,     0,     1,    -1,    -1,    -2,    -1,     1,     0,     0,    -1,    -1,     0,     0,    -1,     1,    -1,     0,     0,     0,    -1,    -1,     1,     2,     1,    -1,    -1,    -2,     0,     0,     0,    -1,    -2,    -3,    -2,    -1,    -2,    -1,    -3,     0,     0,     0,    -1,     0,     0,    -1,     0,    -3,    -1,     0,     1,     1,    -1,    -2,    -2,    -1,    -1,     0,    -2,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,     1,    -2,    -1,    -3,     2,     0,     1,     1,    -2,    -2,    -3,    -1,    -2,    -1,    -1,     0,    -3,    -2,    -2,     0,    -1,     0,    -1,    -1,    -1,     0,     1,     1,     0,    -1,     0,    -2,     1,     0,    -1,     0,    -2,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -2,    -1,    -1,     0,     0,     1,     1,     1,     1,     1,     2,    -1,    -2,    -1,     0,    -1,     1,     0,    -1,     1,    -1,    -2,    -1,     0,     0,     0,     1,     0,    -1,     1,     1,     2,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,     0,     0,     2,     0,     0,     1,     2,     2,     1,     2,    -1,     0,     1,     2,     0,    -1,     0,     0,     0,     1,     1,     0,     0,    -2,    -2,     0,     0,     1,     1,     0,     1,     1,     1,     1,     2,     1,     1,     2,     1,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,     1,     2,     1,     1,    -2,     0,     0,     0,     2,     1,     2,     1,     1,     0,     1,     1,     2,     2,     1,     0,    -1,     1,     1,    -1,     0,     0,     1,     1,     1,     1,     3,     3,    -1,     0,     0,    -3,     1,     3,     2,     1,     1,     2,     1,     1,     1,     1,     0,     0,    -1,     1,     2,    -1,     2,    -1,     2,     1,    -1,     0,     2,     2,     0,     0,     0,     3,     1,     0,     1,     1,    -1,     0,     1,     1,     1,     0,     0,     0,     1,     2,     0,     0,     1,     0,     0,     2,     1,    -1,     1,     3,     0,     0,     0,    -1,     2,     1,     1,     2,     1,     1,     0,     0,     0,     1,     0,     0,     2,     1,     1,     2,     2,     1,     0,     0,     0,     0,     1,     2,    -1,     0,     0,     1,    -1,     2,     2,     1,     1,     0,     0,     0,     0,     0,     1,     1,     1,     1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     1,     0,    -2,     0,     2,     1,     2,     0,     0,     0,     1,     1,     0,     1,     0,     1,     1,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,     0,    -1,    -1,     2,     0,     2,     0,    -1,     1,     0,    -1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,    -2,     2,     1,     0,     0,     0,     0,    -1,    -3,    -2,    -2,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -3,    -2,    -2,    -2,    -1,    -3,    -1,     0,     0,     0,    -2,     1,     1,     0,    -1,    -2,    -1,    -1,    -2,    -1,    -2,    -1,    -2,    -1,     0,    -1,    -1,    -2,    -1,    -2,    -1,    -1,     0,    -2,    -2,     0,     0,     0,     0,    -2,    -3,     0,     0,    -2,    -2,    -2,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -2,     0,     0,     1,    -1,    -1,     0,    -1,     0,     0,     0,    -2,    -1,    -3,     0,     1,     0,    -2,     1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -2,     0,     1,     1,     1,     1,    -1,     0,    -2,     1,     1,    -1,     0,    -1,    -3,    -2,     0,     1,     0,    -1,    -4,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -2,     0,     0,    -1,    -2,    -1,    -1,    -2,    -2,    -1,    -3,     0,    -1,    -1,    -2,    -1,     0,     1,     0,    -2,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     0,    -2,    -2,    -1,    -1,    -3,    -2,    -2,    -3,    -3,    -2,    -3,    -1,    -1,    -3,    -4,    -4,    -4,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -1,    -2,    -3,    -1,    -1,    -3,    -2,    -2,    -2,    -2,    -2,     0,     0,     0,     0,     0),
		    85 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -3,    -2,    -4,    -3,    -2,    -3,    -3,     0,     0,     0,     1,    -1,     1,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,    -1,     1,     1,    -1,    -3,    -3,     0,     0,     1,    -2,    -2,     0,    -1,     2,     1,     1,     2,     2,     2,     4,     3,     2,    -1,     1,     1,     0,     0,     0,    -1,     1,    -3,    -3,    -2,    -1,    -3,    -1,     1,    -1,    -1,    -2,     0,     2,     1,     2,     5,     2,     2,     3,     5,     2,    -2,     0,    -1,    -1,     0,     0,    -2,     2,    -4,    -1,    -1,    -1,     0,     1,     1,     0,    -1,    -2,     1,     1,     2,     2,     3,     3,     4,     1,     2,     1,    -1,    -1,    -2,    -2,     0,     0,     0,    -3,    -1,     2,     2,     1,     2,     1,     1,     0,     0,    -2,     0,     0,     0,     0,     2,     3,     2,     0,     2,     1,     2,     2,     0,     0,     0,    -1,     0,    -4,    -2,    -1,     1,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -2,    -1,    -1,     1,     2,     1,     1,     4,     3,     3,     1,     1,     2,    -1,    -1,    -2,    -4,    -1,    -1,     1,     1,     0,     0,    -1,     1,     1,     0,    -1,    -2,    -2,     0,    -1,     2,     2,     2,     3,     3,     2,     0,     1,     1,     0,     0,    -2,    -2,    -1,    -1,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     0,     2,     0,     1,     2,     2,     2,     1,     0,     0,     0,     0,    -1,    -4,     1,     0,    -1,    -2,     0,     1,    -1,     1,     1,    -1,    -1,    -1,    -3,    -2,     1,     0,     0,     2,     2,     2,     3,     1,    -1,    -1,     0,     0,     0,    -3,     1,    -1,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     1,     1,     0,     0,    -1,     0,     1,     2,     3,     2,    -1,    -1,     0,     0,     0,    -2,     2,     0,     0,     1,     1,     1,     2,     0,     2,    -1,     0,    -2,     0,    -1,     0,    -1,    -2,    -1,     0,     1,     1,     2,     3,    -1,     0,     0,     0,    -2,     0,     0,     0,     2,     0,     0,     1,     1,     1,     0,    -1,     0,     0,    -1,    -2,     0,    -1,     1,    -1,    -2,    -2,    -1,     2,    -1,     0,     0,    -1,    -2,     1,     1,     2,     0,     0,     1,     1,     1,    -1,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     1,     0,     0,    -2,    -2,    -1,     1,     0,    -1,     0,     2,     2,     0,     1,     0,     1,     1,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,    -1,    -2,    -1,     0,     0,    -2,    -1,     1,     2,     3,     1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -2,     0,     1,     0,    -1,     1,     1,     0,    -2,    -3,    -3,    -1,     0,     0,    -2,     0,     1,     3,     1,     3,     2,     0,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     1,     0,    -1,    -3,    -5,    -3,    -1,     0,    -2,     0,     0,     1,     3,     2,     2,     1,    -1,    -1,    -2,    -2,     1,     0,     0,    -2,    -1,    -1,     1,     0,     0,     0,    -1,    -3,    -3,    -2,     0,    -1,     1,     2,     0,     2,     3,     1,     0,     0,     0,     0,    -1,    -2,     0,     1,     1,     0,    -1,     0,    -1,     1,     0,     1,     1,    -1,    -3,    -2,     0,    -1,     2,     1,     2,     3,     1,     0,     1,     1,     0,     1,    -1,     1,     0,     2,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,     1,    -4,     0,     0,     0,    -2,     0,     1,     2,     3,     1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     1,     1,     0,    -1,     1,     0,     0,     0,     0,    -3,    -2,     0,     0,     0,     1,     0,     0,     0,     1,    -1,    -1,     1,     1,     1,     1,     0,     1,     1,     0,    -1,     0,     0,     1,     2,     0,     0,     0,     1,     0,     0,     0,     1,     1,    -1,     0,     2,     1,     1,     2,     1,     1,     1,     0,    -3,    -1,     0,    -1,    -1,     0,     1,     1,     3,     0,     0,     0,    -2,    -1,    -2,     0,     0,     0,     1,     1,     0,     1,     1,     2,     1,     1,     2,     1,     1,     0,    -1,     0,    -1,    -2,     0,    -3,    -1,     0,     0,     0,     0,     1,    -3,    -3,     0,    -1,     0,    -1,     0,     0,     0,     1,    -1,     2,     2,     2,     1,     2,     2,     2,     3,     3,     2,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -4,    -2,    -1,     0,     1,     2,     4,     2,     3,     1,     0,    -1,     1,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -3,    -2,     0,     0,    -1,    -1,    -2,    -3,    -2,    -1,     0,     0,     0,     0),
		    86 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,     0,     1,     1,    -2,     0,     0,     1,     1,     1,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     1,     1,     1,     2,     1,     1,     1,     1,     1,     0,     1,     1,     1,     2,     3,     2,     2,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     1,     2,     2,     2,     2,     3,     2,     1,     2,     1,     0,     0,     2,     2,     0,     1,     2,     2,     2,     2,    -1,     0,     0,     0,     0,    -2,    -1,     1,     2,     3,     2,     1,     2,     2,     1,     2,     0,     1,    -1,     1,     1,     0,     1,     2,    -1,     0,     1,     1,     1,     0,     1,     0,     0,    -1,    -1,     1,     1,     1,     1,     2,     2,     2,     1,     1,     0,     0,     0,     1,     1,    -1,    -1,     0,    -1,     1,     1,     1,     2,     1,     0,     0,     0,     0,     0,     1,     0,     2,     1,     0,     2,     2,     1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,     2,     0,     1,     1,     1,     0,    -1,     0,     0,     0,    -1,     1,     1,     0,     2,     1,     2,     1,     0,     0,    -1,     0,    -1,     0,     1,     2,     0,     1,     1,     0,    -1,     1,     0,    -1,    -1,     0,     0,    -1,    -1,     1,     0,     0,     1,     1,     1,     1,     0,     0,    -1,     0,    -1,    -1,     2,    -1,     1,     1,     2,    -2,    -2,    -2,    -3,    -2,    -2,     0,     0,    -1,    -2,     1,     0,    -1,     0,     1,     0,     0,     1,     0,     0,     0,    -1,    -1,    -2,    -1,     1,     1,    -1,    -2,    -2,    -1,    -2,    -1,    -2,     0,     0,    -1,    -2,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     1,     0,     0,    -2,    -2,    -2,    -1,     1,     0,    -1,    -2,    -2,    -2,    -1,    -1,    -3,     0,     0,    -1,    -2,     0,     0,     0,    -1,    -2,    -1,     0,     1,     1,     0,    -1,    -1,    -1,    -1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,    -2,     0,     0,    -1,    -1,    -3,     0,     0,     0,     0,     0,    -1,     0,     1,     2,     2,     1,    -1,     0,    -1,     2,     1,    -1,    -2,    -1,     0,     0,     0,    -2,     0,    -1,    -1,    -3,    -4,    -1,     0,     0,    -1,     0,    -1,     0,     1,    -1,     0,     1,    -1,     1,     0,     2,    -1,    -1,    -2,     0,     0,     0,     0,    -2,    -2,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     1,     2,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,    -3,    -3,    -1,     0,     0,    -1,    -1,     1,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,    -2,    -2,     0,     0,    -1,    -3,     0,     1,    -1,     0,    -2,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -2,    -2,     0,     0,    -1,    -2,     0,    -1,     0,     0,     0,     0,     1,     1,    -1,    -2,    -1,    -1,     0,     0,     1,     0,     0,    -1,     0,     1,     1,     1,    -1,    -3,     0,     0,     0,    -3,     0,    -1,     0,     0,     0,     1,     2,     2,     1,     0,     0,     0,     0,     1,     1,     0,     1,     1,     0,     1,     1,     2,    -1,    -1,     0,    -1,    -3,    -2,     0,    -1,     1,     1,     1,     0,     3,     3,     2,     0,     1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,     2,     2,     2,     3,     3,     3,     1,     2,     2,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -2,     0,    -2,     0,     0,     0,    -2,    -1,    -1,    -2,    -1,     2,     5,     3,     2,     1,     2,     1,     2,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,    -3,    -2,    -2,     0,     0,     0,     0,    -1,    -2,    -3,    -2,     0,     1,     2,     2,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,    -1,    -4,    -2,    -1,     0,     0,     0,     0,    -2,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     1,     1,    -2,    -1,     2,     1,     0,    -2,    -3,    -3,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -2,    -3,    -3,    -3,    -4,    -2,    -3,    -2,     0,     2,     2,     1,    -1,    -1,    -3,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    87 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -3,    -3,    -3,    -5,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,    -2,    -2,     2,     0,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -3,    -1,     2,     0,     1,     1,     1,    -1,    -3,    -3,     0,    -1,    -2,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -3,    -1,    -2,     0,     0,     0,     0,     1,     2,     1,     2,     2,     2,     1,     1,     3,     0,     0,    -2,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     1,    -2,     0,    -2,    -1,    -1,     0,     0,     2,     0,     3,     3,     3,     4,     1,     3,     3,     1,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     3,     1,     0,    -2,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     2,     0,     2,     2,     1,     2,     0,     1,     1,     0,     0,     0,     0,     0,     0,     2,     0,    -1,    -3,    -2,    -1,     0,     0,     2,     1,     1,     0,     0,     1,     1,     0,     0,     0,     2,     1,     2,     1,     0,     0,     0,     0,     1,     0,     1,     1,    -3,     0,     2,     4,     0,    -1,     1,     0,    -1,    -1,    -1,    -1,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,    -1,     1,    -1,    -1,    -1,    -1,     1,     2,     3,     0,    -1,     1,    -1,    -1,    -2,    -1,    -1,    -1,     0,    -2,     0,    -2,    -3,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,    -2,    -2,    -2,     0,     0,     1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -4,    -2,    -2,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -4,    -1,    -2,     0,     0,     0,     1,    -2,    -3,    -1,    -1,    -2,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     1,     0,     1,     1,     0,    -2,     1,    -1,     0,    -2,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     1,     0,     1,     0,     1,     1,    -1,     2,     1,     1,     0,     1,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     1,     1,     0,    -2,     2,     0,     1,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     1,     0,     1,     1,     0,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,     0,    -3,    -2,     0,     0,     0,    -2,    -2,    -2,    -1,     1,     1,     0,     1,     1,     0,     1,     0,     0,     0,     1,     0,    -1,    -1,     1,     0,     0,     0,     0,    -1,     1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,     0,    -1,    -1,     1,    -1,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -3,    -1,    -2,    -3,    -1,     0,     2,     0,    -2,    -1,     0,     1,     0,    -1,    -3,    -3,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -2,    -2,    -2,    -3,     0,     0,    -2,    -2,     0,     0,     0,    -1,    -2,    -1,    -1,    -2,    -3,    -2,    -2,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -2,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,    -3,     0,    -1,    -1,     0,    -2,    -2,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -5,    -4,    -2,    -1,     0,    -2,     0,     0,     0,    -1,    -3,     0,     0,     0,     1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,    -1,    -2,    -3,    -1,    -1,    -1,    -2,     0,     0,     0,     1,     0,     1,     1,     0,    -1,     0,    -1,    -2,     0,     0,     0,     0,    -1,    -1,     1,    -1,    -1,     1,     1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     1,    -1,    -1,    -1,     2,     1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,     0,    -1,     0,     0,     0,     0,    -1,    -4,    -3,    -3,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,     2,     0,    -1,     0,    -2,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     2,     2,     1,     0,    -1,    -1,     1,     2,     2,     2,     0,     0,     0,    -1,     0,     0,     0,     0,     0),
		    88 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -3,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -2,    -2,     1,     1,     0,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -2,    -3,    -2,    -1,     1,     1,     1,     0,     0,    -2,    -2,    -3,    -1,     0,     0,     1,     0,     1,     1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -3,    -2,    -2,     1,     1,     2,     2,     0,    -2,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     1,     1,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -2,     0,    -1,     1,     2,     1,     0,     1,     0,     1,     1,     2,     1,     0,     0,    -1,    -2,    -2,     1,     0,    -1,    -1,     0,     0,    -2,    -2,     1,    -2,    -2,    -1,     0,     0,     1,     0,    -1,     0,     1,     1,     1,     0,     1,    -1,    -1,     0,     1,     1,     0,     1,     0,     0,     0,    -2,    -1,     0,     1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     2,     2,     1,     0,    -1,     1,     1,     1,     2,     1,     0,     0,    -1,    -1,    -1,    -1,     3,     1,     0,     1,     1,    -1,     0,     1,     0,     0,     0,     0,     1,     1,     1,     1,     0,     0,    -1,     0,     1,    -1,     1,     1,     0,     0,    -1,    -1,     1,     3,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     2,     3,    -2,     0,    -1,    -2,    -1,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,     1,     0,    -2,    -2,    -1,    -1,     0,    -1,     1,     1,     1,     1,     2,    -2,     0,     0,    -1,    -1,     1,     0,     1,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,    -3,    -3,    -2,    -1,     0,    -1,     0,    -1,     1,     0,    -1,     1,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -1,    -1,     0,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     0,    -1,    -3,    -4,    -2,     0,     0,     0,    -1,    -2,    -1,    -2,    -1,    -1,     2,     2,     1,     2,     1,     0,     1,     0,    -1,     0,    -1,     1,     2,     1,     0,    -2,    -3,    -3,     0,    -1,     0,     0,    -1,    -2,     0,     1,    -1,     1,     2,     2,     3,     2,     1,     0,     1,     0,    -1,     0,     1,     1,     1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,     0,    -2,     0,     2,     2,     2,     3,     3,     2,     1,     2,     1,     0,     0,     0,     1,     1,     1,     1,     1,    -2,    -1,     2,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,     2,     2,     2,     1,     0,     0,     0,     1,     2,     2,     0,     1,     1,     0,     0,     0,     1,    -3,    -1,     0,     0,    -1,    -1,     0,    -2,    -2,     0,     0,     0,     1,     0,    -1,    -1,     0,     1,     0,     0,     1,     1,     0,     0,     0,     0,     1,    -1,     0,    -1,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,     1,     0,    -2,     0,    -1,     0,     0,    -1,    -3,    -1,    -2,    -2,    -2,    -2,    -2,    -1,    -1,     0,     1,     1,     0,     1,    -1,    -1,    -1,    -1,     0,     1,     0,    -1,    -2,    -1,    -1,     0,     0,    -1,    -3,    -1,    -1,    -1,     0,     0,    -2,    -1,    -1,     1,     1,     2,     1,     1,     0,    -1,     0,     1,     0,     0,     0,    -2,    -2,    -2,     0,    -1,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,    -1,     1,     3,     1,     1,     2,     1,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,     0,    -1,    -1,    -1,     0,     1,     1,     0,    -1,    -1,     0,     0,     2,     1,     1,     3,     2,     1,     0,     0,    -1,     1,    -1,     1,     1,    -1,    -2,    -2,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     1,     2,     0,     1,     3,     2,     1,     1,    -1,     0,     0,     1,     0,     1,     1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     1,     2,     3,     2,     0,     0,    -1,     0,     2,     2,     0,    -2,    -1,    -3,    -1,    -1,     0,     0,     0,    -1,     0,    -3,    -2,     0,    -1,    -2,    -2,     0,     1,     1,     2,     1,     0,    -2,    -1,     0,     0,    -1,    -3,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     2,     1,    -1,    -1,     0,     1,     0,    -3,    -1,    -1,    -2,    -2,    -3,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,     0,     0,    -1,    -3,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0),
		    89 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,     0,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -2,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -3,    -1,    -1,    -1,    -1,     1,     2,     1,     1,     1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,    -3,     0,    -1,     1,     1,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,    -2,    -1,    -3,    -1,    -1,     1,     0,    -1,     0,     0,    -3,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -2,     0,     1,     0,     1,     0,    -1,     0,    -1,    -1,     0,     1,     1,     0,    -1,    -1,    -1,    -1,    -2,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,     1,     1,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -2,    -1,     1,     0,     0,    -2,    -1,     0,    -1,     0,     0,    -1,     0,    -2,     0,     1,     0,    -1,    -1,     0,     1,     0,    -1,    -3,    -2,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     1,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -1,    -2,     0,     0,     1,     0,     0,    -3,    -1,     0,     0,     0,    -1,    -1,     1,     1,     1,     0,     0,     0,    -2,    -1,    -1,    -2,    -2,    -1,     0,     1,    -2,    -2,     0,     0,     1,     0,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     1,    -2,    -1,    -3,    -2,    -1,    -1,     1,     0,    -1,     1,     1,     0,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     1,    -1,    -1,    -3,    -2,    -2,    -1,    -1,    -1,    -2,     1,     1,     1,     0,     0,    -3,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     1,    -1,     1,     0,     0,    -1,     1,    -1,     0,    -1,    -1,    -2,    -2,    -1,     2,     1,     1,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     1,    -1,     0,     1,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,     1,     0,     1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     1,     1,     1,     0,    -1,     0,     2,     1,     1,     0,     0,    -1,    -1,     1,     1,     0,    -1,     0,     1,    -1,    -2,     0,    -1,    -1,     0,     0,    -1,     0,     0,     2,     2,     2,    -1,     0,     1,     3,     1,     0,    -1,     0,     0,     0,     1,    -1,     0,    -1,     0,    -1,    -1,     1,    -1,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,    -1,    -1,     1,     2,    -1,     0,     0,     0,     0,     2,     1,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     2,     0,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     2,     0,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -3,    -3,    -3,    -2,     0,     1,     1,    -1,     0,    -1,     1,     0,     1,     2,     0,     2,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,     0,     2,     0,     0,     0,    -1,     0,     1,     1,     1,     2,     1,     2,     1,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     1,     2,     0,    -1,    -1,    -2,     0,     2,     2,     2,     2,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -1,     0,     0,     2,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    90 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     1,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     1,     0,     0,     1,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     1,    -1,     1,     1,     0,     1,     0,    -1,    -1,     0,     1,    -1,     0,    -1,     0,     1,     0,     0,     1,     1,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     1,     1,     1,    -1,     0,    -1,    -2,    -2,    -2,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -2,    -2,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     2,     1,     0,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,     1,     0,     1,    -1,     0,     0,     0,    -1,     1,     1,     1,     1,     1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -1,     0,     1,     0,     0,     0,    -2,     0,     0,     0,     0,     0,     2,     1,     1,     1,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -2,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,    -1,     0,     0,    -1,     0,     1,     1,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0),
		    91 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     2,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     1,     1,     3,     2,     1,     1,     1,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     2,     1,     0,    -1,    -2,     1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     2,     2,     2,     0,    -1,     1,     1,     1,     1,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,    -2,    -1,     1,     1,     1,    -1,    -1,    -1,     0,     0,     1,     1,     2,     2,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,     1,     1,     2,     1,    -1,    -1,    -1,     0,     0,    -1,     0,     2,     1,     1,     0,    -1,    -1,     0,     0,     1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,     1,     2,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,    -2,    -1,     2,     2,     1,     0,     0,    -1,    -2,    -1,     0,    -2,     0,     1,     2,     2,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,    -2,    -1,     2,     0,     1,     0,    -1,    -1,    -1,    -2,    -1,    -1,     1,     1,     1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     2,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -2,     0,     0,     1,     1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     1,     0,    -1,     1,     0,     0,     0,     0,    -1,    -2,    -2,     0,    -1,     0,     0,     1,     1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -2,     1,    -1,     0,     0,    -1,     0,    -1,     1,     0,    -2,    -1,     0,    -1,     0,    -1,     1,     1,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     1,     2,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -1,     1,     1,     1,     0,     0,     0,    -2,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -3,    -3,    -1,     1,     1,    -1,    -1,     0,     0,    -2,    -2,    -1,    -2,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     1,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,     0,     1,     0,     1,    -1,     1,     0,     1,     1,     1,     0,     0,    -2,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     2,     1,    -1,    -2,    -1,     1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,     0,     2,     2,     3,     2,     2,     0,    -2,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     1,     3,     1,     1,    -1,     0,     0,     0,     0,    -1,     1,     1,     2,     2,     1,     1,     1,     0,    -1,     0,     1,     0,     1,     0,     0,     0,     2,     2,     2,     1,     1,     0,    -1,     0,     1,     1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     1,     1,     0,     1,     0,     0,     1,     0,     0,     1,     0,    -1,    -1,    -1,     1,     0,    -1,    -2,    -1,    -1,    -2,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     2,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -2,     0,    -2,    -1,    -1,    -1,     1,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     1,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    92 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,    -1,     0,     1,     1,     0,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     2,     2,     2,     0,     1,     2,     3,     2,     1,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     1,     1,     2,     0,    -1,    -2,    -3,    -4,     0,     0,     0,     0,    -1,    -3,    -2,    -2,     0,     0,    -2,    -2,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     3,     2,     2,     3,     1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,    -2,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     2,     1,     1,     0,     0,     0,     1,     0,     0,     0,     1,     1,     1,     2,    -1,    -1,    -2,     1,    -3,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     1,     0,    -1,    -3,     0,    -2,    -1,     0,     0,     1,     0,     1,     3,     1,     0,     1,     0,    -2,    -1,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     2,     1,    -2,     0,     1,    -2,    -1,    -1,     2,     1,     0,     0,     2,     1,    -1,     1,     0,    -1,     1,     1,     0,     0,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,    -1,    -3,    -1,     0,    -1,     0,     1,    -2,     0,     0,    -1,     0,    -1,     0,     1,     1,     1,    -1,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,    -1,    -3,     0,    -1,     0,     0,    -1,     1,    -1,     2,     2,     0,     0,    -1,     1,    -1,     0,     0,     0,     0,    -1,     2,    -1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     1,     1,     0,     1,     1,     0,    -1,    -2,     0,    -1,     0,    -1,     0,     0,     1,     0,    -2,    -1,     1,     1,    -1,    -1,     0,    -1,    -2,     0,    -1,     0,     2,     1,     0,     1,     0,    -2,    -1,    -1,    -2,    -1,    -1,    -1,     1,     2,    -1,     1,     1,    -1,     2,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,     4,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,     1,     3,     2,     2,     2,     0,     0,     0,    -1,     0,     1,     1,     2,     2,    -1,     1,     0,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,    -2,     1,     2,     4,     3,     2,     2,     1,     0,    -1,     2,     2,     0,     1,     1,     1,     1,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     1,     1,     1,     1,     0,     1,     3,     2,     0,     0,     2,     2,    -1,    -1,     0,     2,     1,     2,     1,     0,     1,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     4,     4,     2,     0,     2,     3,     2,     0,     0,     2,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     1,     5,     3,     1,     1,     1,     1,     1,     0,     0,     0,     1,    -1,     0,     0,    -1,     1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     1,     4,     3,     3,     2,     2,     1,     0,     1,     0,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,     1,     1,    -1,    -1,     0,     1,    -1,    -2,     1,     2,     3,     3,     2,     1,     0,    -1,     0,     2,     0,    -1,     2,    -1,     0,     0,     0,     0,     0,     1,     1,     2,     0,     0,    -1,     0,    -1,     0,     1,     3,     3,     4,     2,     1,     1,     0,     0,     0,     0,     0,     2,    -1,     1,     0,     0,     0,     1,     2,     1,     0,     1,     1,    -1,     0,     0,    -1,     3,     5,     3,     3,     4,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,    -1,     0,     1,     1,     0,     1,    -1,     0,    -1,    -1,     0,     1,     4,     4,     4,     3,     3,     1,    -1,     1,     0,     0,     0,     0,     0,    -2,     0,     1,     1,     0,     1,     2,     1,     1,     0,     0,    -1,    -1,     3,     5,     4,     3,     4,     3,     2,     2,    -1,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -2,     1,    -1,     0,     1,     1,     1,    -2,    -3,     0,     0,     3,     4,     5,     4,     2,     3,     2,    -1,     1,     0,     1,     0,     0,     0,    -1,     0,    -2,    -3,     1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,     0,     1,     0,     2,     3,     1,     0,     1,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -2,    -4,    -4,    -3,    -3,    -4,    -4,    -3,    -3,    -3,    -3,    -4,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0),
		    93 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     2,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,    -1,    -2,    -2,    -2,    -2,    -3,    -4,    -2,    -2,    -2,    -2,    -2,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     2,     2,    -1,     0,    -2,     0,    -1,    -1,    -2,    -3,    -3,    -3,    -3,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     2,     0,    -1,     0,     1,     1,     1,     1,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -1,     0,    -2,    -1,     0,     0,     0,     0,     1,     1,    -1,     0,     1,     0,     1,    -1,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     1,     0,     1,     0,     0,    -1,     0,     0,     0,     1,    -1,    -2,    -3,    -3,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,     0,     0,    -2,     0,     2,     2,     2,     1,     0,    -3,    -3,    -3,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     1,    -1,    -1,    -1,     0,    -1,     1,     2,     2,     2,     0,    -1,    -4,    -3,    -3,    -2,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     2,     0,     1,     0,    -1,    -1,     0,     0,     1,     1,     1,     0,    -1,    -2,    -4,    -4,    -3,    -3,    -2,    -1,     0,    -1,    -1,     0,     0,     0,    -2,     0,     2,     1,     0,     0,     0,     0,     1,     1,     1,     1,     0,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,    -2,    -2,     1,     0,     0,    -1,    -1,     1,     1,     2,     1,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     2,     1,    -1,    -1,    -1,     0,     0,    -1,    -1,     2,     1,     0,     0,    -1,     1,     1,     1,     1,     1,     1,     0,    -1,     0,     0,     1,     0,     0,     0,     1,     1,     1,    -1,    -1,     0,     0,     1,     0,     1,    -1,    -1,    -1,    -1,     0,     1,     1,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     0,     0,     0,     3,     1,    -2,    -1,     0,     0,     1,     0,     0,    -2,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     2,     1,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -2,     0,     1,    -1,    -1,    -1,    -2,    -3,    -1,    -1,    -1,     0,     0,     1,     2,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -1,    -1,    -2,    -1,    -1,    -1,    -3,    -2,    -1,    -1,    -2,     1,     1,     2,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -3,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     1,     1,     1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     1,     0,     0,    -1,    -1,     0,     1,     0,    -1,     0,     1,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,     0,     1,     1,     0,     0,     0,     1,     1,     1,     1,     0,    -1,     0,     1,     1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,    -1,     1,     1,     1,     0,     0,     2,     0,    -1,     0,     0,    -1,    -2,    -1,     0,    -1,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,     1,     1,    -1,    -1,    -1,     0,     0,    -2,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    94 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -2,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -1,     0,    -1,    -2,    -1,    -2,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -2,    -3,    -1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -3,    -2,    -1,     1,    -1,    -2,     0,     0,     0,     0,     1,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,     0,     0,    -1,    -2,     0,     1,    -1,    -1,    -2,    -1,    -1,    -1,     1,     1,     1,     0,    -1,    -2,     0,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,     0,     1,     0,     2,    -1,     0,    -1,    -2,    -2,    -1,     0,     3,     1,     0,     1,    -1,    -1,    -2,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -2,    -1,    -1,     0,    -3,    -4,    -1,     0,     1,     2,     3,     3,    -1,    -1,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     2,     0,    -1,    -2,     0,     1,    -1,    -3,    -3,     0,     1,     1,     1,     1,     1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     1,     0,    -1,     0,     1,     1,    -1,    -2,    -1,     1,     0,    -1,    -2,    -2,    -2,     3,     0,     1,     0,    -1,    -2,    -2,    -2,    -1,    -1,    -1,     0,    -1,     1,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,     0,    -1,     0,    -1,    -2,     0,     2,     1,     0,     0,     1,     0,    -2,    -2,     0,     0,    -1,     0,    -1,     1,     1,     0,    -1,    -1,     0,     0,    -1,     1,     0,     0,     0,    -2,    -3,    -1,     1,     0,     0,    -1,     1,    -1,    -3,    -2,     0,     0,    -1,     0,    -2,    -1,     1,    -1,     0,     0,    -1,     1,     0,     1,     1,     0,    -1,    -3,    -2,     0,     1,     0,     0,    -1,    -2,    -2,    -2,    -3,    -1,     0,    -1,     0,    -1,     0,     0,    -1,     0,     1,     0,     0,     0,     1,     1,     1,    -2,    -2,    -2,     0,     0,     0,     0,    -1,    -2,    -2,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,     0,    -2,    -2,    -2,    -1,     1,     1,    -1,    -1,     0,     1,     1,    -1,    -1,    -2,     0,     0,     0,    -2,     0,     2,     1,     0,     1,     0,     2,     2,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     3,     0,     2,     0,     0,     0,     0,     0,     1,     1,     1,     0,    -1,    -2,    -1,     0,     0,     1,     0,     1,     2,    -1,    -2,    -2,    -1,     0,     0,     0,     0,    -2,    -1,    -1,     1,     0,    -1,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     1,     0,     1,     0,     0,    -2,    -1,    -1,    -2,    -1,     0,     0,     1,    -2,     0,     0,     0,     1,     1,     0,     0,     0,    -2,     0,     0,     1,     0,     0,     1,    -1,     0,     1,    -1,    -1,    -2,     1,     0,    -1,    -1,     0,     1,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,    -2,     0,     1,     1,     0,     1,     0,     1,     1,     0,    -2,     0,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,    -3,    -3,    -1,     0,     2,     0,    -1,     1,     1,     1,     1,    -1,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,     1,     1,     1,     1,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -2,     0,     0,     0,     0,     1,     1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     1,     1,     0,     1,     1,     1,    -1,     1,     0,    -1,     0,     0,     0,     0,    -2,    -2,     1,     0,     0,    -2,    -2,    -4,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     1,     1,     0,     0,     0,     2,     1,     0,     0,     0,     0,    -1,    -2,    -1,     0,    -1,     0,    -2,    -3,    -2,    -1,    -1,     0,     0,     1,    -1,     0,     1,     1,     2,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,    -2,    -1,     0,    -1,     0,    -1,     0,     0,    -2,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,    -3,     0,     0,     0,    -2,    -3,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -3,     0,    -1,    -2,    -3,    -2,    -3,    -2,    -2,    -2,    -3,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -1,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0),
		    95 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     1,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,     0,     0,     1,     0,     1,     2,     2,     1,    -1,    -1,     2,     0,     0,     1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     1,     0,    -2,     1,     0,     1,     1,    -1,    -1,     0,     0,    -1,     0,     1,    -1,     0,     1,     1,     3,     3,     1,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     2,     2,     0,    -1,    -2,    -1,     0,     1,     0,     1,     0,     0,     1,     1,     1,     2,     2,     2,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     2,     0,     1,    -2,    -1,     0,     1,     2,     1,     2,     1,     0,     0,     1,     2,     0,     1,     1,     2,     0,     0,     0,     0,    -1,     0,     0,    -1,     1,     1,     1,     1,     0,    -2,    -1,     2,     1,     2,     2,     1,     0,     1,     0,    -1,    -1,    -1,     1,     1,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     2,     2,     1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,    -1,    -1,     2,     0,     0,     0,    -2,    -2,    -1,     0,     0,     0,     1,     1,     1,     1,    -2,    -3,    -3,    -4,    -4,    -6,    -3,    -4,    -4,    -4,    -2,    -2,    -2,    -1,     2,     1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     1,     1,     0,    -1,    -2,    -3,    -3,    -2,    -2,    -5,    -5,    -4,    -5,    -5,    -5,    -2,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,     0,    -1,    -1,     0,     1,     1,     0,    -1,    -1,    -3,    -3,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,     1,     0,     1,     0,    -1,    -1,    -1,     1,     1,     1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     1,    -1,    -1,     0,     1,     0,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     2,     1,     1,     0,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     2,    -1,    -2,    -1,     0,     1,     0,    -2,    -1,    -2,     1,    -1,     0,     0,     1,     1,    -1,    -1,    -1,    -1,     0,    -2,    -1,     0,     0,    -1,     0,     0,     2,     0,    -1,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -2,     0,     0,    -1,     1,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     1,     0,     1,     1,     0,     0,     0,    -2,    -2,     0,     0,     1,     2,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -3,    -2,    -1,    -1,     0,     0,     0,     1,    -1,    -1,     0,     0,    -3,    -2,     0,     0,     2,     2,     1,     0,    -1,    -2,    -3,    -1,    -1,    -2,    -1,    -3,    -2,    -2,    -2,     0,     1,     1,     1,     1,     0,    -1,     2,     0,     0,    -2,     0,     0,     1,     1,     1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     1,     0,     1,     1,     1,     0,     0,     0,     0,    -1,     0,    -2,     0,     0,     0,     0,     1,     1,     0,     0,     0,    -1,    -2,     0,    -1,     0,     0,    -1,     1,     1,     2,     0,     0,     0,     1,     1,     2,     1,     2,     0,     0,     0,     0,    -1,     1,     0,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     3,     1,     3,     2,     0,     0,     0,     1,     1,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     1,     0,     1,     1,     1,     2,     3,     0,     0,     0,     0,     1,     2,     1,     1,    -1,     0,     1,     0,    -1,     0,     1,     1,     1,    -1,     0,     0,     0,     0,     1,    -1,    -2,     0,    -1,     0,     0,     0,     0,     0,     2,    -1,    -1,     2,     1,     2,     2,     1,     0,     2,     1,     1,     1,    -1,     0,     1,     2,     2,     1,     2,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     1,     0,    -3,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0),
		    96 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     1,     2,     1,     1,     1,     2,     3,    -1,     1,     1,     2,     2,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     2,     1,     1,     1,     1,     1,     2,     3,     2,     1,     1,     1,     2,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     3,     0,     0,     2,     3,     1,     1,     2,     0,     1,     2,     2,     1,     0,    -1,    -1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     3,     0,     2,     2,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,    -1,    -3,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -1,     1,     1,     0,    -1,    -1,     0,     1,     0,     1,     0,    -2,     0,    -2,    -1,    -1,    -2,    -3,    -3,    -3,    -2,    -1,    -1,     1,     1,     0,     0,     0,    -2,     1,     0,    -1,    -2,    -2,     2,     1,     1,     1,     0,    -1,    -2,    -2,    -2,    -4,    -4,    -2,    -4,    -3,    -3,    -2,     0,     0,    -1,     0,     0,     0,    -2,     1,     0,    -2,    -2,     0,     0,     1,     1,     0,     0,    -1,    -2,    -3,    -3,    -4,    -3,    -2,    -1,    -4,    -3,    -3,    -1,     1,    -1,     0,     0,     0,    -2,     1,     0,    -1,    -1,     1,     1,     0,     0,    -1,     0,    -3,    -5,    -4,    -2,    -2,     0,     0,     1,    -1,    -2,    -2,    -2,     0,    -2,     0,     0,     0,     0,     1,     0,    -1,     0,     1,     0,     0,     0,     0,    -3,    -2,    -2,    -1,     0,     0,     2,     2,     2,     1,     1,     0,    -2,    -1,    -1,     0,     0,     0,    -1,     1,     1,    -1,     0,     1,    -1,     0,     0,     0,    -4,    -2,     0,     0,     2,     1,     1,     1,     1,     0,     0,     1,    -1,    -2,    -2,     0,     0,     0,    -1,     1,     1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -3,    -2,     0,     1,     1,     1,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     1,    -1,     1,     0,     1,     1,     1,     1,     1,     1,     1,     1,    -1,    -1,     0,     0,    -1,    -2,    -1,     1,     1,    -1,     0,     0,     0,    -2,    -2,    -1,     0,     0,     1,     0,    -1,     1,     0,     1,     1,     2,     2,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     1,    -1,     1,     0,     1,     0,    -1,     0,     0,     1,     0,     0,     1,    -1,     1,     0,     1,     2,     0,     3,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,    -1,     1,     1,     0,     0,     1,     2,     0,    -2,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,     0,     1,     1,    -1,     0,     1,     0,     0,     0,    -2,     0,    -1,     0,    -1,     0,     1,     2,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -1,     0,    -2,     0,    -1,     0,     2,     2,     0,    -1,     0,     0,     0,    -1,     1,    -1,    -2,     1,     0,    -1,    -2,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,    -1,    -1,     0,     0,     0,    -1,     1,    -1,    -1,     0,     1,     0,     0,    -2,    -2,    -1,     1,     1,     1,     0,    -2,    -1,     0,     0,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,     1,     0,    -2,     0,    -1,     0,     0,    -1,    -2,    -1,     1,     3,     1,     1,     1,    -1,     1,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,    -1,    -2,     0,     1,     1,     0,     1,    -1,    -2,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,    -2,    -3,    -2,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -3,    -3,    -3,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -3,    -2,    -2,     0,     0,    -2,    -4,    -4,    -4,    -2,    -1,    -2,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -2,    -2,    -3,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    97 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,    -3,    -3,    -2,    -3,    -3,    -3,    -3,    -2,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -3,    -4,    -4,    -4,    -2,    -2,    -2,    -2,    -1,    -3,    -2,    -2,    -1,    -2,    -1,    -2,    -3,    -3,    -2,    -1,     0,     0,     0,     0,    -2,    -4,     1,    -2,    -1,     0,     1,    -1,    -1,     0,     1,     1,     0,     1,     0,     0,    -2,    -3,    -2,    -1,    -4,    -3,    -3,    -2,     0,     0,     0,     1,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     1,     1,     0,    -1,     0,     0,     2,     1,     1,    -1,    -3,    -2,    -2,    -1,     0,     1,     2,     1,     1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     0,     1,    -1,    -1,     2,     0,    -1,     0,     0,     0,    -1,     0,    -2,    -3,    -1,    -1,     3,     1,     0,     1,     0,    -1,     0,     1,     1,     1,     1,     0,    -1,    -1,     0,     0,     1,     1,     0,     1,     0,    -1,    -1,    -1,    -3,    -4,    -1,     0,     2,    -1,     0,     1,     1,     1,     0,     1,     2,     2,     0,    -1,    -1,     1,     1,     0,     1,     1,     0,     1,     0,     1,    -1,    -1,     0,     0,     3,     0,     1,     1,     0,     1,     1,     0,     1,     2,     1,     1,    -1,    -2,    -1,     1,     2,     1,     0,     1,     0,     1,     0,     0,    -1,    -1,     1,     0,     3,     0,     0,     2,     1,    -1,     0,     0,     1,     1,     1,    -1,    -1,     1,     2,     3,     2,     1,     0,     1,    -1,     1,    -1,     0,     1,     0,    -2,    -1,     2,     0,     1,     2,     0,    -1,    -1,     0,     0,     1,     0,     1,     2,     1,     1,     3,     2,     2,     1,     0,    -1,     0,     0,     2,     0,     1,     1,     1,     2,     0,     0,     2,     0,    -2,    -1,     0,     0,     0,     1,     0,     1,     1,     1,     3,     2,     1,     1,    -1,    -1,    -2,    -1,     0,    -1,     0,     1,     0,    -1,     0,     1,     1,    -1,    -2,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     2,     0,     1,     1,    -1,    -1,    -1,    -2,    -1,     0,     1,    -1,    -2,     0,     0,     0,     0,    -1,    -2,     0,     0,    -1,    -2,    -2,    -1,     0,    -1,     0,    -1,    -1,     0,     1,     2,     0,     0,     0,     2,     1,     1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     1,    -1,    -2,    -1,    -1,     0,    -1,     2,     3,     3,     1,     2,     1,     2,     2,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     0,     0,     2,     2,     3,     1,     2,     1,     2,     2,     0,     1,     0,    -2,     0,     0,     1,    -1,     0,     1,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     3,     2,     1,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     1,     1,     0,     1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     2,     3,     1,     1,     0,     1,     0,     0,     1,     0,    -1,     0,     0,     1,     0,    -1,    -2,     0,     0,     1,     1,     0,     0,    -1,    -1,     0,     0,     1,     0,     1,     0,     0,     0,     0,    -1,    -1,     1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     1,     1,     1,     1,     1,     1,     0,     0,     0,    -1,     1,     0,    -1,    -2,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     1,     2,     1,     0,     0,     1,     0,     1,     0,     0,    -1,     0,    -2,    -1,    -1,    -2,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,    -1,    -2,    -1,     1,     2,     1,     1,     0,     1,     0,    -1,     0,    -2,    -2,    -1,    -2,    -2,    -2,    -1,    -1,    -3,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -3,    -2,    -2,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     2,     0,     0,     0,     0,    -1,     1,     1,     0,     0,     0,    -2,    -2,     0,    -1,    -2,    -3,    -2,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -1,    -1,     0,     2,     0,    -1,     0,     0,     0,     0,     0,    -2,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     2,     1,    -1,     0,     1,     0,     1,     0,     0,     0,     0),
		    98 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,     1,     1,     2,     1,     2,     2,     1,     1,     0,     1,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,     0,     1,     1,    -1,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -3,    -1,     1,     1,    -1,     0,     0,    -2,    -1,     1,     0,     0,     1,     1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     3,     1,     1,     1,     0,     0,     0,     1,     1,     1,     0,    -1,     1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     2,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,     1,     2,    -1,    -1,     1,     1,    -1,    -1,    -2,    -1,    -2,     0,     0,     0,     0,    -1,     0,    -2,     0,     1,     1,     0,     0,     0,    -1,     0,    -2,    -2,     0,    -1,    -1,     0,     1,     2,     1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,     1,     0,    -1,     0,     0,    -2,    -2,     0,     0,    -1,    -1,    -1,    -2,     1,    -1,    -3,    -1,     1,     3,     3,     2,     1,     0,     0,     0,     0,    -2,     1,     1,     0,    -1,    -2,    -3,    -2,    -2,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,     0,     2,     2,     2,     0,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -3,    -3,    -3,     0,     0,     1,     2,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -2,    -3,    -3,    -2,    -2,     0,     0,     1,     0,     0,     0,    -1,    -2,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -1,    -2,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     1,    -1,    -2,    -2,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     1,    -1,    -1,     0,     0,     1,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,     2,     0,     0,    -1,     0,    -2,     0,    -2,     1,    -1,     1,     1,     1,    -1,     0,    -1,    -1,    -3,    -1,     0,     0,    -1,    -2,     1,     0,    -1,     1,     1,     0,    -1,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,     1,     0,     2,     1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     2,     0,     1,     1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -3,    -1,     1,     1,     1,     1,     1,     1,    -2,    -1,     0,    -1,     0,    -1,    -1,     1,     1,     2,     1,     1,    -1,    -1,     0,     0,    -2,    -1,    -1,     0,    -1,     0,    -1,     0,     1,     1,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,    -1,     0,     1,     1,     1,     1,    -1,    -2,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,     1,     1,     0,    -1,    -1,     0,    -2,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     1,    -1,    -1,    -1,    -2,     0,     1,     1,     0,    -1,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -1,    -1,     0,     2,     1,    -1,    -1,     0,     1,     1,    -1,     0,    -2,    -1,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,     1,     0,     1,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     1,    -2,     0,     0,     0,    -1,     0,    -1,    -1,     1,     1,     0,     0,    -1,    -1,     0,     0,     1,     1,     1,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    99 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,     1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     1,     0,     0,     1,    -1,     0,    -1,    -1,    -2,    -1,     1,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -2,    -2,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,     1,     1,     0,     0,     2,     0,    -1,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -2,    -1,     0,    -1,    -2,     1,     1,     0,     1,     0,     1,    -1,     1,     1,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,    -2,     2,     0,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     0,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     0,     0,    -1,     1,     1,     1,     0,     1,     0,    -1,    -2,    -2,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,    -2,    -1,    -1,     0,     0,    -1,     0,     1,     1,     0,     1,     0,    -1,    -3,    -1,     0,    -2,    -2,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,    -1,    -2,    -1,    -1,     0,     0,    -1,    -1,     1,     1,     1,     0,     0,    -2,    -2,    -1,     0,    -1,    -1,    -2,     0,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,    -2,     1,     1,     0,     0,     0,    -1,    -2,     0,    -1,    -1,     0,     0,     0,     0,    -2,     0,     0,     0,     1,     1,    -2,    -2,    -1,     0,    -1,     0,     0,    -1,     1,     2,     1,     2,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     1,     1,    -2,     0,    -1,     0,     0,     0,    -2,     0,     0,     0,     1,     1,     2,     1,     1,     1,     1,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,     0,     1,     0,    -2,    -1,    -1,    -1,     0,     0,    -2,     1,    -1,    -1,     0,     1,     0,     0,     1,     0,     0,    -2,    -1,     0,    -1,    -1,     0,    -2,     0,    -1,     1,     1,    -1,     0,    -1,    -1,     0,     0,    -1,     1,     0,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -2,     1,     0,    -1,    -1,    -1,    -2,     0,    -1,     0,     1,     1,     1,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -2,     1,     1,    -1,    -2,    -1,    -1,     0,     0,     0,     1,     1,     2,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     1,    -1,    -3,    -1,     0,    -1,     0,     1,    -1,     0,     1,     2,    -2,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     2,    -2,    -2,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     1,    -1,     0,     1,     0,    -1,     1,     0,     2,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     1,     1,    -1,     0,     0,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     2,    -1,     0,     1,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,     1,     1,     0,     0,    -1,     1,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     2,     1,     1,     1,     0,     0,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,     0)
        );

 ---------------------------------INFO-
 -- COEF =2.6961303

 -- MIN =-7.9999995
 -- MAX =5.2991276

 -- SUMMIN =-568.40125
 -- SUMMAX =413.2596
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
