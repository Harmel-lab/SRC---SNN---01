----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (   -1,     0,    -1,    -3,    -3,     4,     0,     0,     2,    -3,    -1,     5,    -1,    -8,    -7,     2,    -4,     3,     2,     1,    -5,    -4,    -2,     3,     5,     5,    -1,    -4,    -3,    -4,     0,     1,     1,    -4,     3,     2,     0,     1,    -2,     3,     7,     4,    -7,     5,    13,     6,    -2,    -4,    -4,     3,    -1,     2,     2,    -1,     2,    -4,     3,     5,     1,     5,    13,     1,    -7,     1,    -8,   -21,    -2,    -4,    -2,   -12,   -11,   -18,    -3,    -4,    -7,    -3,    -3,    -3,   -11,    -8,    -7,    -9,     1,    -3,     2,    -5,    -1,    10,    -1,     7,     5,   -15,   -10,    -8,   -14,   -11,   -19,   -12,   -18,   -20,    -6,    13,     1,   -16,   -11,    -8,   -12,    -7,     5,     3,    -3,     3,    -3,     2,     1,    -1,    -7,   -18,     4,   -12,   -26,   -13,   -13,   -20,   -34,    -3,    -1,    -9,    -4,   -18,   -13,   -11,    -2,    -7,   -10,    -7,     2,    -5,    -9,     1,     1,     3,   -10,    -2,     0,    -6,    -4,    -2,    -7,    -5,   -16,   -30,   -18,   -26,     4,    12,    -1,   -12,     1,   -17,   -21,     1,    -3,    -3,    -6,   -23,    -6,    -5,    -5,     5,   -10,    -7,    -7,     0,    -6,    -5,   -10,   -10,    -9,   -32,   -23,    -9,    -3,   -11,    13,    10,     2,   -20,   -17,   -10,     2,   -22,    -9,   -21,    -6,    13,     1,    -9,    -8,    -8,     3,    -4,    -6,     4,    -8,    -9,   -21,   -33,   -32,   -12,    -1,     0,    21,    11,   -20,     0,   -19,   -16,     6,   -12,   -19,    -7,   -20,    13,    15,   -26,    14,     9,    -3,    -4,    -6,    -1,    -4,   -18,   -11,   -32,    -7,    -6,     8,   -11,     5,    23,   -10,     4,   -20,   -25,    -6,   -14,    -7,   -26,    -9,    -6,    -6,    -4,    23,    -2,    -2,    -2,   -16,    -2,   -12,   -30,   -12,    -3,    -7,     8,    -5,    -8,    16,     4,     0,   -16,   -38,    -4,    -2,    -9,   -12,   -20,     0,     4,    -6,    -5,     6,     9,   -10,   -12,    -6,     8,     0,    -3,   -10,    -7,    -4,    -1,   -23,   -25,    -8,   -17,     5,   -17,   -17,    -6,   -15,   -18,    -8,    -7,   -18,     2,     2,    22,   -10,     4,   -12,    -2,    -4,    -2,    -8,    -6,   -15,     2,    10,    -8,    -9,     2,   -13,     4,    30,   -21,   -17,     3,   -15,   -25,    -9,   -14,   -10,    -4,    -2,     7,     4,     0,    -1,     5,     1,     0,   -24,     0,     3,    -5,    11,    -5,   -10,   -25,     3,    15,    25,    -5,     1,    15,     0,   -26,   -17,   -16,   -13,     3,    -1,    11,    12,    -5,     0,     2,    11,   -15,   -13,     2,    -5,   -19,     6,   -17,   -46,   -37,    -3,    13,    22,     6,    -3,    17,    -8,   -15,   -11,    -6,   -20,     1,    -2,     0,     1,    -7,    -5,     9,   -11,   -15,   -12,    -3,     5,     9,    20,    -3,   -32,   -34,    -2,     4,    10,     7,   -18,     1,    -2,    -9,   -13,     3,   -16,    -1,     0,    -4,   -10,    -8,     4,   -16,    -1,   -25,   -13,   -21,    -5,     9,    27,     6,   -42,   -13,    -5,     6,    -2,    -7,   -18,    15,   -14,   -11,     1,   -10,   -12,    -2,    -4,     1,    -5,   -13,     4,     1,   -29,    -9,   -19,   -22,   -12,    12,    13,   -13,   -50,    -1,    -5,    33,   -10,    -6,   -14,   -12,     0,   -12,   -13,    -9,   -28,    12,     0,     2,   -17,    -9,   -22,    -6,   -15,   -14,   -16,   -39,     5,     6,    16,   -11,   -36,   -13,    -1,    17,     6,     0,     9,   -11,    -6,     6,   -12,   -15,   -27,    10,     1,     2,    -7,     5,    -7,   -13,    -6,    -3,   -13,   -20,    14,    14,   -13,   -21,   -42,    -5,    -2,     2,    -6,     1,     0,    -4,     5,   -10,     0,    -2,   -12,    -6,     4,     9,     2,     6,     3,   -11,    -5,   -20,   -15,     4,    11,    13,     0,   -22,   -24,    16,     5,   -14,   -10,     0,   -19,    -8,    -9,    -8,     2,   -36,    -7,    -5,    -2,     0,    -4,    -9,     4,    -4,   -13,   -25,   -20,     6,     2,   -13,   -16,    -5,    -5,     4,     6,   -12,    -1,   -22,   -14,   -16,    -4,    -4,    -6,    -7,     4,     5,     1,    -2,   -12,   -13,    -6,    -6,     1,   -16,    -9,    -6,     5,    -5,     0,    -4,    -4,    10,    -5,    -5,   -14,   -20,   -19,   -11,     3,     2,   -18,     1,     8,     7,    -1,     2,   -10,   -29,     3,     2,     6,     1,   -10,     7,     3,    10,    -4,   -21,    17,    14,    15,   -30,   -12,   -16,   -14,   -10,     3,    -4,    -1,    -5,     7,     2,     2,     2,   -11,   -22,   -10,     4,    -8,    -2,   -10,   -22,    12,     7,    10,    14,   -15,   -14,   -17,   -36,     0,   -22,   -14,    -7,    10,    -1,    -8,   -20,   -11,    -4,     4,    -5,    -5,     1,   -13,    13,     6,     4,   -22,   -26,   -16,   -17,     3,    25,     5,     5,   -22,    -8,    -5,   -17,   -15,     8,    -9,   -12,    -1,    -3,    -5,     2,     1,     4,     2,    -3,   -36,   -14,   -13,   -13,    -6,   -13,   -22,   -25,   -37,   -34,   -42,   -17,   -11,   -13,   -14,   -10,   -18,    -7,   -12,    -9,    -1,     1,    -2,     0,     1,     3,    -4,    -2,    -3,   -17,   -26,     3,    -1,   -16,    -9,    -5,   -13,   -11,   -12,   -12,    -6,   -18,   -27,   -12,   -20,   -12,    -5,     0,    -5,    -3,    -4,     1,     2,    -5,    -1,    -4,    -1,     3,     2,    -1,    -2,    -5,     3,    -2,     2,   -12,     3,     0,    -7,     1,     5,     1,    -3,    -7,    -6,   -10,    -2,     1,    -5,     3),
		     1 => (   -1,    -3,    -1,     5,     1,    -2,     1,    -2,     4,    -4,     2,    -4,    -2,    -5,     2,     3,     1,     2,    -3,     2,    -5,    -3,     4,    -3,     0,     2,    -4,     4,     5,     5,     4,     4,    -5,     5,     1,     2,    -5,    -2,    -2,    -4,    -8,    -5,    16,    12,    -1,    -8,    -5,     4,    -5,    -4,    -1,    -3,    -4,     4,    -2,     4,     3,     1,     0,     4,     1,    -1,     4,     2,   -14,   -14,     0,    -4,    -4,    -5,    -8,   -17,   -19,   -23,   -28,     3,     9,   -25,    -7,    -1,    -4,    -7,     2,     4,     4,    -4,    31,    22,    -1,     3,     5,    25,    20,    13,    13,     7,     3,   -37,   -38,   -39,   -33,    -9,   -10,    -3,     4,   -20,     9,     2,   -13,    -1,     3,     4,     0,    -1,    21,    18,     9,    -6,    -4,     0,     0,    -4,   -14,   -35,   -34,   -41,     4,    17,     2,     3,     6,     8,     5,     9,   -10,   -42,   -22,   -35,   -21,   -20,     1,    -5,    20,    28,     9,     2,    -9,   -10,   -48,   -21,   -18,   -30,   -41,   -23,    -3,    29,    -2,    -3,    -1,    10,    12,   -12,   -17,   -40,   -30,   -22,   -21,   -17,    -2,    -2,     0,    11,    10,    -9,    -1,     4,   -39,     3,     3,   -30,   -31,   -16,   -23,    -9,    -2,     9,    -1,    11,   -11,   -13,    -7,   -42,   -29,   -11,    -2,    -6,    -4,    -1,    -9,     9,     5,     1,    -8,   -16,   -43,   -10,   -22,   -35,   -26,    -5,    17,     7,     8,    -3,    19,    -4,   -16,   -11,     0,   -26,   -28,   -12,   -12,    -9,     0,    -6,    -6,    -6,    -4,    -6,   -14,   -16,   -30,   -27,   -13,   -49,   -45,     1,    11,     9,    17,    11,     6,   -10,   -17,    -9,   -15,   -25,   -29,   -16,   -16,    -3,     4,    -1,    -6,     7,    -6,     1,   -23,   -11,    -9,   -14,   -35,   -64,   -15,    -3,    -8,     0,    20,     4,   -20,   -14,   -29,   -11,    -7,   -16,   -27,   -14,     1,   -16,     1,     6,    -3,    -7,    -3,    -3,   -20,   -26,   -17,   -23,    -3,   -33,   -26,   -13,     4,    24,    20,    -3,   -20,   -18,   -26,   -10,   -10,   -13,   -28,   -31,    -1,    33,     1,    -1,     5,     8,     9,     2,   -13,   -15,   -26,   -42,   -22,   -35,   -10,   -14,    -1,    30,     2,   -26,   -15,    -8,    -9,     5,    -8,   -17,   -31,   -28,    -2,    28,     1,     1,    -9,    22,     5,    -6,    -8,    -6,   -40,   -34,   -20,   -19,     1,    -9,    20,    -4,    12,   -41,   -44,   -15,    19,    26,    27,    18,    -8,     0,    -4,    17,     2,    -4,    -1,     7,    11,    -8,   -10,    -3,   -20,   -46,   -21,   -11,    -7,     6,    23,    -9,     8,   -38,   -44,     4,    17,     2,    -2,   -34,   -19,     1,     9,     3,    -4,     4,    11,    10,    13,   -25,   -15,   -10,    -5,   -29,   -20,     8,    -4,   -16,    23,     1,   -17,   -38,    -3,    23,    26,    32,    18,   -10,   -15,    31,    30,     1,     4,     2,    12,    29,    12,    -3,    -7,    -3,    17,     2,    -7,    17,     1,   -10,    -9,   -24,   -18,   -30,   -11,   -24,    -4,    35,    14,   -18,   -41,    10,     6,    -3,     2,     4,     4,   -13,   -10,    -3,     7,     2,    17,    11,     9,    20,     8,     9,   -16,    -8,    -6,   -36,   -30,   -32,    -3,    26,    17,    32,    39,   -10,    -7,    -2,     3,    -3,     6,   -14,     5,     2,    15,     5,    12,     4,     5,     8,    -3,     6,     7,    -8,   -16,   -12,     7,    14,    18,    30,    33,    37,    23,    -1,    -6,   -14,   -11,    -2,    -1,    -9,   -10,   -12,   -14,    -6,     5,   -16,     5,    -8,    -3,    12,   -18,   -38,   -30,     7,    19,    22,    13,     3,     3,    -1,    11,    20,     3,    14,    -2,    -4,    16,    16,   -19,    15,    19,     5,     2,   -17,    -4,     9,     8,    11,   -23,   -28,   -43,    -7,    13,    -4,    -4,    -7,   -22,     2,    21,    27,     6,    14,    -1,    -3,    17,     5,     0,    27,    11,   -17,    -1,    -7,   -18,     7,    -1,    11,   -12,   -32,   -36,    -9,   -10,    -4,    21,   -22,   -13,     0,    10,    10,    11,     0,    21,    14,    -6,    -2,     1,   -22,   -36,   -12,     1,    -7,     1,    -6,    10,   -15,     0,    -8,   -31,   -33,   -27,    -9,    12,     7,     7,    10,    14,    14,     3,     3,    15,    17,     2,     0,     2,   -19,   -43,    -8,    -1,   -11,     8,   -12,    -3,    -5,    12,   -14,   -10,   -27,     3,    19,    30,    11,    19,    14,    17,    26,    41,     5,    -4,    -4,    -5,     2,   -15,    -3,   -14,   -17,    17,   -10,    -5,    10,     0,     2,     8,    -3,     5,     5,     9,    25,    30,     2,    -2,    -7,    13,    20,    39,    -2,     0,     2,    -4,    -6,   -13,   -22,    -7,   -19,   -12,   -19,   -34,   -10,   -16,   -38,    14,    12,    -5,     6,     4,    50,    34,     5,    -3,     5,    -9,     7,    10,    -1,     3,     3,    -1,    -2,     0,    -2,    -3,    -5,   -17,    10,   -33,   -18,   -27,   -22,   -23,   -37,   -14,   -21,   -14,   -16,   -20,   -17,   -10,    -9,    -6,     1,    -5,     4,    -2,    -4,    -2,    -4,    -9,   -17,   -21,   -11,   -13,   -16,     6,    -3,   -27,   -25,   -34,   -35,   -27,   -19,    -4,    -9,    -5,    -4,    -1,     3,    -5,     2,    -4,     1,    -2,    -1,    -5,     3,     4,     2,    -3,    -2,    -3,    -4,    -5,    -7,     3,     3,     6,    -2,    -3,    -2,    -5,    -4,     0,     2,    -4,     4,     5,     1,     3,     3),
		     2 => (    0,    -4,     2,    -4,    -4,     2,     3,     2,     0,     4,     1,    -5,    -1,     1,     0,     2,     1,    -5,    -2,     1,     1,     3,     0,     2,     1,    -4,    -2,    -2,     0,     3,     0,    -1,     4,     3,    -4,     4,   -10,   -14,   -10,    -8,    -4,   -22,   -16,    -6,    -1,     6,    -1,    -5,    -6,    -3,    -4,    -9,     2,     2,     5,     3,     2,    -4,     1,   -13,   -15,     1,     4,   -26,    -7,   -11,   -11,   -19,   -10,   -50,   -15,    -3,    -8,   -12,   -21,   -25,   -19,    -4,   -11,     2,     6,    11,     3,     4,    -2,     4,    -8,   -21,   -20,    -1,    22,    -9,    -3,    21,    21,     3,   -22,   -28,   -16,   -28,   -26,   -10,    13,    -9,   -29,   -17,    -3,   -11,   -14,     6,    -4,    -4,    -4,     5,    -2,    12,    -7,   -13,    -3,    21,     5,    -2,   -21,   -16,   -13,   -31,   -32,   -21,     8,     8,     2,   -10,    11,    16,    -4,   -24,     4,     3,   -13,    -5,     0,     4,    -7,     3,    26,     6,    -1,    -1,    -5,    -8,   -24,   -34,   -36,   -34,   -27,   -13,    -5,     3,    16,    18,    13,    21,     5,   -18,   -15,     1,   -14,    -3,     5,     5,     8,     2,     4,    -6,    -7,    12,     6,    -8,    -9,   -13,    -6,   -35,   -27,   -23,   -13,    21,     8,    15,    -6,     6,     3,   -28,   -24,    24,   -15,    -3,     3,     3,    21,     1,    -1,   -13,    -2,    14,    -2,     5,     0,    10,     7,    15,   -13,   -13,   -11,    -8,   -27,    -7,     9,     6,     3,   -47,    -6,    34,   -17,    -2,   -26,    24,    22,   -14,   -10,     8,    -1,    -8,   -13,   -27,     3,    18,     0,     8,    11,   -32,   -40,   -14,   -17,     4,    11,    -4,    -2,     5,     6,    17,   -25,    -6,     1,   -12,    25,   -12,   -22,    -4,    -5,     0,   -17,   -12,     8,    -9,   -16,     2,     8,     5,   -12,   -11,    -4,    20,     6,    10,     8,    -5,    -4,   -24,    17,    -8,    -5,    -9,    21,   -27,   -14,    13,    12,    18,    -2,     0,     6,     1,    12,    26,    48,    15,   -18,    -9,     3,    23,     8,    11,     4,   -22,   -12,   -17,    12,   -13,     3,   -19,   -14,   -18,    12,     3,    12,    26,    23,    13,   -13,   -10,   -27,    -9,     2,     1,     0,   -22,    -2,    14,    -1,     6,     5,   -23,    -1,    -7,     7,   -21,    -4,     1,   -41,   -11,    21,    15,    13,    13,    -1,     7,     1,   -30,   -35,   -18,   -15,   -13,   -18,   -16,   -14,     6,    10,     2,    -2,   -36,    -6,     5,    29,    -2,    -1,     1,    -3,    16,    -5,   -19,   -26,   -27,   -48,   -14,   -11,     0,   -18,   -33,   -20,   -25,   -14,    -2,    -3,    -4,   -10,   -19,    -8,    -8,    12,    17,    45,     6,    -4,    -2,    -7,     2,   -25,   -36,   -12,   -17,   -30,   -35,   -27,     9,    12,   -22,   -33,   -13,    11,     8,    -6,   -13,   -32,   -22,     5,     8,     1,    17,    34,    12,     3,    -6,     3,     7,     8,    -7,   -18,   -40,   -20,   -23,     8,     4,    19,    10,    -1,    10,   -10,    11,    10,     1,    -6,     0,     3,     6,     9,     7,    12,    20,    -2,     2,     3,    11,    18,     7,   -11,     2,    -9,    -5,     5,     7,    12,     0,    21,    25,    22,    34,    -2,   -24,   -43,   -24,   -11,    -7,   -10,     6,    22,    18,     4,    -7,    14,    16,     1,    13,    -1,   -14,    -2,    -8,    12,    -9,    25,    -1,     2,     1,     7,    -5,   -12,   -20,   -11,    -4,     4,    -5,     2,    -3,    19,    29,     3,     1,   -17,    32,    19,    33,    22,    -2,   -13,    -5,    -3,   -15,    -7,    10,     8,    20,    10,    -2,    -6,    -8,     1,    -8,     1,    -3,    29,     5,    26,    46,     3,    -4,    -4,    28,    37,    17,    15,     5,    -3,    -9,    23,    12,    11,    -5,    -4,     8,    14,    11,    -3,   -21,   -11,    -2,    16,    10,    32,    18,    34,    36,    -3,     4,     6,    15,    19,    20,    22,    17,     6,     1,    -2,     0,   -15,     0,     0,    19,    12,    -9,    -6,    -1,   -11,    -1,    -9,    16,    30,     8,    33,    -5,    -1,     7,     4,    -3,    19,    28,    -5,   -10,    -6,    -6,   -10,   -17,   -17,   -38,   -18,     6,     3,    14,    32,    25,    13,   -23,    -2,    20,    22,    21,    29,     1,     0,    -4,    14,     8,    23,     0,   -19,   -22,   -16,   -14,   -19,   -25,   -31,   -40,   -17,     2,    -6,    15,    14,     6,   -14,    -6,    -4,     5,    19,   -13,   -18,     0,    -5,     1,     9,    10,    12,     4,    -3,    -8,    -5,   -19,   -26,   -23,   -36,   -28,   -22,     5,   -33,   -59,   -19,     2,    -3,     3,   -15,   -18,    -5,     9,    -5,    -3,     4,     4,   -13,     9,   -15,   -19,    -5,   -12,    -4,   -38,   -40,   -36,   -34,   -39,   -18,   -16,   -45,   -66,   -34,    10,     4,    10,   -14,    -7,    14,     1,    -2,    -4,    -1,     2,    -3,   -10,   -20,   -28,   -28,   -23,   -27,   -32,   -34,   -18,   -12,   -31,     6,   -10,   -25,   -23,   -50,   -44,   -22,     3,   -16,   -20,    -8,     3,     4,    -1,     1,    -4,    -1,     2,   -15,   -16,   -16,   -18,   -13,   -40,   -20,    -7,   -10,   -17,    -9,   -24,   -23,   -30,   -39,   -42,   -30,   -26,   -26,    -1,    -5,     3,     5,     0,     3,     3,     1,     2,     1,    -4,     0,     0,    -4,    -3,   -17,   -13,    -3,   -14,   -11,   -12,   -11,    -7,    -8,   -11,   -30,   -33,   -11,     0,     1,    -1,     3,    -2),
		     3 => (   -1,    -4,     0,     5,     0,    -3,     3,     4,     5,     0,    -4,    -3,    -2,    -6,     0,     0,     5,     4,     4,     2,    -1,     0,     2,     4,     4,     5,    -2,    -3,     3,     2,     4,     1,     5,    -3,    -4,    -2,    -4,    -3,     1,    -3,    -8,    -2,    -5,    -9,   -13,   -11,     3,     2,     3,     3,     0,     0,     0,    -4,    -4,    -3,    -2,     4,    -5,     4,    -2,     4,    -6,    -6,    -5,   -19,   -20,    -6,   -17,   -22,   -13,   -16,   -28,   -34,   -29,   -16,   -42,   -36,   -40,   -13,    -3,     0,     1,     3,     5,    -3,     3,    -5,    -5,   -12,    -6,   -14,   -15,   -15,   -22,   -16,    -2,    -5,   -19,   -20,     3,    23,    14,   -10,    -5,   -10,   -29,   -38,   -18,    -3,    -2,    -3,     1,     5,    -5,     8,    23,    10,     1,    13,    17,    27,    23,    -2,     1,    10,    19,     4,   -17,    -6,    14,     1,    -5,   -34,   -15,   -64,   -42,    -3,   -11,     2,     2,     1,     2,    -7,     8,   -11,   -14,   -20,     6,   -17,     9,     9,     2,    -2,    -4,     1,     0,     9,    16,     6,     6,    17,     7,    -9,   -15,   -11,   -11,    -1,     4,     4,     3,    -4,   -13,    -5,    -3,     0,    12,     1,     3,    -3,     9,    31,    13,    -1,    -4,     0,     2,    19,   -20,   -11,     4,     0,    -1,   -17,   -21,    -3,     3,     8,     0,   -19,   -10,    25,     2,    -2,     5,    -1,    12,    20,     4,   -11,     6,    13,    19,    -2,    -3,     1,    20,    -5,   -15,   -32,   -19,   -28,   -19,    -5,     4,    -2,     4,    30,    14,     7,   -14,    16,    -4,   -25,    15,     9,    22,     6,     0,   -10,    -5,     7,    -2,     2,    11,    13,    -6,   -50,   -57,   -15,   -23,    -4,    -5,   -13,    37,    31,     7,   -33,   -10,    -4,   -13,    -4,   -21,   -16,   -39,   -47,   -74,   -33,     8,     3,     7,    12,    14,     7,     3,   -36,   -73,   -30,   -33,     2,     1,    -9,    49,    21,   -18,   -36,   -42,   -59,   -50,   -54,   -49,   -88,   -72,   -65,   -27,    -8,     2,    -9,    -6,     4,     4,    17,    11,   -13,   -66,   -18,   -18,    -5,     1,    -7,    -7,   -13,   -27,   -37,   -58,   -41,   -58,   -78,   -54,   -46,   -23,    18,    26,    27,     3,     9,     0,    13,    32,    21,    15,   -37,   -33,   -29,   -12,     0,    -4,    -2,   -19,   -27,     8,   -10,    -8,   -26,   -12,   -25,   -11,     4,    27,    25,    18,    -7,     2,    -9,    14,   -24,    -5,    -3,    -8,   -12,     2,    -4,    -6,    -5,     2,     0,   -25,     5,    31,    19,    -1,   -13,     3,   -11,     7,    22,    12,    18,    -9,    -2,    -1,   -18,   -21,   -31,   -21,    -3,   -10,    -1,   -19,   -20,    -9,    -6,    -7,     6,    -2,    -1,     5,    27,   -10,   -18,    27,     8,    -2,     9,     9,     9,    -2,     2,    -2,    -5,    -3,   -14,   -25,    -6,   -20,   -24,   -28,   -50,   -14,    -8,    -9,    15,    19,    -7,    17,    -6,   -34,   -44,   -27,   -17,     4,     8,     0,    21,    20,    -6,    -6,     3,    -5,     1,    -9,    -3,   -27,    -3,   -20,   -16,    39,     1,    -3,     2,    17,    21,    12,     0,   -54,   -40,   -58,   -34,   -19,     4,    -4,    12,    -7,   -12,     2,     1,     0,    10,     5,    13,   -21,   -12,   -32,   -17,    14,    -4,     0,     7,    25,    -3,   -25,    -8,   -37,   -13,   -42,   -77,   -93,   -38,   -42,   -41,   -23,   -16,    11,    10,    11,     1,    -6,    12,     3,   -17,   -31,   -32,   -14,    -6,    -9,     6,    33,     8,   -19,    14,     5,    23,    -3,   -10,   -32,   -22,   -47,   -45,   -18,     8,    -8,     0,    -6,    10,    17,    12,    -3,   -41,   -58,   -21,   -14,   -12,    -4,    -5,   -22,    38,     6,     6,    11,     4,    11,   -10,    -9,   -21,   -17,    10,    -1,    -1,    -5,    -6,    -1,    -1,    -5,   -11,   -19,   -26,   -43,   -18,   -15,    -9,    -4,     3,   -40,    29,    25,     2,    -1,     0,    15,     2,    11,     9,     9,     9,    -8,   -15,    -1,     1,    -8,    -8,    -2,   -18,   -30,   -39,   -35,   -10,    -9,    -2,   -10,     5,    -5,    14,    30,    -2,   -12,     8,    23,     1,    16,     7,     3,   -14,   -10,   -18,   -21,     6,    -4,   -25,   -12,   -11,   -21,   -42,   -32,   -12,     0,     3,    -2,    -8,    -3,    12,     9,    14,   -10,   -17,    -4,   -13,    -1,    -3,   -15,   -10,   -14,    -8,    -4,    12,   -23,    -4,   -24,   -28,   -41,   -39,   -32,   -14,    -3,    -3,    -5,     3,    22,    20,     3,    27,   -17,     5,   -12,    -4,    -9,     5,    -6,     0,     9,    -2,    30,    -2,     0,    27,   -14,   -32,   -54,   -41,   -18,   -28,    -2,     0,    -1,     0,    -4,     9,   -11,   -12,     3,   -10,   -10,     6,    -8,   -12,   -12,   -25,    -7,   -17,   -15,   -25,   -10,   -31,   -33,   -28,   -33,   -13,   -17,    -3,     2,     0,    -1,     1,     2,   -20,    -8,    -3,   -15,   -25,   -16,    -3,     7,   -24,    -2,    -5,   -13,   -37,   -37,   -34,   -13,    -8,     0,   -12,   -30,   -19,     2,    -7,     3,     1,    -3,    -4,    -1,   -15,    -5,     4,   -14,   -25,   -37,   -41,   -15,   -25,     9,    25,    16,     2,   -17,   -20,   -13,   -15,   -26,   -16,   -21,    -3,     4,    -3,     2,    -4,     3,     3,     3,     1,    -2,    -1,    -6,     1,     1,   -11,    -2,    -8,     1,    -6,   -15,    -2,   -16,   -13,     2,    -3,   -11,    -3,    -4,    -3,    -1,     3,    -3,    -1),
		     4 => (    2,    -2,     1,     1,    -3,     4,     3,    -3,    -2,    -2,    -4,     0,    -7,    -8,    -9,    -3,    -3,    -4,    -1,     4,     2,     0,     2,     0,    -5,    -3,    -3,    -1,     4,    -1,     1,    -5,    -1,     1,   -14,   -18,    -6,    -8,   -17,    -7,   -19,   -33,   -15,   -15,   -17,   -13,    -5,     2,   -12,    -7,   -11,   -14,     2,     1,     4,    -2,     3,     1,    -3,     4,   -18,    -5,   -19,   -22,   -32,   -14,   -15,   -35,   -21,   -22,   -13,   -13,   -30,   -25,   -23,    -6,   -30,   -27,   -24,   -20,    -6,   -17,     5,    -3,    -3,     1,    -2,   -14,   -36,   -18,   -26,   -15,   -16,   -22,   -12,   -22,   -24,   -21,   -20,   -22,   -36,   -43,   -21,    -5,     2,    -3,    -9,    -6,   -20,   -13,    -4,    -2,    -3,    -3,    -9,   -33,    -5,     5,    25,     7,   -11,   -31,   -21,   -10,    -9,   -29,   -49,   -38,   -22,   -35,   -19,    39,    18,     5,    24,   -14,   -17,    -9,   -15,    -4,    -3,    -2,   -17,   -12,    -3,     5,    22,    -8,    -5,   -10,   -10,    -9,    -7,   -42,   -49,     6,   -20,     7,   -16,     6,     3,     4,     5,   -28,   -12,    -8,    -8,    -4,     3,    -1,    -2,    -4,   -12,   -11,    23,   -20,     9,    16,     4,   -17,   -33,   -69,   -64,   -36,    -9,     6,    24,     0,    -1,     5,   -22,   -29,   -32,    -8,    -1,   -12,     3,   -19,    -4,     3,    -6,    -9,    11,    -2,     5,     6,     9,     9,   -31,   -55,   -77,   -31,   -13,    36,    24,    26,    10,    -4,   -19,   -28,   -27,    -1,    -7,   -28,   -18,   -43,     3,    -4,    10,    10,    14,    -4,     9,    24,    -4,    -8,     3,   -60,   -54,   -23,    33,    23,    14,    -8,   -20,    10,    -3,   -11,   -16,     3,   -26,   -38,    -3,   -28,     5,     5,    27,    12,   -33,    -6,    18,     3,    13,    15,    22,   -30,   -42,    -2,    48,     8,     5,     0,   -24,    -9,   -10,     3,   -29,     6,   -24,   -19,     4,   -15,     0,    12,     9,    -4,   -58,   -14,     8,    20,    -4,    10,    20,   -31,   -34,    22,    22,     3,    17,    13,   -15,   -30,   -19,   -37,   -38,     8,    -2,   -12,     1,   -22,     8,     4,    14,     4,   -21,    -4,     8,     6,    13,    14,     3,   -46,   -47,     4,    12,    -1,     7,   -11,   -28,   -29,   -14,   -27,   -11,     8,    -9,   -29,     3,   -13,    10,    14,    14,    15,     4,     4,   -20,   -12,    11,     0,     4,   -13,   -31,    14,     2,     3,    -1,     5,   -19,     0,    20,    43,    42,    34,   -32,   -23,     0,   -11,   -19,     0,    23,     8,    -7,    -1,    -6,    11,    21,    -1,    -3,    -4,   -11,   -14,     8,    -2,    14,     1,     5,    21,    40,    20,     6,    -3,   -31,     1,    -4,    -3,   -20,     2,    11,    32,     5,    20,    10,    -4,    -2,    -6,   -10,    -5,   -22,     2,    -9,     6,     8,    20,     3,    28,    23,    -5,    12,   -11,   -18,    -2,     4,     5,     5,    -5,    25,    -3,    -3,    21,     0,     3,     0,     7,     3,    18,    13,    18,    14,     6,     8,    20,    -1,    -5,     9,   -17,   -24,   -25,    10,    -4,    -5,    -3,   -28,    15,    26,   -13,   -16,    22,     1,    -8,     4,     2,    -3,     7,    19,    16,    -2,   -11,    13,     0,    -3,     9,   -19,   -26,    -4,    -8,   -11,     1,     0,    -4,    26,    19,    39,     0,   -25,     5,   -16,     3,   -23,   -16,    -8,   -11,     5,   -17,   -22,   -21,    -3,   -37,   -13,     6,   -11,   -15,     1,    -6,     3,     3,   -19,    -3,    19,    22,    28,   -20,   -23,   -25,   -14,    -5,   -15,   -21,   -13,   -10,   -12,   -36,   -26,   -12,   -24,   -26,   -10,     3,     4,    -7,   -10,   -14,     4,    -1,    -2,     0,    -7,    10,    -3,   -31,    -5,   -34,   -18,    -6,    -4,    -3,   -20,    -1,     5,    -4,   -24,     9,   -18,    -6,    -9,    26,     8,     2,   -12,   -19,    -5,     0,     0,     0,    -6,   -21,   -46,   -30,   -27,    -6,   -22,   -27,   -17,    20,     7,    -3,     5,    -3,    -4,    -5,    15,     1,   -12,    -8,    -1,    -4,    -3,   -41,    -6,    -5,   -14,   -13,    -8,   -27,   -18,   -29,   -22,   -21,    -8,   -23,    -9,     3,     4,    -7,    12,   -22,     6,   -16,    -9,   -14,   -21,   -32,    -8,     9,     2,   -34,   -19,    -3,    -6,   -12,    -5,   -13,    -6,     0,     2,   -25,     5,   -35,   -25,     1,     4,   -12,    -4,   -13,    -2,   -11,    -7,   -22,   -19,   -28,     5,    15,    -2,     4,     8,    -3,    -4,    -5,    -7,   -14,     0,   -10,    15,    15,     3,   -43,    -5,   -14,   -14,   -13,   -10,   -15,     1,     1,    20,   -20,   -25,    -5,   -11,     7,   -12,     9,     2,    -3,    -3,     5,    -2,     3,   -35,    -9,   -14,   -10,    -2,    -8,   -20,    -9,   -18,   -13,    30,    -5,    19,    18,    25,   -23,    -3,     4,    -3,    -2,   -30,     1,    -9,    -3,     2,    -3,    -2,    -4,    -3,   -21,   -57,   -33,   -24,   -16,   -24,   -22,   -22,     4,     9,   -19,    -2,     9,     2,   -12,    -4,    13,   -15,     7,   -14,    -6,    -7,     5,    -4,    -2,     4,    -7,    -9,    -4,   -15,   -26,     6,    -5,   -30,   -51,   -44,   -34,   -15,   -26,   -45,   -11,   -28,   -35,   -45,   -42,   -35,    -8,   -13,    -1,     4,    -3,     5,     0,    -2,    -2,    -3,     2,   -15,   -13,   -18,   -19,   -16,   -33,   -18,   -14,   -38,   -11,   -17,   -22,   -17,   -24,   -29,   -25,   -20,    -6,    -3,    -1,     1,     4),
		     5 => (    3,    -1,    -2,     3,     4,     0,     1,     2,    -3,     4,     3,     0,    -1,     1,     0,     4,    -3,    -4,     2,     4,    -5,    -1,     2,    -1,     3,     5,     3,     4,     5,     2,     4,    -3,     3,    -5,     1,     1,     3,     5,     3,    -3,   -10,   -10,   -10,    -9,    -6,   -10,    -3,    -3,    -6,    -1,    -1,     0,    -4,     3,    -4,     5,     4,    -3,    -1,    -5,    -5,    -3,     2,     3,    -6,    -2,   -17,   -35,   -32,   -44,   -15,    17,    15,    19,    28,    23,    29,    22,    21,    24,   -11,    -6,     1,    -5,     4,     4,    -3,     8,    19,    -4,   -12,    -9,    -7,   -25,   -29,   -22,    -9,   -22,    18,    -8,   -33,   -26,    -3,    -6,     9,    14,   -10,    -4,    13,    11,    15,     5,     2,    -7,   -10,     2,   -25,   -25,   -32,   -37,   -52,   -17,   -40,   -27,   -26,     0,    27,     2,    10,    -1,     0,    -3,     5,    14,    20,    22,    27,    54,    14,    -4,    -1,    -4,    -5,    -4,   -23,   -22,   -46,   -45,   -54,   -28,    -4,    -2,     9,     1,     3,    -7,     8,    20,    12,     3,    39,    33,    18,    32,    35,    51,    24,    -8,     2,    -1,    10,    -8,   -24,   -41,   -42,   -26,   -13,   -24,    -6,     4,    25,     2,     0,     2,    11,    18,    38,     5,    31,     0,     3,    31,    11,    25,    17,     4,    -2,     5,    -4,   -14,   -20,   -27,   -12,    -3,    -8,     2,     0,    23,    15,     5,    -9,   -13,     4,    14,    17,     1,    17,    -1,   -18,    -3,   -11,    10,    12,     8,    -5,    -6,   -15,   -12,   -16,   -10,   -25,   -12,   -19,   -27,     9,    28,    15,   -20,   -18,   -31,   -61,   -33,   -31,   -81,   -38,   -44,   -31,   -12,    -7,    -4,     9,     2,     0,    -8,   -30,   -34,   -31,    -4,   -29,   -34,   -29,   -15,   -14,    -8,   -10,   -18,   -33,   -76,   -96,  -110,  -119,  -115,   -81,   -62,   -56,   -31,   -19,   -16,     1,     5,     2,    -6,    -2,   -18,    -3,    -9,   -18,   -12,    -2,   -12,   -15,     3,   -15,     3,   -24,    -7,     2,   -23,   -69,   -71,   -69,   -57,   -54,   -37,   -21,     0,     3,     3,    -3,    -1,    -2,   -11,    -4,   -12,   -21,   -21,   -16,   -19,   -15,    -9,    -9,     0,   -11,   -10,     9,     3,    10,   -11,   -34,   -58,   -42,   -19,   -22,    -4,     7,    -9,     3,    -3,     0,   -11,    -3,    -9,    -9,   -17,   -10,   -17,    -8,     8,     7,     6,     7,     3,     5,   -11,   -10,     1,   -11,   -20,   -30,   -22,    -8,    -7,     0,   -14,    -2,     0,    -4,    -5,    -2,     9,   -13,     3,   -21,     8,    16,    29,    12,    -6,    11,     3,    -2,    -6,   -15,     5,     2,    11,   -12,    -8,   -17,     1,    -2,    -8,     9,    -5,    -3,     3,    17,   -17,   -28,   -24,    -5,    -8,    18,     2,     1,   -10,     4,   -19,    16,     3,     3,   -18,     0,     3,     0,     1,    -7,    -5,    -9,    -8,    -1,   -14,    -9,    -7,    15,   -17,   -28,   -21,   -24,   -13,   -13,    -7,    10,   -12,   -23,    -6,   -18,    10,    -7,    -5,   -13,     4,    -2,     6,     5,    -4,    -5,    -2,     0,     3,   -13,     4,     0,   -25,   -26,   -40,   -41,   -65,   -52,   -32,     6,     4,   -17,     7,     6,    33,    -7,    11,     7,     9,    12,   -16,   -21,   -13,   -14,   -14,    -3,   -10,   -27,     6,   -13,   -16,   -19,   -40,   -19,   -51,   -69,   -23,   -28,   -37,   -29,     8,    -9,   -14,    29,    15,    18,    11,    -8,   -12,   -30,   -15,    -6,    -9,    -1,    -7,     2,    14,     1,   -13,   -21,    -6,    16,   -10,    -3,   -19,   -51,   -27,    -2,   -12,     7,     0,    20,   -10,    -2,     8,    -2,   -10,   -29,     4,   -25,   -19,     1,    -1,    21,    -2,     3,   -17,    -4,    -7,    11,    17,     5,    16,    11,     7,    10,    -5,    10,    -4,     8,     7,     7,   -10,     1,   -17,   -26,     2,    -7,   -10,    -3,    -2,    14,     7,    49,    -2,     6,    -2,    26,    18,     2,     7,   -19,    21,    19,     8,     2,    -1,    -9,    15,    11,   -13,    16,   -29,   -19,   -13,    -4,     2,     2,    -6,   -13,    -7,    31,    26,     1,    -5,     6,     1,     9,    17,     8,    11,    -4,     8,    10,   -11,   -17,    11,    17,    20,    18,     2,   -10,   -15,    -1,    -4,     3,     2,   -19,     4,   -14,    -9,   -14,    -8,   -11,    -8,    26,     5,    12,   -11,    -2,   -10,     2,    -5,     8,     3,    24,   -10,    -9,   -12,   -17,   -15,    -1,     1,     1,    -4,     9,    12,   -15,   -14,     6,     3,    27,    14,     4,   -23,    -9,    -9,    -1,    28,    -4,   -28,   -24,   -20,   -24,   -19,     3,     9,   -39,   -41,     5,    -1,    -5,    -1,   -17,    -2,    22,    19,    55,    27,    -5,    16,    33,     0,     9,     6,    20,   -17,   -27,   -13,   -21,   -24,    -5,    14,    18,    -3,     1,   -12,   -14,     4,    -4,    -1,    -2,    21,   -10,    -2,    19,    26,     7,    22,    18,    15,     8,     3,   -13,    -6,   -11,   -27,     6,    13,     3,     6,    14,     3,    -3,     2,    -2,    -3,    -3,     3,     5,     0,   -10,   -12,    -6,    -2,     1,    -5,    11,    10,     9,    -8,   -10,    -6,    -4,    -6,    -7,    -3,     4,     3,     9,    -4,     2,     2,     3,     0,     0,    -2,     3,    -4,    -2,     0,    -5,     3,    -1,    -4,     5,    -2,     1,     4,    -6,     2,    -5,    -5,    -7,    -9,    -7,    -7,    -7,     5,     2,     0,     3,    -4),
		     6 => (   -3,    -2,     3,     3,     3,    -4,    -3,    -3,     2,     3,     2,     3,    12,     6,    -1,     1,     1,    -1,    -3,     1,    -1,     2,    -3,    -2,     2,    -2,     3,    -2,     4,     4,    -4,    -4,     3,     1,     8,    10,    18,    25,    22,     9,    23,    16,    -8,     1,    10,    20,     1,    16,    19,    16,    14,    19,     5,     3,    -3,     3,     4,     2,     7,    15,    22,    13,    15,    17,     4,    -3,   -13,    18,    29,    13,    13,    36,    20,     9,    12,    -5,    -6,    -2,     3,    -1,     7,     8,    -2,    -4,     3,    -2,    -1,    44,    24,    -6,    21,    30,    -6,     5,   -13,     8,     8,    20,     9,    -9,    -8,     1,   -17,    -2,    14,    -1,    -3,    -7,    -6,     1,     4,    -5,     0,     3,   -15,    21,    -2,    11,    12,    -9,     2,     1,     9,    13,   -16,    -3,    -4,   -21,   -13,   -13,   -17,    27,    22,    10,   -12,   -26,   -14,   -15,    -3,     9,    -3,     2,     4,    -8,    -1,   -30,   -23,    -9,   -16,    18,     1,   -14,    11,    16,    -7,   -10,   -24,     6,     8,    14,     6,    -1,   -14,   -22,   -16,    -7,     5,    10,    -4,    -5,     6,   -22,   -20,   -38,   -31,    -5,   -15,     0,   -24,    18,    25,     4,    -3,    -8,    -7,   -19,     8,    -2,   -22,    -2,   -26,   -34,    -7,    -9,    14,    -4,    -1,    -5,     2,   -21,   -18,   -48,   -31,   -15,    -7,    -7,     5,    28,    20,     2,    12,   -16,   -20,   -18,   -48,   -38,   -38,   -22,   -33,   -41,   -24,   -17,    10,   -24,     2,    -1,     5,   -22,   -16,   -52,    -7,    -9,   -23,    13,     6,    -5,    21,     4,   -17,   -35,   -33,   -56,   -51,   -49,   -33,   -37,   -62,   -48,   -40,   -28,    -9,   -22,     4,    -3,    -9,   -13,   -12,   -55,    -2,     4,    -4,   -17,   -14,     2,   -10,   -23,   -21,   -42,   -40,   -57,   -57,   -50,   -30,   -55,   -51,   -36,   -10,   -10,   -13,    -8,    -4,     2,    -7,   -15,   -26,   -50,   -30,     2,    12,     0,   -15,    -2,    11,   -17,   -50,   -46,   -11,    14,    -2,   -24,   -17,   -13,   -24,   -10,    -8,    15,   -18,   -21,     3,     0,     3,   -30,   -22,    -8,   -21,     0,    17,   -12,    -3,     5,    11,   -40,   -36,   -10,    12,    16,    13,   -15,     0,   -34,   -17,   -23,   -22,    -4,   -30,   -16,     3,    -5,     5,   -17,   -21,   -23,   -12,    19,    12,    -4,   -15,     1,   -14,   -54,   -16,    -3,    21,     8,    -1,    15,    17,    -3,   -12,   -16,    23,    -7,   -18,   -17,     2,     1,   -12,    -9,   -35,   -29,     0,    25,    12,   -31,   -23,     1,   -10,   -23,   -18,     2,    -5,    -5,    -2,    20,    31,    14,    -6,     8,     5,    -8,   -18,    13,     1,     2,    -3,   -23,   -41,   -15,    21,    14,     6,    -8,     9,    24,    -6,    -6,    11,    -5,     9,   -15,    14,    13,     7,    16,    21,     7,    -5,     2,   -12,    -4,     2,    -1,    -6,   -20,   -30,     1,    30,    17,    -5,     0,    -6,    32,     4,   -15,    21,    -8,     1,    -9,    12,     3,     3,    12,    25,    11,     0,     8,   -25,   -32,    -5,    -5,    -6,   -17,   -11,    18,    36,    -5,    -6,   -28,    15,    26,    -5,   -17,    26,    -5,    -6,     0,    -5,    -5,     9,    22,    15,     2,     6,     0,   -31,   -27,     5,     0,     1,   -11,    -1,   -11,    16,     9,   -15,   -16,    -1,    11,     5,    -5,     4,    -3,    -7,   -16,     8,   -11,   -16,    19,    22,     2,    27,    24,   -12,   -26,     3,     0,     5,   -18,     0,    -9,     7,    16,     0,   -22,     3,    -3,    20,     7,    14,   -21,    -8,   -19,    -6,    10,    -6,    24,     9,    19,    16,    32,   -16,   -27,    -4,    -1,    -3,   -18,    14,   -28,   -21,     9,    -3,   -13,   -17,     3,    14,    13,    20,    17,     2,     1,   -14,     7,   -15,    -9,   -21,    17,     7,    22,    -8,    -2,     3,    -6,     0,   -19,     9,   -12,   -20,     0,   -29,   -12,    -8,     0,   -11,     2,    28,    30,     7,     2,    21,    -6,    -7,    -8,     9,    16,    21,    27,    -1,     3,    -2,     1,     0,    -2,     2,    -8,     4,    -2,   -24,   -29,    -5,   -20,   -32,   -24,    19,    20,    -7,     8,    -3,     5,    14,   -15,    15,    27,    10,     5,    10,     2,     4,     3,    -4,    -8,    -8,   -11,    13,   -33,   -58,   -58,    -4,   -15,   -17,   -17,   -21,   -12,   -31,   -20,    11,   -21,   -21,   -21,     7,   -10,   -47,   -31,    10,    -4,    -4,    -3,    -5,    -1,   -16,     0,   -15,   -19,   -24,   -11,    29,     8,   -44,   -35,   -40,   -43,   -43,   -53,   -49,   -11,   -13,   -31,   -26,   -38,   -43,   -14,   -14,     1,     3,     2,    -3,    -3,    -5,    -6,    -7,    -2,    -8,    -9,   -16,     0,   -11,   -25,   -39,   -28,   -17,   -26,   -29,   -48,   -21,   -22,   -10,   -14,   -23,   -16,     1,    -1,     0,    -2,     4,    -3,    -1,     3,    -6,    -8,     2,    -9,    -4,     8,    12,     3,    -1,    -2,     0,    -8,    -1,   -14,   -22,   -16,   -15,   -24,    -2,    -3,     1,     0,    -3,     2,    -3,     2,    -1,    -3,    -2,    -5,    -3,     0,     2,    -6,    -2,    -6,     0,     1,     2,     0,    -2,    -3,    -7,    -5,    -4,     2,     4,     2,    -2,     0,     1,    -1,     1,     4,    -3,    -1,    -5,    -3,     2,     0,     2,    -2,    -1,     4,    -1,     3,     3,    -2,    -2,     3,    -3,     1,    -6,     3,     1,    -2,     3,    -1),
		     7 => (    1,     1,    -3,    -1,     5,    -4,    -4,     5,     1,     4,     1,     2,    -2,    -3,     1,    -2,    -3,     2,    -2,     3,     2,    -1,     4,     4,     0,    -4,    -2,     3,    -1,     2,    -2,     0,     1,    -5,     1,     1,    -2,     4,    -6,   -11,    -4,   -10,   -12,   -12,   -21,   -22,   -14,    -4,    -2,     6,     7,    -3,     5,     1,    -4,     2,     0,    -4,     3,    -2,    -3,    -4,     1,    -8,   -12,    -4,   -23,   -42,   -20,   -12,    -9,    -6,   -11,    -6,     0,    -2,   -10,    -2,    -4,     8,     2,    -5,     2,    -1,     4,     1,     1,    -5,    -1,   -16,   -24,   -19,   -24,    -3,    -5,   -16,   -28,   -36,   -18,   -16,   -16,    -8,     0,   -11,    -7,    -5,   -13,    -8,    -2,     1,     5,    -4,     3,    -2,    -4,    -2,    -9,   -10,   -10,   -31,   -40,   -20,   -41,   -11,     5,    -3,   -21,   -32,   -38,   -42,   -28,   -22,   -16,   -13,   -27,   -38,   -26,   -23,   -15,     0,     1,    -2,    -1,   -31,    -9,    22,    33,    19,    30,     9,   -15,     6,     6,     9,    18,    10,     4,    -6,   -23,   -30,   -49,   -33,   -29,   -45,   -67,   -46,   -13,     5,    -4,     3,    -6,   -22,    -3,    15,    16,    16,     7,    -2,    16,     0,    24,    10,    11,   -12,   -18,   -12,   -23,     0,     1,   -10,   -26,   -25,   -51,   -27,   -28,    -9,    -2,    13,     0,     7,     7,    15,     7,    -1,    -2,   -16,     4,   -15,    11,    -6,   -17,   -28,   -14,   -17,   -25,   -23,    -5,   -21,     6,     8,    -9,   -30,   -32,   -12,   -15,    28,    14,     2,    25,    33,     0,    16,     4,    10,     5,   -18,   -12,    -9,   -12,    10,     7,     6,    -3,    -4,     2,     1,    -3,   -13,     1,   -43,   -40,   -15,     0,    21,     5,    15,    23,    31,     9,     6,    35,    10,   -17,   -22,   -17,    -2,    -4,     6,   -12,     0,    12,    -5,    11,    11,    13,   -10,   -14,    -1,    30,    41,     3,    -3,     3,   -10,    11,    -4,    16,    21,    18,    -1,    -2,     4,   -12,    -3,   -10,    -6,    -5,    13,    20,     9,    15,    11,     7,    -5,     0,    20,    13,    36,     0,   -12,     7,    21,    -2,    -9,    26,    38,    24,    19,     2,     0,     1,     4,     5,    -4,   -12,    23,   -12,    23,    12,    -9,   -15,   -18,    -9,   -29,    -8,    27,     0,     5,     5,   -14,   -23,   -40,    -2,    -2,     4,     1,   -16,   -13,   -12,   -29,   -17,    -4,   -11,   -20,     2,     0,    -1,    -4,   -13,    -9,    -6,     5,    21,    33,    -4,     8,    20,   -25,   -27,   -31,   -11,   -10,   -23,   -29,   -34,   -31,   -48,   -52,    -7,    -5,    -1,    -7,    20,     8,    13,    -8,     6,    29,    12,    12,   -23,   -20,    -8,    -7,    -7,   -22,   -20,   -33,   -23,   -33,   -54,   -42,   -38,   -38,   -45,   -25,     4,     3,    10,    -3,    12,    20,    26,   -13,     4,    -5,   -15,   -37,   -26,    -6,    -1,     0,   -12,    -3,   -36,   -17,   -15,   -45,   -24,   -17,    -2,    -5,     7,    -1,    14,    17,    -9,     9,     6,    -7,    27,     4,    14,    -6,    -9,   -45,   -18,    -8,    -4,    -8,    -9,    -7,   -25,   -22,   -23,   -30,     2,    18,    18,    17,    19,    12,    12,   -17,   -14,    -1,    -5,     6,    -1,     8,    14,   -15,   -51,   -50,   -21,   -13,    -3,    -4,    -2,   -17,   -16,   -20,   -28,   -35,    -1,     5,   -21,    -1,     1,     9,    10,   -16,   -12,   -23,     8,    12,     5,    -7,     9,   -12,   -20,     4,    -5,   -10,     6,    -6,    24,   -12,   -24,   -39,   -43,   -28,   -17,   -46,   -30,    -5,    24,    26,   -24,   -24,   -18,    -7,    -5,   -20,   -15,   -23,   -12,   -21,   -19,   -10,    16,    -8,    -3,     9,     4,    -7,   -19,   -49,   -26,   -28,   -23,     7,   -15,   -13,    -1,    -6,   -16,   -13,    -5,   -24,   -15,   -10,   -12,   -21,   -17,   -23,   -39,    -5,   -20,     0,     4,    -6,     1,    -9,   -27,    -5,     3,    13,   -10,    -6,    -5,    -4,     6,     7,   -22,   -27,   -21,   -34,   -34,   -26,    -9,     2,     9,    -1,   -17,    -8,   -32,    -3,    -6,    -5,    -2,   -28,   -20,    21,    25,   -13,     8,     0,    -7,   -15,    -8,     8,   -48,   -32,   -44,   -47,   -28,   -31,   -25,    -4,    -6,   -23,   -19,    -5,    -8,    -7,   -11,    -9,    -7,   -43,    14,    23,    21,    26,    32,     9,     9,     1,   -11,   -19,   -31,   -30,   -32,   -26,   -36,   -26,   -28,     3,     8,   -47,   -27,    -3,   -10,     1,     0,     4,   -12,   -50,    12,    -3,    16,    42,     3,     1,    -7,    11,   -16,   -11,   -30,   -14,   -34,   -57,   -44,   -41,   -39,    -3,     1,   -21,   -16,    -2,   -23,     1,    -5,     0,    10,    -3,    20,    31,    21,     7,    26,     4,   -10,     8,    -8,    10,   -18,   -14,   -49,   -50,   -41,   -26,   -35,     3,   -10,   -37,    -5,   -14,    -4,     4,    -4,    -1,    -8,    19,   -20,     4,    -1,     9,   -11,   -22,    -4,    13,    -5,   -27,   -35,   -27,   -32,   -18,   -12,   -17,   -44,    -4,    -7,   -29,     5,     1,    -6,    -4,     5,     3,    -2,   -22,   -26,   -28,    -7,    14,    24,     9,   -13,    -1,     8,    15,   -17,    -6,    -1,   -10,     5,    -2,   -13,    13,    19,     9,    -7,     1,     4,    -4,     0,    -2,     0,     4,    21,    19,    -4,    -2,    -5,     0,    13,     9,    -9,    29,    19,     2,     7,     4,     4,    -4,     6,    23,    17,    21,    -1,     3,     1,     1),
		     8 => (   -2,     2,     1,     2,    -2,     3,    -3,     0,     4,    -3,    -1,     4,    -1,    -1,    -1,    -3,    -4,    -3,    -2,    -2,    -5,    -3,    -3,    -3,     0,     0,    -2,     3,     3,    -3,    -3,     3,     1,     4,     4,    -4,     3,     5,     1,     1,    -1,    -6,    -4,    -5,   -14,   -12,    -6,     3,    -3,     0,     3,     2,     0,     4,     4,    -2,     2,    -4,    -4,     4,    -5,     4,    -2,    -1,    -5,   -14,   -36,   -31,    -9,    -8,    -5,   -15,   -20,    15,    24,     8,   -15,   -15,   -14,   -15,    -5,    -7,     4,    -1,    -1,    -5,   -11,   -10,    -8,   -14,    -9,   -28,    20,    15,    -9,   -23,   -21,   -16,   -15,     6,     4,     4,    32,    16,     0,   -11,    21,    28,    -1,    -7,   -10,     5,     1,    -3,   -10,   -15,   -27,   -36,     0,    15,    -4,   -22,   -19,    11,    -6,    -1,     6,     7,     9,     3,    -5,     1,   -11,     0,    12,   -13,   -22,    17,    19,    -1,    -2,    -3,    -7,   -16,   -16,   -27,     1,    -2,   -27,   -15,    -9,     0,    -3,    11,    -2,     8,   -10,   -27,   -34,    20,    -4,    20,     2,    -9,    -9,    -3,    -9,    -7,     3,     0,   -16,   -28,   -20,     4,    -4,   -13,   -22,   -10,     5,   -11,    -9,    -9,   -24,     0,   -14,   -14,   -15,     9,     1,    -8,    -8,   -21,   -19,   -13,    -3,    -2,     3,   -22,    -6,   -10,    -2,    -3,   -10,   -11,    -2,    -4,   -17,    -4,   -12,   -27,   -16,     7,    -5,   -19,   -14,     3,     1,    -5,   -20,   -17,   -17,    -1,     6,    14,    -9,   -16,    -5,    -3,   -11,    -2,   -19,    -8,     3,     9,   -24,   -19,   -12,    -3,   -10,   -10,   -16,   -22,   -12,     3,     4,     8,   -26,   -30,    -9,     2,    30,    15,    -2,    -6,   -16,     2,    -8,    -8,   -16,     7,    -1,   -10,   -25,    -3,    -8,   -15,   -23,   -21,   -11,   -12,   -24,    11,     5,   -26,   -29,   -25,   -20,    -1,    10,   -15,     4,    -7,   -14,     0,    -7,     5,   -14,   -14,    -4,     1,    11,    31,   -10,   -13,     7,     3,     3,     3,     8,    13,     1,   -10,   -20,   -31,   -14,   -18,     4,     6,     0,    -6,    -7,   -15,   -11,    13,     8,     0,     8,    19,    11,     3,   -12,   -21,    -9,    -6,    10,    -5,     2,   -18,   -20,    20,   -13,   -13,    -6,   -40,    -2,   -20,    -3,     1,   -14,    -1,    15,    20,    13,    -4,     5,    17,    13,   -19,   -11,   -21,   -17,   -22,   -12,    -9,    -1,   -21,    -3,    11,    12,    18,     6,   -34,   -36,   -27,     5,    -2,   -19,   -29,     4,    11,    -7,   -26,    13,    40,    15,    12,    -4,   -13,   -18,    -2,     2,   -31,    -9,     1,    10,    24,    18,    18,    -3,   -31,   -47,     6,     0,     1,    -1,   -35,   -17,    -5,   -10,   -29,     6,     4,    -4,     1,     5,    -2,   -12,   -12,   -43,   -19,    14,    21,    21,    17,    -9,   -27,   -38,   -29,   -45,     0,    -5,     2,    -8,     9,     4,   -18,   -15,   -13,     2,    -3,    11,    17,    -2,    -2,   -16,   -35,   -13,    -7,   -14,     5,    -6,   -24,   -28,   -15,   -11,     0,   -23,   -18,     2,    -2,    -4,    18,    -3,   -15,   -18,   -16,   -40,   -27,    -8,    10,    13,   -14,   -10,    -9,    -1,    -4,    -2,   -15,    -4,     6,   -14,    -4,     3,    -5,   -26,   -14,     2,    -3,    -9,    13,   -12,   -17,   -22,   -12,   -35,   -63,   -24,     6,    19,    -3,    -3,     3,     4,   -11,   -26,   -24,     4,   -11,   -12,   -11,   -10,    -5,     3,    -8,    -5,     2,   -11,   -13,    -7,   -14,   -18,   -19,   -12,   -21,    -1,    -2,    10,     7,   -11,    13,    10,    -8,    -7,    -8,     2,   -15,    -8,   -16,    -6,    -3,    -4,   -12,     3,    -2,    -9,    -7,    -4,   -12,   -25,   -30,     9,    10,    -1,    -7,    12,     8,    -6,    17,   -15,    -4,     0,     1,   -17,   -15,   -12,   -10,     0,    -1,   -15,   -17,     4,    -3,    -7,     0,   -11,    -9,   -29,   -32,    -7,     8,    -6,    -6,    -5,    10,   -14,     3,   -22,   -23,    -8,    -2,   -30,   -12,    -3,     1,     0,     0,   -11,    -1,    -9,    -4,   -10,    -1,   -13,   -16,   -23,    -5,   -18,   -17,   -10,     8,    26,     8,    10,     4,   -12,   -11,    -8,   -10,   -17,   -14,    -8,    -8,   -12,    -6,   -15,    -5,    -8,   -12,    -5,    -7,   -10,   -32,   -36,   -20,   -13,   -12,   -29,   -14,    15,    11,    12,   -19,    -2,     1,    -1,     1,    -8,     0,    -1,    -1,    -7,    -5,   -14,    -1,    -3,     1,   -12,    -3,    -4,   -17,   -31,   -40,   -13,    -2,   -15,    -1,   -14,    -6,   -20,    -9,     4,   -14,   -12,     1,     9,    10,     3,    -6,     1,    -1,   -16,    -1,     5,    -3,    -2,    -4,    -7,   -11,   -11,   -19,   -15,   -14,   -35,   -12,   -15,   -16,    -8,    13,    10,   -10,    17,    10,     1,    -3,    -7,    -8,   -27,   -19,    -7,     4,    -2,     4,    -7,    -2,    -7,   -18,   -12,    -6,   -12,   -13,   -20,   -25,    -4,     7,    -6,    11,    -3,    -3,    11,    10,     4,   -20,    -7,    -8,    -1,    -8,    -3,     2,     1,    -2,    -2,    -7,    -6,   -12,   -19,    -7,    -5,    -9,   -15,   -31,   -37,   -30,   -31,   -45,     1,    -4,    -5,   -38,   -34,   -19,   -13,     5,    -4,    -2,     5,    -3,     1,    -2,    -3,     2,    -7,    -2,    -6,    -3,    -1,    -9,    -2,   -11,     3,   -10,     0,    -1,     0,     2,    -1,    -2,    -1,     2,    -5,    -3,     2,     4,    -2,     3),
		     9 => (   -1,    -3,     3,    -3,    -2,    -5,    -3,     4,     3,     1,    -4,     0,     1,     0,     5,     5,    -2,     0,    -5,     3,    -1,    -3,     3,     2,     5,    -5,    -1,     0,     5,    -2,     4,     3,    -4,     3,    -6,    -2,     4,    -1,    -2,    -3,   -13,    -7,    -2,    -1,    -5,    -5,    -9,     4,     0,    -7,    -3,    -5,    -1,    -1,    -2,    -2,     0,     1,     3,    -3,     2,     4,    -1,    -1,    -3,    -5,    -7,    -1,    -1,    -2,   -14,    -2,    -6,    -2,    -5,    -1,   -13,     6,    -5,    -6,    -5,     5,     0,    -3,     0,     0,     3,    -8,    -1,    -8,    -6,    -1,   -16,    -7,   -10,   -22,   -14,    -5,   -12,   -12,   -14,    -6,    12,    -7,   -12,   -17,   -13,     1,    -7,    -6,     1,    -2,     0,    -4,     0,    -8,    -7,     2,   -21,    -5,    -6,    -2,    -9,   -11,   -30,   -39,   -44,   -43,   -23,    -3,    15,   -21,   -32,   -23,   -16,   -14,   -13,   -28,   -20,     2,     0,     3,    -4,    -6,     1,    -5,    -9,   -11,   -29,   -16,   -25,    -7,    -8,     9,   -11,   -17,   -35,   -37,   -36,   -31,     4,   -16,   -21,   -24,   -15,   -13,   -31,     2,    -5,    -6,     0,    -7,     8,   -13,    -5,   -31,   -24,   -23,   -31,   -12,   -14,   -23,    -8,    -9,    -9,   -23,     1,   -16,     7,    14,     0,   -10,   -14,   -17,   -21,   -20,    -2,    -7,   -12,   -11,   -16,   -27,   -29,   -35,   -40,   -55,   -45,   -35,   -17,   -14,   -18,   -34,    11,     7,    -3,    -4,    42,    16,    16,    11,    -7,   -20,    -8,   -13,   -16,    -6,     4,     0,   -19,   -15,   -19,   -26,   -30,   -43,   -14,   -28,   -12,    -6,   -27,   -10,     3,    16,    16,     2,     3,    -3,    -2,    17,     7,   -13,   -19,    -9,    -4,    -9,    24,    -2,   -11,   -17,   -10,    -4,   -33,    -6,    -7,   -11,   -14,   -26,     5,    21,     4,     1,    -5,    14,   -17,     3,     8,    -1,    14,    13,   -40,   -19,     0,    -6,   -16,   -14,    -2,   -12,   -22,   -28,   -11,    -1,    -4,     9,   -12,     8,    -5,   -19,   -19,   -16,   -36,   -33,   -16,    -7,   -13,    -4,    23,    48,   -17,   -29,     5,   -40,    -9,    -6,   -11,   -18,   -17,    -5,    23,    12,    16,    -6,     5,    -8,   -21,   -36,   -40,   -46,   -21,    -8,    12,    -5,    11,     5,    34,    45,    -3,   -25,     2,    -4,     4,   -24,    10,   -12,   -21,    -2,    10,     6,    18,    -9,   -27,   -19,   -34,   -24,   -10,   -35,     0,    -1,    22,    -6,    14,    18,    -7,   -34,   -29,   -29,    -4,    -7,   -10,   -17,    11,   -15,    -2,     7,     4,    11,    26,     2,     2,     5,   -15,    13,    25,     2,    -1,    27,     9,    29,     5,   -10,   -23,   -15,   -16,     2,     0,    -7,     2,   -16,    13,   -14,    -1,   -11,    25,    26,    23,     0,    11,    12,    10,    16,     3,     4,    -1,    12,    -8,   -29,   -11,   -36,   -32,    -7,     4,     1,    -3,     3,   -29,   -19,    14,   -15,   -21,   -17,     5,   -13,     4,    12,    13,    28,     1,     8,    -3,     1,    16,     7,   -23,   -28,   -39,   -30,   -24,    -5,    26,    -5,    -5,    -7,   -19,   -17,     9,   -10,    -3,    -1,   -14,    -7,     6,     9,    -9,     5,   -19,   -22,     1,    11,     5,    -3,   -34,   -12,   -11,   -36,   -18,    -2,    -4,    -2,     2,    -5,   -16,    -5,   -13,   -15,   -10,    14,   -14,   -24,   -17,   -13,    -9,    -5,   -12,    -6,    -1,    18,    13,   -14,   -17,    -8,   -18,   -36,   -15,    20,    -2,    -7,     0,     3,   -17,    -7,   -33,   -24,     0,    13,   -16,   -26,    -6,     7,   -10,    -6,    11,   -13,    -3,    -8,     8,     2,   -15,   -12,    -3,   -13,    -8,    23,   -13,   -13,    -1,    -4,   -19,   -12,   -35,   -30,   -13,   -11,   -22,   -33,   -21,   -27,    -3,   -14,    -3,   -17,   -19,   -13,    -5,     1,   -33,   -15,    -2,    -6,     7,    27,   -18,   -13,     3,     0,    12,   -10,   -26,   -15,   -45,   -34,    10,   -13,   -30,    -5,    17,    12,    -6,   -20,    -6,    -2,     1,    -7,   -19,   -17,   -13,    -3,     7,    24,    -5,    -4,    -1,    -4,    -4,   -13,   -27,   -13,   -31,   -23,     8,    11,     2,   -12,    -6,   -15,   -12,   -37,     2,    -9,    -8,     7,   -18,   -14,   -19,    -8,     5,    19,   -20,    -2,     4,     3,   -16,   -26,   -31,   -26,   -41,   -13,     8,    13,    15,    10,    -5,   -17,   -27,   -20,   -12,    -8,   -29,     1,     4,   -17,    -9,     1,     8,    -2,   -11,    -4,     0,     3,   -14,   -18,   -40,   -20,   -25,     4,    22,    16,     5,   -17,    -5,   -25,   -25,    -7,     2,    -4,    -6,    -5,     5,    -1,     3,   -16,    -5,     8,   -10,     4,     3,     4,    -8,   -14,   -18,     0,     2,    12,     5,    16,     6,    -6,     0,   -25,     5,   -18,   -16,    -1,   -14,     9,     2,    -1,     8,     0,    -3,    -2,    -7,    -1,    -5,     4,    16,    -7,     7,    -3,    -8,    -2,    10,     5,    16,    -2,    14,    -1,   -15,   -14,     5,    20,    13,     3,    -7,   -10,   -13,    11,     3,    -2,    -2,     2,     4,     5,     0,    27,    13,    -5,    15,    13,   -10,     1,     8,    24,     4,    19,    15,     9,    28,    35,    18,    13,    26,     4,   -11,     8,    -6,     1,     2,    -4,    -3,     3,     4,    -2,    -8,    -5,     7,    27,    24,    17,    16,    34,    18,    15,    12,    13,     6,    12,    19,    26,    -9,   -12,    -6,    -7,     5,    -1,    -5,    -2),
		    10 => (    3,     4,     2,    -5,     2,    -2,    -4,     1,     4,    -3,     2,    -1,    -4,     1,     0,     1,     1,    -2,    -4,    -2,     1,    -2,     0,     2,    -4,     0,     0,     3,    -1,    -5,    -3,    -4,     3,     5,    -2,     2,     4,    -6,    -5,     5,    12,     1,    -8,    16,    21,    23,     0,     3,     3,     0,     0,    -2,    -1,     0,    -3,     3,     4,     5,    -6,    19,    17,    -5,    -4,     4,    -7,    -8,   -15,    -2,     0,   -11,    -5,   -23,    -3,   -28,   -23,   -25,   -20,    -7,   -23,   -14,   -11,    -3,    -5,     5,     4,     2,     3,    -1,    -5,     0,    -6,    -2,     9,   -15,   -39,   -23,     2,     5,    -3,   -19,   -16,   -32,    -4,    -1,     2,   -18,   -19,   -11,    -2,     4,   -35,     0,     4,     4,    -5,    -7,     5,   -25,   -17,   -21,   -14,   -26,   -28,   -22,   -40,   -42,    -9,     8,   -20,     6,    -9,     0,    -3,     1,     8,     6,   -18,   -27,   -29,    -3,    -3,    -5,   -11,    -4,     4,   -30,   -15,   -30,    -9,     0,   -35,   -14,   -26,   -17,    -2,    -5,   -13,    -1,   -12,    -3,   -35,   -16,    17,     2,   -28,   -18,   -24,   -18,     1,     2,   -20,    -3,    -6,    -3,   -13,   -12,     4,    -4,   -11,     2,   -10,     2,     1,   -11,    -8,     0,     5,     2,   -16,    12,    22,   -13,   -28,   -28,    -2,    -4,     0,   -24,   -13,    -8,    -5,     2,    -4,   -20,    -3,   -10,    -3,     4,    -4,   -10,    -8,     4,   -13,     3,    14,     5,   -28,    -1,    -9,   -12,   -40,   -29,   -20,    11,    43,   -34,    17,     8,    -6,    -7,    -7,   -23,   -12,   -11,     0,    -2,     7,   -39,     6,    17,     0,    23,    16,   -20,   -28,    -6,   -12,   -13,   -40,   -16,   -30,    -5,     3,    -7,    26,    -3,    -5,     6,   -16,     5,     9,    -9,     4,    -3,     1,     0,   -11,   -13,    17,     9,    14,    -7,    15,    -8,   -18,   -18,   -17,   -37,   -32,     0,    -1,     2,    15,     8,    -4,    -2,    -5,    -8,    -7,    -3,     6,    -2,    -1,    -8,     4,   -33,   -12,    12,    -2,    -1,    -8,   -17,     2,    -5,   -24,   -22,   -26,    -2,    -3,    51,   -17,   -17,   -19,     4,     8,   -16,   -33,   -28,    -4,     3,    -7,     8,   -21,   -37,   -29,    -5,     9,    13,    -2,   -30,   -31,   -23,   -31,   -30,   -18,     2,     1,     7,    -8,   -22,    19,    21,     5,   -13,   -46,    -5,     8,     3,    17,    -2,   -29,   -39,   -16,     3,    17,    22,     7,   -24,   -29,   -12,   -24,   -31,   -11,    -4,    -3,    12,    14,   -18,    37,    18,    11,     3,   -17,    15,     8,    -5,     2,   -20,   -48,   -65,   -25,     2,     5,    24,    33,   -21,   -11,    13,     3,    -2,   -19,    -8,     3,     3,    -5,   -25,     2,    21,   -17,     5,    12,    12,     6,    27,    22,    -5,   -35,   -27,   -22,   -16,    13,    33,    29,   -22,     0,    19,    -2,   -12,   -11,    -6,     4,    -3,   -17,   -30,   -20,   -12,   -12,    -4,    10,     4,    13,    24,    49,   -19,   -49,   -25,    -9,    -2,    26,    -6,    12,   -27,    -2,    12,    -7,    -7,   -40,    -7,     4,     2,   -14,   -18,   -13,    -5,   -20,   -21,    15,    -4,    -8,    12,    15,   -35,   -51,    -5,     8,    10,    11,     9,   -21,   -35,   -24,    -7,   -16,   -23,   -34,    32,     3,    -8,   -16,   -22,    -5,   -15,   -27,    -9,     6,    -7,     1,     0,     7,   -29,   -28,    -3,    10,     8,    -9,     8,    -3,   -34,   -13,   -15,   -16,   -20,   -20,    50,    -1,    -7,   -18,   -18,   -17,   -35,   -22,   -12,     1,    -6,     8,     4,   -20,   -25,   -17,     2,    26,     8,     5,   -11,   -16,   -21,     0,   -17,    -9,   -15,   -24,   -12,     1,    15,     0,   -14,   -19,   -21,   -30,   -12,    19,     3,    -1,     4,    -4,     5,   -11,    -9,   -24,   -13,    16,    -8,    -9,     2,   -15,   -17,    -2,   -27,   -15,    -6,    -5,    18,    -7,   -16,    -5,   -20,   -35,   -15,     7,     3,    13,    15,    18,    11,    -3,   -31,   -23,    -5,   -16,     2,    -9,     7,   -18,    -6,   -21,     2,    12,     4,     4,     1,    -9,   -21,   -25,   -12,   -22,   -15,     1,     5,    26,     3,    24,    10,   -16,   -15,   -13,   -13,     3,    12,     1,   -11,   -19,    -3,     0,     6,    62,    14,     3,    -5,   -20,   -33,   -27,   -15,   -25,   -19,   -10,    17,    -1,    -1,     1,   -26,     6,    12,    13,   -15,   -28,    -5,   -26,   -21,   -15,    -9,    -3,    10,    34,    14,    -5,     3,    -2,   -22,   -26,   -42,   -18,   -14,   -16,    18,    34,    11,     6,    -6,    -3,   -17,     3,   -10,     0,    -5,   -26,   -21,    -6,    -7,     0,     1,   -28,     1,    -3,    -1,    -8,     0,    13,     9,   -27,   -35,   -38,   -28,   -25,   -15,    -4,   -18,   -24,   -15,   -17,    -7,    12,   -32,   -20,   -17,   -12,    -4,     4,     6,     3,     3,     5,    -1,    -6,     0,   -19,   -16,   -18,   -28,    -8,   -14,   -36,   -42,   -70,   -68,   -70,   -54,   -32,   -26,   -26,   -25,   -32,   -25,   -14,   -12,     1,    -1,    -2,     2,     5,    -4,     2,     4,   -13,   -18,   -45,   -13,   -18,   -35,   -23,   -26,   -18,   -19,    -7,   -25,   -24,   -25,   -33,   -29,   -26,   -21,   -10,   -11,     1,     2,     2,     2,    -1,    -4,    -4,     4,    -2,     3,    -4,    -8,   -10,     1,    -2,    -2,     0,    -5,    -6,    -7,    -4,     0,    -4,    -1,     2,    -5,    -1,    -5,     2,    -3,    -3,     1),
		    11 => (    1,     1,    -4,    -5,     4,    -4,     5,     3,    -1,     2,     5,    -5,    -3,    -4,     4,    -4,     1,     3,    -3,    -1,     1,    -4,     2,    -4,     4,    -1,     4,    -4,     1,    -1,    -4,     5,     0,    -4,     1,     2,     5,     0,     0,    -5,    -3,    -9,     0,    -7,   -10,    -8,    -1,    -4,     1,    -4,    -3,     3,    -3,     4,    -2,    -4,    -4,    -5,    -4,    -4,    -4,     1,     3,     1,    -8,    -4,     7,     5,     1,    -3,    -5,   -16,   -37,   -45,   -36,     9,    12,   -15,    -7,   -12,    -4,    -4,     1,     1,     3,    -5,    13,     2,    -3,    -4,    -5,    17,    15,    20,    16,     4,     3,     0,     4,   -23,   -37,   -28,    -4,   -13,   -12,   -20,     5,    15,   -15,     0,    -1,     4,    -2,     4,    12,    10,     5,    10,    14,    13,    -5,     1,   -14,   -11,   -10,   -14,   -15,   -29,   -22,   -11,     4,     9,    20,     0,     0,    -8,   -23,   -18,   -26,   -21,    -1,    -2,     1,    22,    17,    17,    -4,     1,   -26,   -14,   -22,   -24,   -10,    -8,   -44,   -48,   -31,     3,     9,     5,    -1,    19,    16,     7,     4,   -16,   -19,    -2,    -1,     0,    -3,    20,    34,    -6,   -13,    -3,   -29,    18,    14,    -2,   -44,   -50,   -64,   -52,   -25,   -16,     0,    -5,    -6,     4,     0,     4,   -13,   -21,   -15,   -10,     2,    -7,   -12,     1,   -15,   -17,   -13,   -16,   -33,     0,    21,     2,   -28,   -40,   -44,   -35,   -12,    -7,    13,     0,     2,    -3,    -3,     6,   -28,   -42,   -25,    -7,     0,   -18,   -14,    -4,    -7,   -10,   -10,   -20,   -20,    -7,     2,   -27,   -22,   -25,   -44,   -21,    -1,     9,     6,    -1,     9,    -6,    -1,    -3,   -28,   -34,   -26,    -8,    -3,     1,   -13,    -5,    -7,   -11,    -9,   -10,   -10,    -2,   -37,   -41,   -43,   -70,   -62,     0,    16,     3,     7,    -4,    -5,    -7,     2,    -1,    -7,   -21,    -8,   -15,    -3,     2,    -6,    -2,     0,     0,   -23,   -24,   -33,   -20,   -36,   -36,   -48,   -59,   -29,    -2,    27,     4,    -9,    -3,    -1,     8,     6,    -2,     5,   -10,   -12,    -9,    -4,     2,     6,     3,    -7,     4,   -10,   -27,   -30,   -24,   -31,   -19,   -28,   -21,   -14,    32,    12,    11,    33,    -7,    -1,     3,   -18,   -27,   -17,     2,   -15,     2,    -2,     1,   -14,     8,    -1,    10,     3,   -22,     2,   -36,   -23,   -25,    -9,   -15,     9,    24,     1,    12,     4,     8,   -24,    -2,   -20,    -4,   -14,     2,    -7,     0,    -4,     1,   -11,     0,     1,   -12,    -6,   -12,    -9,   -20,    -9,    -5,   -16,     4,    24,    15,     4,    15,    10,   -10,   -55,   -24,   -24,    -8,   -10,    -5,    -1,     1,    -3,    -2,    -2,     0,     6,    -8,    -6,     0,    -3,    15,    18,    -7,    -1,    17,     6,     8,    14,   -22,   -30,   -64,   -70,    -9,    10,    -1,    -5,   -12,    -7,    -3,     1,    -5,    13,    24,    -2,   -26,    -1,     4,    35,    14,    11,     2,    -5,     5,     4,    12,     4,   -20,   -58,   -71,   -42,    -6,     7,     1,   -46,   -34,   -22,     0,     3,     0,     5,    -7,     7,    -6,   -15,     1,    14,    13,   -21,    -2,    -7,    -1,   -17,    11,    11,    -5,   -41,   -39,    -5,    11,    13,    27,    38,   -15,   -23,    -7,     0,     0,    -1,   -13,     0,   -29,   -13,     7,    -1,     1,    -6,    16,    14,    -2,     3,   -19,     5,    -2,     7,    15,    19,    34,    42,    39,    30,    -2,   -43,   -16,     1,    -1,    -3,    -1,   -18,   -48,   -30,     4,     3,    -2,    -6,    14,    -6,    -3,     2,    -6,   -14,    -2,     7,    11,    11,    -2,    24,    19,     0,     8,    -3,    12,    -2,     4,     4,   -17,   -29,    -9,     2,     8,     6,    -3,    -9,    -4,    -3,   -19,   -38,   -29,   -19,   -28,   -22,   -14,   -12,    -7,    14,    19,    19,    20,    -1,     6,    -2,    -2,     0,   -14,     7,    15,    13,     3,     6,     1,   -11,    12,   -14,   -27,   -28,   -19,    10,   -13,   -29,   -18,   -19,    -7,    16,    15,    28,     0,     4,     8,    11,    12,     2,     0,    -4,     0,    -2,     5,     4,    -8,    -8,    -3,   -10,    -5,    -9,     6,    15,    11,   -16,   -14,   -20,    -9,     5,    28,    23,    11,     3,     4,    15,    12,     1,     1,     6,    26,     8,    -1,     7,    15,    -9,   -14,   -22,    -2,   -19,    17,    20,     0,   -17,   -22,   -20,   -20,     3,     4,     5,     1,     5,     2,     1,     0,    -7,    13,     2,     2,     2,     1,    22,    12,    -7,   -19,     4,     8,    10,    17,     6,   -11,   -14,   -17,    -8,    -2,    -3,    -4,    13,    25,    30,     2,    -1,     2,     3,     8,   -23,   -17,   -23,   -31,    -6,    19,    -4,   -14,    18,    28,     3,     3,    -2,     1,     0,    -8,    -1,     4,     5,     3,   -15,     4,     1,     3,    -1,    -2,     4,   -11,   -20,   -20,    -6,   -41,   -10,     8,    -8,     7,    21,     6,   -30,   -19,   -15,   -27,   -16,   -10,    -5,   -15,   -11,   -10,   -11,    -3,     0,    -3,    -1,    -4,    -1,    -3,   -19,   -14,   -15,   -22,   -28,   -23,   -16,    -8,   -15,   -15,   -12,   -13,   -18,   -20,    -8,     1,    -3,    -3,    -2,    -3,     2,    -1,    -4,    -4,     3,     0,    -5,     3,    -2,    -3,     1,     2,     2,    -3,   -16,    -7,    -4,    -2,    -9,    -5,     4,     2,    -5,     0,     0,     0,     4,    -3,    -2,    -2,    -4,     4),
		    12 => (    5,    -4,     5,    -3,     1,    -1,    -1,     5,     1,     3,    -4,     3,     3,    -4,     9,     5,    -5,    -3,     2,    -2,     1,     2,    -3,    -3,     1,     1,     3,    -3,    -5,    -4,    -3,    -3,     0,     0,     1,    -7,   -16,    -6,    -7,    -9,    -8,   -13,    -4,     4,     5,    -2,    -5,   -16,   -10,    -9,    -1,     5,    -1,     2,    -5,    -2,     4,    -2,    -6,   -15,   -10,     4,    -1,    -5,     1,     4,     6,    16,     5,    -8,    -6,   -15,   -17,   -10,     5,     6,     3,     3,   -14,    -5,    -8,     3,     3,     3,     0,     5,    -6,   -29,     1,   -15,    -7,   -14,    -2,    15,    29,    21,    16,     4,     1,     2,    -1,    -1,    -8,     0,     3,     5,   -14,   -25,   -13,   -12,    -4,     2,     0,    -1,    -2,   -11,     3,     8,    18,    25,     2,    -1,     7,    22,    21,    25,     0,    -4,    -1,   -11,    -3,   -17,    -9,   -14,   -16,   -15,   -27,   -22,   -22,    -5,     5,     4,   -17,    -2,     1,    10,    18,    34,    16,     8,     7,     2,     6,     6,   -11,    -8,   -12,    -9,   -11,    -5,     2,     5,    -7,   -13,   -23,   -10,   -12,    -5,    -5,    -3,     0,     0,    -3,     1,    24,    20,    13,    12,     4,     1,    -6,    -1,    -8,   -11,    -8,    -7,    -3,   -14,    -2,     6,     4,   -15,     0,    22,   -11,     1,     3,    -4,    -2,    -2,    -6,     5,     1,     7,    -1,   -13,    -9,     0,    -7,   -10,    -6,     5,     6,   -16,   -14,   -18,     2,    10,    -6,   -16,     7,    26,   -34,   -14,   -15,    10,    -6,     1,    -4,     1,    -6,     3,   -17,   -21,   -10,   -12,    -3,     2,    -1,     3,     4,    -5,   -12,    -6,    -4,    -1,    -5,     6,     4,    -3,   -32,   -16,     3,   -14,    17,     0,    -7,    -6,   -11,    -9,   -14,   -19,   -10,   -12,    -2,    -5,    18,     3,   -12,    -4,   -10,    -8,    -3,     6,     6,    -1,    -9,   -18,     0,   -12,     3,    -2,     5,    -4,   -16,    -6,   -12,   -21,   -30,   -26,   -29,   -11,    -3,    -9,    -8,     1,   -18,    -5,   -20,    -5,   -17,     6,    10,   -10,   -19,    -8,     9,   -18,    -2,   -10,    -6,   -17,   -13,   -10,     1,   -28,   -30,   -30,   -27,    -9,    -2,     3,     8,    -7,   -20,   -13,     6,    -3,    -9,    -8,    -5,    -8,   -14,    -7,    -1,    -8,    -2,    -7,   -18,   -19,    -8,    -4,   -13,   -16,    -7,    -8,    -7,     4,    14,    -1,    -3,    -5,   -11,    -6,   -11,     1,   -18,   -20,    -8,   -17,   -21,     1,     8,     4,     3,    -6,   -10,   -13,   -14,   -21,    -7,   -18,   -12,    -5,     0,    -4,    -1,    -3,    -4,    -6,   -13,   -11,     5,     0,    -7,    -7,   -15,   -17,    -5,     6,    17,     1,    -1,   -12,    -9,    -5,   -15,   -23,    -4,   -15,   -11,   -12,   -11,   -18,   -17,   -11,    -9,   -14,   -18,   -19,     1,    -5,    -4,   -22,   -16,   -15,    -5,    13,    21,    13,     1,   -15,   -10,     1,   -12,     2,   -12,    -8,    -1,   -13,    -7,   -10,   -14,    -2,    -5,   -15,   -28,   -20,    -1,    -1,     2,    -9,   -15,   -18,     8,    20,    26,    19,     2,    -7,    -3,    15,    13,    -1,    -7,   -10,    -6,    -5,     5,     2,     5,     5,     3,   -10,   -15,   -14,   -17,   -11,    -8,    -6,   -12,   -15,     2,    16,    31,    21,    -4,    -4,     5,    16,    13,    -4,    -2,   -18,    -8,    -5,    -9,    -9,    14,     3,    -9,    -9,   -19,   -18,   -11,   -18,   -21,   -13,   -13,   -23,     0,    25,    20,    24,     4,     0,    -5,     4,    16,     0,   -17,    -7,     0,     3,    -2,   -13,    -1,    -4,    -1,    -3,   -21,    -9,   -17,   -15,    -7,    -8,     2,    -1,    15,    14,    16,    19,     1,    -2,    -1,     7,     4,    -8,    -3,    -7,    -3,    -8,     3,     6,     1,     2,   -12,    -9,    -2,    -6,    11,   -25,   -10,     7,    12,    18,    18,    20,    34,    37,     2,    -7,     4,    -2,     7,     7,    -5,    -6,    -9,    -1,     2,    12,    -1,    -7,   -10,   -13,    -6,    -9,    10,   -16,    -3,     9,    15,    21,    23,    12,    11,    -4,     2,     2,     8,    11,    -6,     4,    -2,   -11,   -15,   -12,   -11,    -4,   -11,    -8,   -13,    -8,    -2,     3,    -5,   -10,     5,    12,    22,    21,    11,    -3,     4,    -7,     0,     3,     2,     6,    11,    -7,    -4,    -9,    -4,    -8,   -15,    -8,    -5,    -5,     7,    -9,     8,    -7,   -12,     0,     2,     9,    20,    19,     5,    15,   -16,    -8,    -1,     2,     2,     5,     4,     0,    -3,     0,     7,   -10,    -5,    10,     1,     4,     6,     5,     1,   -15,   -19,   -14,     3,     8,    21,    25,     1,    12,    -8,     3,    -2,     5,   -10,    -5,   -10,   -11,   -11,    -2,    -6,    -4,   -14,     1,    10,     1,    12,    -1,   -15,   -10,   -10,    -1,   -12,    -5,   -13,     9,     7,     4,     1,    -1,    -3,     2,   -18,    -5,    -2,    -3,     1,    -3,   -12,   -16,   -18,    -6,   -15,   -28,   -11,   -13,   -19,    -3,   -13,    -1,   -13,   -12,   -14,   -10,    -7,    -3,     1,     4,     0,     4,     1,     2,    -9,   -16,   -11,   -12,   -15,   -22,   -20,    -9,    -7,   -13,   -26,   -19,   -40,   -43,   -37,   -30,   -16,   -12,   -20,   -14,     1,    -1,     5,    -5,     3,     2,     2,    -1,     0,     3,    -6,    -7,   -11,    -6,   -12,   -14,    -7,   -22,   -14,   -13,   -15,   -13,   -17,    -6,   -11,    -7,   -11,     4,     1,    -2,    -5,     5),
		    13 => (   -2,    -5,     4,    -2,    -4,     1,    -5,    -4,     4,     2,     4,    -3,    -5,    -5,    -1,     0,     3,     5,    -1,     2,     5,     2,    -2,    -5,     3,    -1,    -2,     2,     2,     1,    -3,     4,     1,    -2,    -4,    -1,     4,     0,    -3,     2,     0,    -3,    -7,    -4,    -9,    -3,     4,    -2,    -4,     0,    -3,     2,    -2,    -3,     5,     1,     2,     2,     0,    -2,     4,    -2,     3,     0,   -11,   -22,    17,    11,    20,    -7,    -8,   -10,    -5,     1,    -3,    -2,   -11,    -7,   -16,    -9,     0,     0,     2,     4,     0,     3,    -2,     2,     1,    -8,     4,    -6,   -13,   -20,   -24,   -15,   -19,   -49,   -71,   -55,   -44,    -6,     6,    -1,   -18,   -16,   -13,   -22,    -2,    -3,     0,    -4,     5,    13,     1,     7,   -18,   -22,   -14,   -10,    21,   -13,    12,    22,   -18,   -11,     1,    -6,   -19,    16,     5,   -18,    -8,    14,    -9,   -10,   -18,    -9,    -7,     0,     3,    -1,    19,     0,    26,    31,    17,    14,   -13,   -19,     0,     0,    -3,    -7,     4,     0,   -11,    -8,    -6,    -4,   -27,   -26,   -12,   -22,    -9,   -22,   -11,    -4,    -1,    -1,     5,     8,    21,    24,     8,     1,    -9,     0,    -2,    17,     0,    15,     8,     5,    -2,    11,     1,   -47,    -3,   -16,   -33,   -18,    -7,    -9,    -2,    -5,    -4,     4,     9,   -12,    30,   -11,    27,     8,     3,    14,     3,    10,     2,     9,     9,   -23,   -12,     0,     4,   -12,    -8,     0,   -31,   -21,   -13,   -12,   -15,    -5,    -2,    -4,     7,   -13,    28,     6,     4,     9,     0,    33,    18,    10,    -8,    -3,   -12,     0,    -2,     8,    13,   -10,   -21,     2,   -18,   -47,   -29,    -9,   -20,     4,     4,   -14,    18,     8,    21,     2,    31,    36,    17,    16,    -1,   -29,   -21,    -4,     4,    12,    -1,     3,     2,    11,     4,    -7,   -35,   -35,   -39,   -14,   -11,     0,     4,   -17,    20,    30,    26,    15,    18,    10,   -31,   -45,   -61,   -31,   -25,     6,     9,    20,    -5,    29,    -2,     3,     5,   -10,   -26,    -1,   -21,   -14,   -13,     1,     4,   -10,     2,    29,    11,   -15,   -30,   -49,   -77,   -41,    -9,   -10,    13,    27,     2,    -3,   -16,   -13,     5,    -2,     8,    -2,   -35,   -25,   -14,   -12,    -4,    -1,    -3,    -2,    24,    27,   -18,   -39,   -63,   -38,   -39,     3,    22,    14,    20,    16,     4,   -14,   -24,   -19,   -19,   -39,   -24,   -50,   -25,   -39,   -17,    -1,     1,    -7,    -4,     2,    -7,    -9,    -6,   -25,   -39,   -31,   -16,     2,    20,     6,    11,     6,     6,   -19,    -8,   -14,   -22,   -21,   -30,   -33,   -13,    -9,    -8,   -17,   -13,    -7,    -5,     9,     2,    12,     0,   -19,   -22,   -14,    24,    -1,     6,    -3,     4,    -2,    15,    -8,    -8,   -10,   -27,     7,   -19,   -17,   -20,     8,    -2,   -38,   -18,   -10,    -8,     9,     8,    20,   -12,   -17,    -9,    -6,    -4,    12,    19,    37,     1,     4,     6,    10,    -1,   -21,   -22,     0,     2,    18,   -22,    25,    -3,   -19,    -8,   -12,     5,     3,    10,    19,   -22,   -30,   -18,   -12,     8,    25,     1,     1,    19,    18,    14,    -6,     1,    -4,    -1,   -14,     5,    29,    12,    14,    -5,   -28,   -28,   -12,     3,     6,    10,    20,   -23,   -43,   -42,   -36,   -16,    -9,   -26,    -4,     5,    13,     2,     2,    13,     3,    -4,     4,   -10,    22,    24,     2,   -13,   -43,   -20,    -8,    -7,    -1,    17,    35,    -8,   -25,   -35,   -45,   -72,   -96,   -79,   -83,   -80,   -60,   -40,   -53,   -14,    32,     3,    10,    11,     8,    37,    20,   -15,   -34,   -17,   -14,     0,    -6,   -29,    19,    16,    18,   -15,   -18,   -30,   -42,   -64,   -70,   -64,   -55,   -44,   -49,   -26,   -11,     5,    22,    21,    15,    24,    27,    -5,   -22,   -29,   -15,     2,     5,   -20,   -11,    -5,    18,     7,    -5,    -2,   -22,   -22,   -19,   -16,    -4,    -6,   -26,   -30,    -5,    -1,    15,    14,    -5,     3,    50,    -3,   -22,     1,     2,    -3,     3,    13,    15,    11,    -2,    15,     9,    -2,    -6,     3,    -1,    10,    13,    -9,    -5,   -13,    -2,     9,     5,    23,   -13,   -14,    -4,   -17,   -20,    -6,     3,     4,    -3,    21,    19,    27,    16,     8,    13,    23,     9,    -3,   -10,    -1,    13,   -16,     2,    -3,   -15,     6,     3,    10,     8,    -1,     9,   -33,   -24,     0,    -4,    -1,     2,    21,    28,    25,    -2,     1,    10,     9,     6,    -5,    11,   -10,     9,    -9,    -7,   -10,   -10,   -26,     0,   -19,    -8,   -20,    -1,   -22,    -4,     4,     4,     5,     5,     7,    -3,    31,    20,     8,    29,    20,     0,    21,    16,     9,    -3,     6,   -10,   -12,     4,    -6,   -19,   -32,     2,    13,     3,   -21,     1,    -1,     0,     4,     1,    -5,   -17,     6,    23,     6,    12,    19,    11,    -4,   -11,   -17,   -22,   -27,   -17,    -6,   -31,   -31,   -31,   -22,   -18,   -11,   -55,   -24,    -5,    -4,     1,     4,     0,     4,   -12,     2,     1,   -16,    -7,   -23,   -26,   -30,   -31,   -26,    10,    -9,   -20,    22,    -1,     6,    -4,    -3,     2,   -15,    -2,    -1,    -4,     3,     0,     5,    -5,    -1,    -3,    -6,     3,    -3,     4,    -1,   -25,   -18,   -13,     1,   -16,   -10,   -12,    -6,    -1,    -8,   -18,   -21,    -4,    -9,    -3,    -1,    -4,    -4,     2),
		    14 => (    0,    -5,     4,    -4,     3,     3,     3,    -5,     0,    -3,     0,     0,   -14,    -9,     0,    -1,     1,    -4,    -2,    -4,     3,     0,    -3,     5,     5,     3,     3,     3,     2,    -2,     4,     3,     2,     0,    -1,    -9,    -4,    -7,   -15,   -14,   -19,   -13,    -5,   -42,   -35,   -27,    -8,    -6,   -15,    -8,    -4,    -4,    -3,    -1,     0,     3,     4,    -5,    -2,   -15,   -42,     1,    -3,   -14,   -23,   -17,   -34,   -33,   -34,    -1,     8,     8,   -33,   -22,   -11,   -11,   -31,   -16,     3,    -2,    -3,   -21,    -1,    -4,    -1,     0,     1,   -15,   -42,   -33,   -14,    -6,    -7,   -13,   -30,   -33,   -22,     1,    12,     1,   -25,   -31,     0,    15,    22,    18,    -8,   -21,   -33,   -18,     2,     0,     3,    -2,    -6,   -29,   -13,   -16,    -9,     7,    13,    19,    -2,   -32,   -33,     2,     3,    -5,    -9,    -9,    12,    -3,    18,     4,    -3,   -17,   -32,   -20,   -24,    -4,     0,     3,   -12,    -5,   -11,     0,    12,     8,    21,    11,    -3,   -27,   -28,   -18,    -1,   -12,   -21,     5,     6,    14,    -2,    -3,     1,    -1,   -10,    12,   -27,    -7,    -3,     0,   -20,    -8,    13,    14,     4,     6,     1,   -12,     2,   -11,    12,    10,    24,    48,    48,    36,    23,    20,     4,    23,   -12,    -3,    -7,   -14,     2,   -11,    -1,   -36,    -9,     6,     7,    10,    22,    22,     1,     8,     9,    -3,    12,    14,    12,    31,    36,    29,     3,    -6,     1,    -1,     2,     2,   -10,     6,    -5,   -37,   -17,   -42,    -4,     3,     1,     3,    26,    17,    21,    -4,   -19,    -3,   -11,    -2,    -8,     5,     1,    -9,     0,     1,    -4,     3,    -4,    -2,     6,    13,    -3,   -31,    -2,   -19,   -22,     2,     0,     5,    -1,    -3,    -4,   -32,   -32,    -6,   -18,   -28,   -33,   -15,   -12,   -13,    -1,   -14,     1,    14,     4,     5,   -11,    -6,   -12,   -23,     2,   -15,     3,    -1,   -11,    -7,   -15,   -11,   -17,   -19,   -13,   -12,   -16,   -41,   -45,   -29,   -25,   -16,     3,    -7,   -18,    17,    -7,   -32,   -38,   -24,   -14,    -7,    -1,   -14,   -12,     0,   -18,     1,   -15,    -8,   -19,   -19,   -15,   -19,     1,   -16,   -37,    -3,   -14,     6,     6,     9,    -7,     9,   -16,   -47,   -44,   -30,   -19,   -30,    -3,     2,     3,     8,    -9,     7,    12,    -2,    10,    11,    12,     4,    17,    13,   -22,    10,     8,    -2,    -2,     8,    12,    36,     9,   -10,   -27,   -17,   -35,   -38,    -3,    -6,   -16,    -1,    19,    -4,     0,    -3,    13,     8,     1,    17,    10,    -6,     7,    28,    14,    16,    17,    20,    14,     9,    -7,    -7,   -28,   -12,   -26,    -1,    -3,    -7,   -42,    -8,    19,    -6,    -5,    -2,    -5,     0,   -14,    -6,   -19,    -7,     4,    27,     7,    18,    27,    18,    20,     6,     1,   -11,     3,   -16,    24,     4,     3,     1,    21,     5,    15,   -25,   -11,     1,    -7,   -18,   -39,   -23,   -14,    13,    22,    37,    34,    29,    29,    -3,     1,     6,     8,    -9,   -21,   -23,    25,   -20,     2,    -1,     3,    13,    14,   -18,   -19,   -10,   -14,   -23,   -31,    -4,     6,    29,    43,    35,    40,    10,    26,   -10,     2,    -4,    -8,   -12,   -10,     3,     3,    -8,     5,    -1,    10,    -9,    30,   -24,   -10,   -11,    -3,   -22,    -5,    11,    30,    29,    25,    29,    40,    12,    19,   -16,    -8,    -3,     3,     2,   -16,     3,    17,   -21,   -27,    -4,    -1,    -4,    25,   -17,   -10,   -13,   -44,   -10,     6,    10,    22,     4,    26,    24,    28,    10,    -2,   -20,     4,     2,    -4,    28,   -24,   -30,    -8,    -3,    -1,    -7,   -17,    19,    -1,    -5,     2,     2,    -3,    10,    13,    34,     0,   -17,    14,    15,    -2,   -13,    15,     6,    -7,     5,    -2,    -2,   -18,   -15,    -9,    -3,     3,     2,    -8,   -17,   -28,   -23,   -18,     3,    21,    16,    20,    20,    17,    18,    -5,     8,    29,     3,    21,    10,    16,     7,     3,    -2,   -24,   -36,   -20,     1,    -4,    -7,   -27,   -13,   -32,    -3,   -36,    -2,    10,     6,     1,   -12,   -26,   -24,    26,    18,    10,     8,    -4,    10,     7,    -7,    12,     5,    -8,   -54,   -31,     2,    -5,    -8,    -5,   -22,   -66,   -31,    -6,    -4,     3,   -32,     2,   -11,   -15,    -7,    -6,    14,    -2,   -21,    -9,     8,    -5,    10,     1,    12,   -16,   -28,   -12,    -9,     1,     0,    -1,   -37,   -56,   -49,    15,    -1,   -21,   -23,   -10,   -16,   -17,    -8,     7,    -8,   -10,    -9,     6,    19,     3,    -9,   -18,    -2,   -12,    -4,    -7,    -3,     4,     0,    -6,    -7,   -40,     7,    -2,   -14,   -27,   -22,   -24,   -14,   -11,     3,    -4,   -14,     1,   -13,     1,    27,   -16,   -23,    -6,     6,   -25,    14,   -18,     2,     1,     5,    -1,    -2,    26,    19,   -24,   -28,   -22,    -1,   -24,     7,    -2,    15,     7,     6,    -3,   -19,   -11,    -7,   -23,   -30,   -10,    12,    -7,   -20,   -20,    -4,    -4,     3,     4,   -19,    28,     2,   -16,   -38,   -22,   -20,   -26,   -16,   -45,   -34,   -39,   -40,   -27,   -39,   -30,   -15,   -42,   -64,   -67,     1,    -2,    -2,    -4,    -1,     2,     1,    -3,     1,    -4,    -7,   -10,   -17,   -20,   -19,   -35,   -27,   -20,   -23,   -40,    -5,   -22,   -29,   -17,   -23,   -27,   -22,   -27,    -2,    -3,    -2,     2,     3),
		    15 => (   -2,    -5,     0,     5,    -3,    -2,     2,    -4,     4,     4,    -1,     0,     2,    -1,    -1,    -2,     5,     5,    -2,    -1,    -5,    -2,     3,     0,     1,    -4,     0,    -2,    -3,     0,    -2,     0,     4,     5,    -5,     3,     5,     1,    -4,    -5,   -11,   -13,   -11,    -8,   -11,   -19,   -11,    -7,    -9,    -4,     2,     1,    -1,    -5,     0,    -4,    -5,    -5,    -3,    -6,    -3,     4,    -6,   -15,   -13,   -27,   -13,    -4,   -12,   -21,   -26,   -34,   -15,    -9,     2,     0,    -6,   -15,    -3,     3,    -8,    -5,    -5,    -2,     1,    -1,   -10,     9,     4,   -11,    -1,   -21,   -22,   -21,   -22,   -11,    -9,   -23,   -23,   -36,   -42,   -23,   -10,    -4,    -4,     7,     7,    -5,   -10,   -12,     3,    -4,    -4,     1,    -6,     6,    -6,    -5,    -3,     8,    -9,     5,   -21,   -17,   -29,   -29,    -6,     7,   -22,    -9,   -12,    -9,   -19,    -4,   -12,     9,    10,   -12,   -22,   -23,     1,    -4,    -7,     0,    -3,     6,    13,    11,   -20,   -19,     5,    -4,   -14,   -26,     3,     8,    -7,   -16,   -15,   -12,     4,    -5,   -22,   -31,   -24,    -6,   -11,   -15,     3,    -6,    -2,   -13,   -10,    12,    10,    -3,   -14,   -16,   -11,     4,    -9,    -2,    17,   -13,   -21,   -28,   -22,    -3,    -3,   -11,    -2,    -5,   -14,    -1,    -1,    17,     3,    -7,    -6,   -19,    -4,     5,     5,   -13,   -16,   -26,     4,     3,    -9,   -18,     7,   -17,   -25,   -25,   -49,   -46,   -40,   -15,    -2,    -7,     7,     6,     7,    13,    -1,   -22,   -21,   -22,   -16,    19,     0,    -7,   -32,    -9,    13,   -16,    -6,     2,   -21,   -41,   -22,   -18,   -40,   -37,   -20,   -17,   -16,    -5,     2,   -17,   -37,    -1,    -1,    -5,    -8,   -19,   -11,    15,   -16,   -30,   -11,    -2,     8,     0,     1,   -33,    -8,   -29,     8,     8,    10,   -11,   -15,    -2,    -9,     4,    24,     7,    -8,    -6,    -3,    -8,    -2,    -4,   -18,    -8,    -2,   -23,    -4,    -3,    11,     2,    -7,    16,    -5,     7,    23,    24,    26,    27,    21,    12,    15,    45,    29,    37,     9,    -7,     2,    -4,    -6,    -6,   -10,   -12,    13,   -12,    -2,     3,     9,    21,     2,    -7,    -6,    -5,    20,     2,    15,    17,    31,    36,    40,    43,    11,    19,     1,     1,    -4,    -1,    -3,   -15,   -26,   -10,    -2,    -9,    -3,    21,    21,     4,     7,     0,    13,     2,    -7,    -4,     1,     7,    36,    19,    30,    22,     5,    19,    41,    -5,    -3,    -3,    -3,    -8,   -32,    -6,   -17,   -15,     8,     6,    17,     4,     3,    -5,   -11,   -34,    -7,    -5,   -50,   -31,   -20,   -27,    -4,   -10,    -4,     2,    36,   -11,     0,    -3,   -11,   -24,    15,    12,    -5,    -2,    21,     8,    10,    25,    10,    14,   -32,   -35,   -28,   -25,   -16,   -35,   -12,   -18,    -9,   -17,   -22,   -24,   -13,     1,     5,     4,    -7,   -14,    35,    -2,     7,    -4,    -7,    14,    -4,     5,    25,    -2,   -24,   -19,   -31,   -31,    -9,   -22,   -15,   -10,   -14,   -23,    -3,   -35,    -7,   -10,    -6,    -9,    -9,    -2,   -30,   -19,   -31,   -12,   -23,   -15,    -7,    -8,     1,     0,    -8,    -4,    -3,    -1,    -4,   -20,   -25,    -7,   -25,    -6,   -13,   -32,   -16,   -12,    -4,    -5,    -8,   -12,   -18,   -25,   -28,   -42,   -35,    -7,   -31,    -1,    -7,   -23,     3,    -2,   -11,    -2,    -1,    -9,    -2,    -8,   -33,    15,   -21,   -37,   -20,   -33,    -3,     1,    -7,     4,    -2,    -4,     0,    -7,   -26,   -14,   -12,    10,     8,   -15,   -23,   -27,    15,     8,     2,   -16,    -4,   -14,   -15,     9,   -14,    -8,   -21,   -17,    -2,    -4,    10,   -21,    -4,   -21,    14,    13,   -16,    -9,    -3,     4,    -8,     0,     9,     4,    19,     4,    12,     2,    -8,   -21,     7,    19,    -8,   -25,   -23,   -20,    -3,   -13,     8,   -21,   -16,   -11,    12,    20,    -3,     8,    17,   -11,    -3,     5,   -15,     2,    15,    13,    -6,    -5,   -16,     6,    17,     4,    -6,    -2,   -30,     5,     0,    -4,    -3,    -2,   -15,     8,    20,    22,     4,    -1,     5,   -13,   -21,     8,   -17,     7,     7,    -2,    16,     2,    14,    11,    -1,    -2,   -24,    -5,   -23,    -3,     0,     4,    -4,    12,    -2,    -6,     8,    -7,    11,     1,    11,    10,    22,     7,    11,    12,     2,     8,     0,     8,    14,     4,    -8,    -4,   -20,    -2,    -8,    -2,     1,     3,    10,    -9,   -17,   -23,    -8,    -5,    18,     8,     8,     4,    13,    26,    17,    -9,    -3,     3,   -15,     8,    11,    -8,   -16,     2,    -2,     1,    -4,    -1,    -5,    -3,   -11,    -2,    -3,   -22,   -22,   -20,    17,    20,    14,     7,     3,    -7,    16,     6,     5,    17,    -8,     6,     3,   -22,   -11,     6,    -2,   -23,    -7,     5,     1,    -4,    -4,     4,   -12,   -30,   -15,   -36,   -22,   -33,   -22,   -15,   -21,   -29,   -20,   -12,   -25,   -33,   -21,   -16,    -8,    -6,    -9,    -5,    -2,    -3,     4,    -3,    -1,     4,    -3,    -6,    -5,   -21,   -27,   -25,     0,   -11,     7,    -7,   -20,   -37,   -34,   -35,   -28,   -15,   -22,    -5,    -7,     3,     1,   -12,    -1,     3,     2,    -4,     4,    -3,    -2,    -4,    -7,    -1,    -4,    -7,     0,     2,     1,    -3,    -5,    -6,   -30,   -14,   -10,    -3,    -2,   -12,   -14,   -19,   -19,    -6,    -3,    -3,     0,    -3),
		    16 => (    3,    -4,     4,     0,     4,    -2,    -2,     0,     5,    -1,     0,    -2,     8,     1,    -3,     1,    -1,    -3,     4,     3,    -1,    -1,     1,    -3,    -2,    -2,     3,    -4,    -1,     2,     2,    -3,     2,    -4,     1,    14,     4,     4,     4,     6,    18,     8,   -13,     1,     8,     7,     3,     1,    22,     4,     7,     4,     3,     1,     0,     5,    -2,    -2,     9,     2,     5,     6,     9,    11,    11,    -6,    -8,    -2,   -18,   -14,     8,     7,    30,    34,     3,   -17,   -23,    12,    20,    14,     6,    -6,     0,    -1,    -4,     0,    -5,    -1,     7,    15,    -3,    -2,    -1,   -10,    -7,    -4,   -22,    -6,    15,    17,    31,    13,    -5,     7,    27,    13,   -11,    -4,     2,     0,    -1,    -4,     3,     1,   -14,   -13,    25,    22,    -4,    -5,   -13,    -8,    -7,   -20,   -23,   -10,   -20,     2,    -5,     1,   -13,    -6,     2,   -20,     3,   -18,   -16,    -9,    12,    12,     4,    -1,    -9,    -2,    28,    25,     3,    -3,    -5,    -2,   -26,   -41,   -14,   -25,    -6,    -7,    12,    11,    -8,    -5,   -32,   -26,    -2,   -18,    -3,     0,    11,     5,     2,     0,     2,   -13,    17,    14,    -3,    -1,    -7,   -12,   -36,   -39,   -24,    -5,     5,    21,     2,   -23,    12,    11,    -5,   -32,    -6,    -6,     1,    -2,    -5,     6,     4,    -2,     0,   -25,    12,    17,    -1,   -13,   -10,   -16,   -29,   -38,   -22,     2,     4,   -29,   -17,   -31,   -18,     2,     3,    12,    14,     2,    -4,     7,     2,    -8,    -1,     1,    -4,   -24,    13,    15,     4,    -1,   -15,   -18,   -27,   -41,   -10,     5,     4,   -20,   -11,   -19,   -29,   -19,    -9,    22,     9,    -7,    -5,    -2,   -17,   -24,     2,     0,    -2,   -12,    23,    19,     3,     7,    -9,   -20,   -22,    -5,     7,    11,    -5,     4,   -20,   -14,   -23,   -20,   -19,   -19,   -17,     2,    -5,     2,     0,    -7,     4,    -4,    -8,   -15,    22,    24,    -6,    -9,   -14,    -6,    -4,   -16,    11,     0,    -2,   -32,   -20,   -23,   -41,   -30,   -24,   -28,   -15,     2,     5,     2,    -8,    -4,    -3,     3,     1,   -18,    29,    27,    -5,    -7,   -13,   -22,   -17,     5,    -2,   -11,   -16,   -23,   -15,   -28,   -37,   -30,   -20,   -31,   -24,     5,     7,     2,    -5,   -11,     2,    -1,    -4,   -13,    16,    23,    -7,   -17,   -16,    -8,    -2,    22,     7,   -12,    -9,     0,   -22,   -34,   -24,   -14,   -11,   -28,   -23,    15,    13,     0,   -14,   -10,     2,     1,     5,   -12,    17,    17,    -1,   -10,    -9,   -12,    -2,    10,    -3,    -3,     6,     8,    22,     6,   -12,   -12,    -7,   -21,   -19,     8,   -15,   -19,   -14,     0,     3,     4,    -4,    -3,     0,    13,    10,     2,    -4,   -27,     1,    -2,    -1,    -8,   -15,    -4,    17,   -14,   -23,     0,    12,   -16,   -17,    -3,    -9,    -9,    -9,    -5,     5,     0,    -5,   -15,    -5,     4,     6,     0,   -11,   -19,    -1,     2,    -1,   -35,    -5,    -5,     6,    22,    -1,    23,    18,   -14,    -4,    -7,   -13,   -14,    -7,   -19,    -2,     5,    -3,   -16,    -6,     7,    -2,    11,     9,   -20,    -2,    25,    22,   -19,    -6,   -24,    -4,     6,   -14,    12,    -1,   -21,    -9,   -16,    -8,    -5,   -10,    -8,     2,     5,     2,   -17,   -11,    -5,     3,     6,     7,   -21,    13,    32,     8,   -36,   -32,   -12,     3,   -14,    -3,    10,    -2,   -17,   -15,    -7,   -14,   -25,    -4,   -14,     4,     0,     0,     4,   -13,     0,     0,     0,   -23,   -18,     1,     4,    14,     1,   -26,   -19,     0,     9,     7,     9,   -27,   -16,   -23,   -19,   -23,   -26,    -4,   -13,     2,    -2,     1,     1,    -6,   -12,   -15,   -15,   -17,   -24,    -3,    26,    15,    16,    -1,    -9,   -17,    12,     5,     6,   -16,   -11,   -20,   -18,   -19,   -14,   -14,    -6,     3,    -3,    -4,    -4,    -1,    -8,   -12,   -19,   -21,   -32,   -27,    -3,     8,    17,    -4,     1,    -6,    19,    -3,    10,     6,   -11,    -9,   -10,    -7,    -7,    -2,     0,    -2,     1,     3,    -2,     4,    -4,    -6,   -14,   -18,   -29,   -27,   -27,     0,    13,     2,    -4,   -10,    -5,     0,    -2,   -23,   -13,    -7,    -6,   -11,   -13,    -1,     3,     4,     0,     0,    -7,     1,    -5,     5,     0,   -14,   -32,     4,   -11,     0,     4,    15,    16,   -10,   -23,   -26,     8,    -5,    -7,     2,    -7,   -20,    -5,     4,     2,     3,    -4,    -3,    -7,     2,    -3,     0,    -5,    -5,   -21,   -25,   -14,     4,    -7,     2,    -7,    -9,   -10,    -2,     3,   -10,    -7,     2,    -2,    -2,    -6,     4,     1,     4,     2,     0,    -5,    -7,    -8,    -6,     0,   -12,    -7,   -13,     4,     7,     7,     0,    22,    38,    16,   -25,   -38,   -10,    -1,    -1,    -2,    -3,    -7,     0,     1,     2,    -5,     0,    -4,     3,    -5,    -4,    -4,     1,    -7,    -5,     2,    11,     7,    -5,    -2,    -7,    -3,    -4,    -7,   -13,    -2,    -6,    -8,     1,     4,     3,     1,    -1,     2,     2,     1,    -2,    -2,     4,     2,     2,    -1,    -4,    -6,    -3,     2,     3,    -5,     1,     0,     2,    -4,    -2,    -8,     1,    -1,     4,     4,    -5,     3,    -2,    -3,     4,     4,     1,    -1,    -4,    -2,     2,    -3,    -2,     3,     0,     1,     1,    -6,    -3,     0,     3,    -2,     1,     1,     2,    -3,     4,     0,     0,     0),
		    17 => (   -1,     1,    -3,     3,     0,    -3,    -4,    -5,     3,     3,    -4,     4,     1,     5,     4,    -4,    -1,    -3,     4,    -2,    -3,     2,    -3,     5,    -2,     1,     1,     3,    -2,     0,     5,    -1,     5,     4,     1,    -2,    -2,     2,    -4,   -20,   -18,   -13,    -3,   -15,   -17,   -12,     1,     2,     3,     3,     0,    -3,     5,     1,     2,    -1,    -1,     3,     1,   -11,    -8,     1,    -5,    -1,    -7,    -5,    -5,   -15,    -9,    -8,     0,   -11,   -12,    -2,    -2,     3,    -3,     1,    -5,     0,     4,     2,     5,    -1,     3,     0,     3,   -17,    -3,    -6,    -7,   -13,   -18,   -14,   -11,    -8,    -9,   -13,    -7,   -14,    -4,    -4,    -7,    -5,    -5,    -8,   -23,   -10,    -1,    -7,     5,    -4,     2,    -1,    -4,    -2,   -23,   -11,    -3,   -31,   -30,   -15,   -31,   -51,   -44,   -40,   -31,   -16,    -9,    -2,     2,    -3,   -20,   -24,   -13,   -25,    -6,   -11,    -6,     1,     3,     5,    -2,    -5,   -24,   -12,    -8,     7,     6,    -4,   -20,   -12,     3,     1,   -27,   -33,   -37,   -68,   -78,   -73,   -69,   -41,    -4,   -25,   -16,   -12,    -5,    -3,    -4,     4,    24,    25,    -2,    -4,    -1,   -13,   -12,   -23,   -32,    11,    18,    10,   -11,   -40,   -30,     0,    -4,    -3,    -9,    25,    15,     5,   -18,   -20,   -33,   -10,    -4,    47,    43,    28,     4,    -4,     0,    21,    -5,     0,     4,   -13,    10,    -3,   -14,   -21,   -21,    -6,    -2,    -7,   -16,     3,    -5,    12,    10,    -2,   -25,   -11,   -30,    50,    15,     5,   -10,   -16,   -13,    -5,   -21,    -3,    20,     2,     8,   -17,   -14,    -9,   -14,     9,    11,     1,    -6,   -18,    -8,    19,    31,     9,   -19,   -16,     2,    28,   -21,    -2,     8,     1,    12,    -5,   -11,     4,     4,    10,     5,     1,    22,    -2,   -14,     8,    17,    14,     3,     5,     5,    11,    35,    -5,   -32,    -1,     4,    21,    15,     4,     9,     4,    19,     8,     9,    -1,     2,    19,    18,    25,    -2,   -21,   -15,     7,     0,    13,    20,    18,   -14,   -10,   -15,   -11,   -26,     8,    -1,     4,    18,    23,     9,    28,     6,   -11,   -20,    20,     7,    34,    38,    -2,   -31,   -20,   -12,    -5,    28,    14,    19,    -7,   -18,     0,    -9,   -22,   -11,     4,     5,     7,    11,    15,     2,    14,     6,    21,    13,    10,    22,    12,    23,   -61,   -66,   -11,    10,     9,    15,     0,     8,    -9,   -20,   -20,   -12,   -16,    -3,    14,     1,     8,    23,    -6,    -5,    23,    16,    22,    18,    -3,     3,     2,   -14,   -84,   -57,   -29,    13,    -2,    16,   -14,     0,     9,   -18,   -33,    -2,   -27,    -7,    -4,    -5,    16,    44,    17,   -12,    26,     8,    -7,    -3,    17,    25,     6,   -39,  -110,   -51,   -19,    11,    -3,    22,    12,    -3,    -5,    -5,    -3,     1,   -16,   -12,    -3,    -5,     0,    12,    17,   -40,    10,    15,    13,   -18,   -11,    28,   -14,   -96,   -67,   -36,   -15,    14,    13,     9,    20,     1,    -7,     2,   -16,   -22,   -22,    -2,    -8,    -6,    -6,     7,     6,   -20,   -15,     3,    27,    -4,    -2,    31,   -41,   -93,   -12,     1,    -6,    -7,     4,    17,    16,   -19,    -2,    13,   -12,   -12,   -20,    -1,   -19,    -5,     2,    13,    -7,     3,   -13,     4,    -2,   -16,   -31,   -47,   -64,   -51,    -5,     6,    -4,    -6,   -11,    16,   -14,     5,    -3,    15,   -47,   -62,   -10,     0,   -23,    11,    -4,    27,   -41,   -17,    -4,    10,     2,   -24,   -48,   -80,   -21,    -7,    13,    23,    -4,     8,    11,    11,   -13,    15,   -11,   -17,   -60,   -57,     6,     0,    -7,    -4,    15,    10,   -33,    -5,     6,     8,   -50,   -50,   -59,   -62,   -20,    -2,     1,     5,    -1,    -7,   -12,     9,     1,    -9,   -24,   -38,   -44,   -27,    19,    -1,    -5,     0,    18,    -2,   -19,   -11,   -11,   -20,   -48,   -48,   -63,   -14,    23,    16,   -12,     0,   -16,   -11,     3,   -13,    -4,   -16,   -38,   -33,   -47,   -17,     1,    -2,    -1,    -3,     0,    -7,   -23,   -46,   -12,   -42,   -39,   -36,   -14,    32,    10,   -11,   -17,   -10,   -29,   -16,    -2,    13,     3,    -2,    -8,    -1,    -7,    62,     3,    -5,     2,     0,     5,    -5,   -12,   -30,     3,     3,     0,     5,    11,     2,     7,   -13,     0,     3,     1,    -6,     3,     6,    12,     3,   -10,    -1,    -7,    -4,    -1,   -13,    -2,     2,     2,    -5,   -30,   -16,    17,    22,    14,    15,    -1,     8,   -32,     1,    10,     0,     0,   -13,   -10,    11,   -20,   -10,    -4,   -43,   -27,    -5,    -9,    -4,    -3,    -3,     0,     7,     7,    -1,    21,    -8,   -24,    15,    -2,     4,     8,     6,     0,    14,    -8,   -13,   -10,   -31,   -19,    -9,     7,   -35,   -35,    -8,   -29,     4,     1,     3,     0,    -4,    -1,   -35,   -44,   -17,   -12,     0,    -4,     7,     6,    10,     2,    15,    -1,     9,    13,   -21,    -7,    -9,     9,    -2,   -22,    10,    -5,    -4,     2,     2,     1,     4,    -2,   -39,   -36,   -30,   -32,   -13,   -20,   -19,   -24,     4,    19,    21,     3,    13,    -6,     0,     9,    -8,   -10,    -6,     0,   -10,     3,     0,     1,     4,     4,     2,    -2,    12,    11,     4,    10,    19,     7,    11,     5,    -6,    -4,     5,   -10,   -11,    23,    22,   -18,    11,    35,     9,    19,    -2,     4,     0,     0),
		    18 => (    3,    -4,     1,     0,     4,     0,     1,    -4,    -1,    -3,    -5,    -3,    -1,     4,    -2,     2,     2,     1,    -2,    -4,     1,     3,    -4,    -4,     1,     2,    -4,     2,     3,    -4,    -1,    -2,    -3,     4,    -3,    -2,     3,    -4,     2,     1,    -5,    -8,   -12,   -22,   -35,   -16,    -6,    -8,    -6,   -11,    -9,     0,     4,     4,    -3,     0,     4,    -1,    -6,     0,     0,    -2,   -13,    -8,   -10,   -29,   -37,   -20,    -5,     1,    -7,   -25,   -16,    -6,     7,   -13,   -39,   -32,   -36,   -11,    -8,    -7,     4,     3,    -3,     2,   -15,   -16,     0,   -13,   -17,   -41,     7,     4,    -5,   -17,   -19,   -29,   -43,    -2,     6,     4,    15,     9,    36,    30,    13,    12,   -13,    -5,   -11,     1,    -1,     4,    -2,   -25,   -23,   -38,    -1,     0,   -16,   -26,     4,   -12,   -34,   -28,    14,     1,     5,    -5,    -5,    12,    26,    29,    17,    11,     0,    36,    16,    -6,    -4,     2,   -19,   -26,   -39,   -13,    -2,     3,    10,    -3,    -1,     0,   -14,   -13,   -12,     4,     0,   -16,   -21,    -8,    26,    14,     7,    33,    33,    15,   -13,    -1,     1,     1,   -14,   -23,    -6,   -21,     6,     9,    10,    -3,    -7,   -13,     9,    -1,     5,    -1,   -23,   -25,    -8,    13,     1,   -11,   -24,     8,    -3,    40,     3,   -20,    -2,   -27,   -15,    -5,    -1,   -24,     9,    27,    -1,   -14,   -10,    -6,     2,     0,     3,     9,   -23,    -5,    17,     7,   -13,     2,    11,    12,     9,    -3,    -4,   -23,    -9,    -8,   -15,     8,    26,   -10,    19,    20,   -19,    10,    -5,     3,     4,    21,   -10,   -33,   -14,   -11,   -12,   -27,     3,    24,    14,    -3,     5,    16,    14,     7,    -2,     5,    -4,    16,     8,   -24,   -10,    -7,   -11,    -8,     8,    19,    -7,    -8,   -24,   -33,    -1,    -5,   -19,     9,    10,     8,     4,    20,     4,     5,   -23,   -54,     2,    -5,    -7,   -16,    -2,   -23,   -17,   -27,     5,    15,    19,     4,    -5,   -19,   -21,   -20,     4,    20,    -8,   -10,    -6,    -9,     0,    13,     1,   -38,   -20,   -42,    -1,    -4,   -15,   -20,   -20,   -14,    -7,     3,   -12,    14,     0,    23,    19,    -4,    -8,   -14,    -1,   -11,    -8,   -34,   -17,   -40,   -19,    18,    35,     4,    32,   -25,     1,     2,   -23,    26,   -13,    24,     3,     7,   -23,   -11,     0,   -17,    10,    18,    -4,   -14,   -15,     0,     6,    15,   -24,    -6,    21,    42,    40,    12,     9,   -44,     0,    -1,   -22,    21,    -7,   -13,   -41,   -16,   -19,   -21,    -4,    -4,     4,    11,     3,    -4,   -27,     6,    -3,    11,    15,    34,    49,    43,    21,   -12,   -13,     7,    -7,     0,    -1,   -36,     0,   -34,   -17,   -16,   -28,   -35,    -1,   -15,     0,    22,     7,     3,   -25,    18,   -23,    10,     0,    23,     4,    35,    21,   -12,   -29,     0,     0,     3,    -5,    13,    -4,     8,     3,   -10,     1,   -31,    -8,     4,    13,     6,    -1,   -10,    14,   -43,   -15,     7,   -15,   -31,    -8,    25,    26,     0,   -36,   -24,    -1,    -4,   -10,    18,   -25,    24,    -6,     6,   -20,   -23,   -11,    -3,    21,     4,    -3,     5,   -21,   -10,    -8,   -27,   -35,   -26,   -18,    13,     5,     9,   -27,   -20,    -1,    -3,   -11,    11,   -37,    -6,    -3,    15,   -12,   -18,     2,    16,    18,   -13,    20,    18,    -7,    -6,   -36,   -30,   -15,   -27,   -17,     0,    -3,     3,    -5,   -13,    -8,    -3,    -5,   -14,   -26,   -12,    -7,   -16,   -19,    19,    14,    28,   -13,   -44,    -9,    21,     1,    -5,   -10,    11,    -8,   -44,   -11,     2,   -28,     3,    -2,   -14,     2,    -4,   -10,   -10,   -30,   -12,   -11,   -26,    21,     7,    23,    22,   -21,   -41,   -19,     7,     5,    16,   -19,    -5,   -13,   -26,    -2,   -17,   -19,     1,   -17,    -7,     0,     4,    -5,   -13,   -45,    -5,   -22,    15,    11,    10,    20,    26,     4,   -12,    -5,     3,     1,   -11,     0,     3,   -14,   -13,   -14,   -18,     0,     5,   -21,     2,    -4,   -15,   -12,    -2,   -38,   -46,     4,     8,     9,     9,     2,    -3,     8,   -19,   -17,    10,   -22,   -11,     7,   -11,   -43,   -24,    -3,   -16,    -7,    11,   -25,     0,    -6,    -5,    -7,   -18,   -27,   -55,   -26,     7,    -7,     3,    -1,    12,    -5,    12,   -15,    -4,   -40,     0,     4,   -38,   -59,   -27,   -16,   -16,     3,    13,   -35,    -1,     1,     1,   -14,   -25,   -31,   -38,   -14,     1,    22,   -15,   -25,     3,    12,     6,     8,   -19,    -6,    24,   -26,   -57,   -52,   -24,   -25,    -8,    12,    10,   -34,     2,    -2,    -1,    -4,    -3,   -34,   -46,   -25,    -2,    12,     1,    -3,     5,    21,    21,    11,    -5,    10,   -19,   -28,   -34,   -17,   -13,   -16,    -5,   -13,   -28,   -26,     1,     0,    -2,   -17,   -10,   -16,   -24,    -9,    -5,   -19,   -19,    21,   -25,   -29,   -12,    -5,    14,   -10,     0,     8,    16,    15,    -7,   -17,    -8,   -23,   -12,   -13,    -2,    -2,    -1,     4,    -3,    -6,   -18,   -27,    -3,     2,   -15,   -36,   -26,   -21,   -28,   -41,   -38,   -15,    -7,    -2,    -8,   -14,   -15,   -14,    -4,    -2,     2,     4,     2,    -1,     1,    -4,     3,    -9,    -3,    -1,   -13,   -15,    -7,    -7,    -7,    -3,   -10,    -8,     1,    -3,    -4,     1,    -2,    -3,    -3,    -5,     2,    -1,    -3,     4,    -1),
		    19 => (   -2,     2,    -1,    -2,     0,     1,     0,    -3,     3,     5,    -2,    -3,    -3,    -2,     4,     0,     4,     3,    -1,    -1,     2,     2,     0,    -2,    -4,     1,    -5,     5,     2,     4,    -3,    -1,     3,    -1,     5,    -3,    -5,    -4,     0,     6,    -6,    -7,     0,   -12,   -11,   -16,    -6,    -5,     1,    -6,    -1,     1,     4,     3,    -4,    -1,    -4,     4,     5,    -1,     0,    -1,    -2,    -1,    -1,    -6,    -3,    -4,     2,    -2,   -12,    -6,    -1,    -4,   -11,    -2,    -9,     3,    -3,    -5,    -5,    -5,    -3,     4,     1,     3,    -3,    -1,    -5,   -22,    -1,    -3,   -16,    -1,    -3,    -1,    -2,    -1,   -14,   -32,   -16,     7,    33,    12,   -19,    -9,   -11,    -1,    -3,    -7,    -4,     4,    -4,    -1,    -5,    -6,    -1,   -12,   -13,     0,    -6,     2,     4,    -4,   -17,   -22,   -29,   -46,   -51,   -52,   -31,   -38,   -46,   -24,   -23,   -28,   -18,   -26,   -13,    -3,     2,     2,    -9,    -3,    -5,    -3,    -6,    -2,   -21,    -3,    -9,   -19,   -44,   -50,   -65,   -64,   -51,   -43,   -14,   -13,     2,    -6,   -19,   -37,   -27,   -20,   -24,     3,    -3,    -8,   -15,   -15,    10,    -2,   -13,   -14,   -16,   -34,   -27,   -60,   -67,   -36,    -2,    -8,    -3,    21,    17,   -16,    -5,   -10,   -21,   -33,   -18,   -16,   -20,   -23,     2,   -13,   -18,    -8,   -11,    -8,   -15,   -21,    -8,   -47,   -67,   -39,   -13,    10,    10,    29,    25,   -13,    14,    -2,    19,   -15,    -9,     9,   -28,   -20,   -17,   -13,   -21,   -14,   -16,     3,    -5,     0,    31,   -13,    -2,   -21,   -27,   -14,     9,    11,   -11,   -19,    -1,     5,     8,    16,   -28,     1,    24,    17,   -32,   -33,   -17,    -6,    -1,   -15,    16,    15,    18,     4,    -6,   -14,   -38,   -12,     6,    11,    14,     0,   -26,    -1,   -28,   -47,   -16,     0,   -16,   -15,    39,   -15,   -17,   -35,    -6,   -14,     1,   -21,   -38,    17,    20,     6,   -17,   -32,   -14,     9,    11,    20,     6,     4,     3,    -2,   -22,   -27,    -1,    -1,    -9,     3,     0,   -17,    -7,   -28,   -22,   -13,     1,    -9,   -15,     3,    -4,    -3,   -10,    -2,   -13,   -11,    -3,    18,     2,    12,     0,    -3,     6,   -11,    17,     2,    -8,     3,     5,   -12,    -8,   -11,   -23,   -12,     0,     0,     9,     3,     7,   -17,   -20,    -2,    -3,   -12,     8,     4,     6,     1,    42,    27,    18,    -4,     4,   -27,   -50,    -9,   -28,    -8,   -19,   -32,   -26,   -28,     3,   -10,    -9,    -8,    -6,   -12,     2,   -19,     3,    -9,    22,    30,    16,    13,    12,    14,    -8,     1,    -7,   -62,   -58,   -20,   -28,    -8,     2,   -15,   -13,     1,    -6,    -5,   -15,    -9,    -7,    -5,    -7,     4,   -15,   -15,     2,     4,     0,     4,    19,     7,    -3,    -4,     0,   -52,   -36,   -26,   -16,   -10,     3,     0,    -1,    -4,    -3,    -2,   -20,    -5,    -9,   -20,    -2,    -1,     4,   -12,    10,     4,     7,     8,    15,    10,    25,     9,    15,   -69,   -46,   -14,   -21,     9,    10,    -7,    28,     4,     1,    -4,   -14,    -1,    -5,   -42,   -30,   -11,     2,     2,    39,    17,    15,   -17,   -12,    -2,     2,     4,   -58,   -80,   -24,    21,     7,     2,    32,   -19,    -7,     2,     3,    -7,   -11,    -5,    -7,   -37,   -35,   -19,   -24,   -12,    17,     8,   -24,     0,    19,    -2,   -12,   -16,   -37,   -37,    13,    27,   -23,   -14,    25,    -9,   -21,    -1,    14,    -2,   -13,    -9,   -14,   -15,   -11,   -49,   -52,   -20,    -3,   -11,   -30,     6,    11,    10,   -26,   -19,   -31,   -32,    24,    24,     3,    -6,    -1,     2,   -25,   -15,     0,   -13,   -16,    -7,   -22,   -30,   -24,   -37,   -64,   -51,   -39,   -37,    -4,     3,    -7,    -4,   -26,   -13,   -35,    -7,    12,    32,     4,   -11,    -6,     0,   -10,   -13,    -2,     1,   -12,   -12,   -22,    -3,   -14,   -42,   -31,   -16,   -23,     0,     0,   -14,    -2,   -29,   -21,   -20,   -26,    19,     6,    -6,    -5,    -7,    19,    11,    -4,    -3,    -5,     0,   -15,   -15,   -19,    -9,     7,    -8,     3,    -3,    -3,   -13,     3,    -5,    -8,     1,   -10,   -30,   -17,    21,    21,    -2,     0,    22,   -33,    21,   -14,    -5,     0,     3,   -11,   -23,    -2,     7,   -15,     2,     9,     2,   -11,     4,   -18,   -26,   -14,   -12,   -13,   -40,   -16,    15,    30,    -1,    -9,    20,    30,    -1,     2,    -3,    -3,    -3,    -8,    -7,   -23,     4,    -7,    21,     4,     6,     3,   -21,    -7,   -15,   -20,   -27,   -16,   -25,   -21,    11,    37,     5,    -1,    -8,    21,   -15,     2,     2,     0,     0,    -5,   -16,   -11,     9,     2,    15,    -3,     4,    -5,   -18,    -2,   -13,   -16,   -21,   -12,    -9,   -32,   -18,    12,    -3,    -1,     2,   -21,   -13,   -17,    -4,    -5,    -1,    14,    -5,    24,    -7,     1,    18,     2,   -25,   -15,    15,    -9,     8,   -19,   -13,    43,    14,   -18,   -11,     7,     8,    -6,     7,   -26,   -22,   -16,     1,    -5,    -2,     2,    28,    31,     3,    -4,    19,    -5,    12,   -11,    17,    30,    13,    28,     6,    53,    48,     2,   -33,     2,    12,    -9,    -8,     1,    -5,     0,    -4,    -5,     5,    -1,    -2,    -1,    -3,     3,     2,     1,     2,    17,    34,    29,    29,    37,    22,    13,    -6,   -10,    -6,   -10,    -8,     2,    -5,     2,     1,     2,     4),
		    20 => (    1,    -4,    -2,     0,    -4,    -5,     3,     4,    -1,     3,     1,    -5,    -4,    -6,    -4,    -6,    -2,     3,     3,     5,    -4,    -1,    -4,    -2,    -2,     0,     5,    -3,    -5,    -5,    -2,     1,     4,     5,     0,    -9,   -15,   -20,   -21,     6,     5,     1,    -2,    18,    11,    10,    -5,    -2,    -2,    -1,    -5,    -2,    -4,     2,    -4,    -2,     1,     3,    -1,     7,    14,    -5,    -7,    -2,   -11,   -20,   -13,    -2,     2,    -8,   -22,   -17,     2,    -1,     3,    -4,    -1,    -5,   -21,   -18,    -7,    -7,     1,     4,     0,     3,    -4,     8,     1,   -18,   -11,    -4,   -21,   -39,   -13,   -14,   -13,   -31,   -22,    -9,    -9,     3,   -10,    -6,   -26,   -25,   -19,   -31,   -13,   -15,   -22,     1,     2,     0,    -8,   -14,   -13,   -34,   -12,    -8,   -11,    -7,     0,     1,   -20,   -16,   -13,    -7,    11,    17,    12,    12,    -7,   -19,   -16,   -19,     2,   -38,   -16,     5,     1,    -1,   -11,    -5,     6,   -17,    -7,   -20,   -19,    -1,     5,     3,    -7,   -12,     3,     8,    25,    19,    24,    12,    -7,    -5,   -30,   -23,    -3,   -34,   -17,     0,    -1,    -3,   -13,     0,    -3,     0,    -3,    -8,   -21,   -17,    -5,    -6,   -14,     2,    -5,    13,    17,    16,    20,    10,    20,     9,     0,    -3,   -10,   -21,    -6,    12,    -4,   -15,   -23,   -16,   -11,    -7,     1,     3,   -24,   -12,    -7,    -3,    -6,     2,     9,     1,     4,    12,     3,     8,    12,    -7,     9,     2,     0,     9,   -19,     3,     9,   -30,     4,   -13,   -18,    -9,   -20,   -11,   -21,   -15,   -13,    -1,     1,    -2,    -7,   -14,    -8,     2,    10,    -4,     3,    12,     3,     2,    -3,   -13,   -18,    -4,    -6,    -6,     5,    -3,   -18,   -17,   -30,    -7,   -19,   -15,   -19,    -1,    -7,   -10,   -26,   -21,   -11,   -18,   -24,   -23,   -15,   -15,   -11,   -11,    -5,   -26,   -28,     0,    -4,     4,    14,    -1,   -20,   -27,   -12,    -1,   -18,   -19,   -24,   -28,   -32,   -31,   -15,   -21,   -14,   -10,   -22,   -20,   -37,   -40,   -12,    -9,   -15,   -11,   -21,    -4,    -3,    23,   -23,     3,   -17,    -7,     9,   -11,   -32,   -24,   -24,   -26,   -25,   -15,   -16,    -8,   -15,   -10,    -9,    -6,   -14,   -19,    -3,    -9,    -7,   -11,    -8,    -4,    -2,     4,   -30,     8,   -10,    -2,    -2,   -12,   -11,    -3,    -9,    -2,     2,     4,     3,    -4,    -1,    -5,     6,     2,     2,    -2,     4,    -6,    -8,   -15,   -13,    -7,     1,     7,    -1,     5,    -2,    -4,     3,    -6,   -15,    -1,   -12,    -6,    -4,     3,    -1,   -17,    -9,     0,    17,     2,   -15,     1,     4,     6,    -2,    -3,   -21,   -15,     2,    -2,    -7,   -19,     3,    -1,    -3,     5,     5,    -3,   -27,   -17,   -13,   -10,   -29,   -24,   -18,    -3,    -2,   -19,    -7,    -4,    -1,   -15,    -6,    14,   -23,    -3,     3,     3,    -6,   -27,     9,     7,   -17,     5,     6,   -19,   -27,   -31,   -19,   -46,   -46,   -21,   -16,     0,    -4,    -4,     9,     1,   -13,   -19,    -4,     3,   -29,   -10,     4,    -1,   -15,    -5,    21,     0,   -16,   -18,    -3,   -28,   -36,   -26,   -37,   -43,   -28,    -1,     1,    11,     4,     0,    13,    -8,   -13,    -2,     9,     8,   -38,     6,    -1,    -2,   -16,    -4,     5,     0,     6,     3,    -3,    -2,   -23,   -21,   -12,   -13,    -8,    12,     6,    14,    -3,     8,    -5,   -11,    -7,    11,     8,     3,   -35,     7,    -7,    -3,   -12,    -4,     9,    -6,     5,     5,     6,     5,    -6,   -17,   -22,   -16,    -1,    19,    14,    11,    -2,   -10,   -10,    -9,     3,     9,     2,    -2,   -21,   -14,     2,     3,     0,    -1,     3,     3,    -5,    15,     9,     9,    -6,    -6,    -1,   -19,     0,    12,     1,   -20,   -30,   -19,    -2,    18,     9,     3,    18,   -33,   -13,   -11,    -3,     8,     8,     4,     2,     4,    -7,    -6,    -4,    -8,    -1,    -8,    -9,   -17,    -3,    -1,   -12,   -25,   -11,    -3,    -2,    -5,    -2,    10,     9,   -10,    -5,    -5,     4,     3,    -7,     0,    -3,    -2,    -6,    -4,     1,    -1,    -7,   -24,   -16,   -28,   -13,     3,   -10,   -13,     1,     3,     3,   -17,    -4,    11,    10,     0,     7,     3,     0,    -5,   -19,     0,    10,     1,    -2,    -3,    -4,    -2,   -21,    -7,   -11,    -6,    -1,   -20,    -3,   -17,     0,     0,   -11,    -1,     9,     5,     3,    -5,     1,     2,    -4,     0,   -17,   -16,   -14,    -9,    -5,    -5,   -22,   -17,    -5,     4,     3,     2,   -11,    -8,    -6,     3,     9,     5,    -6,     9,    11,     4,   -27,   -19,   -11,     1,    -3,     2,    -2,   -12,   -14,     7,   -21,    -8,    -9,   -17,   -38,   -27,   -20,   -19,   -23,   -16,   -11,     6,    -3,    -1,    -8,    -7,    -7,   -11,   -10,    -3,    -3,     3,    -3,     2,     1,   -15,   -26,   -15,   -15,   -13,   -13,   -10,   -16,   -28,   -30,   -36,   -32,   -23,   -25,   -10,    -7,   -30,   -19,   -18,   -21,   -12,     1,    -1,     4,    -2,     1,    -3,    -4,     3,   -19,   -25,   -30,   -14,   -10,   -18,   -19,    -4,    -9,   -18,   -17,   -24,   -21,   -30,   -31,   -34,   -25,   -24,   -19,    -7,     4,     1,     0,     1,     0,    -1,     1,     0,    -1,     2,    -9,   -16,   -15,   -11,    -2,     2,    -2,   -11,     3,    -6,    -7,   -12,    -8,   -12,    -4,    -9,   -12,    -7,    -3,    -1,     5,    -4),
		    21 => (    4,    -2,    -5,     2,    -3,    -4,     2,    -4,    -4,    -4,    -4,     5,     4,     4,     0,     3,    -1,    -4,     3,    -1,     3,    -1,    -2,     0,     4,     0,    -2,    -5,     3,     3,     2,     4,    -3,     1,     3,    -1,     5,    -2,    -4,     4,     0,   -12,    22,    23,    -4,   -18,    -7,   -10,     1,    -3,    -2,     4,     3,     2,    -3,    -5,     2,     1,     1,    -4,    -5,     1,    -3,    -2,    -4,   -24,   -23,   -16,   -39,   -11,   -22,   -21,    -4,   -21,   -11,    -6,    -7,   -28,   -35,   -20,   -15,    -7,     2,    -2,    -1,    -5,    35,    22,    -3,   -19,    -4,    22,    19,    22,     6,   -31,   -21,    29,    -5,   -28,   -22,    -8,    -9,   -18,    -6,   -48,   -32,   -20,   -18,    -6,     4,     3,    -4,    -5,    31,    30,     4,   -10,    -1,    29,    29,    26,    18,    -8,    -3,    10,    -3,     0,   -23,   -24,    -7,     2,   -13,   -32,   -16,   -17,   -17,   -36,   -38,   -29,    -3,     1,    28,     4,     8,    15,    15,    29,    10,    23,    38,    39,    20,    20,     3,   -11,   -13,    -9,   -14,     5,   -11,   -23,   -18,    14,     3,   -60,   -27,   -25,     0,     1,   -13,     2,    13,     5,    19,    35,     9,    11,    43,    19,     7,    15,     3,     0,    -6,     0,    -2,     1,    -3,   -21,   -13,    16,     1,   -27,   -33,   -16,    -2,   -25,   -34,   -29,   -43,    17,    26,    42,   -13,   -16,    19,     6,    18,    -9,    19,     0,     9,     7,   -19,   -15,    14,   -12,    16,    14,    -8,   -22,   -54,   -34,    -6,   -24,   -32,   -46,   -44,    -4,    28,    30,   -16,   -35,    17,   -18,     6,    23,    16,    12,     4,    17,    22,     8,    -8,    -3,    11,    -4,   -27,   -23,   -58,   -23,     4,   -10,   -32,   -44,   -31,   -15,     0,    21,    -8,   -10,   -20,   -27,   -11,    28,     5,     6,    -3,    21,    29,    -6,     4,     9,     2,   -16,   -23,   -24,   -22,   -33,     1,   -15,   -28,   -41,   -33,   -20,   -19,     1,    14,   -16,   -23,   -28,    -6,    17,     0,    -2,    28,    32,     9,    -6,    -2,   -15,   -19,   -28,   -32,   -20,   -36,     3,     0,    -2,   -11,   -25,     2,    -7,   -11,    27,    10,     2,   -14,   -20,    -5,     6,     1,     4,    36,    53,    15,    -1,    22,   -26,   -34,   -27,   -34,   -29,   -36,    30,     2,     4,   -43,   -18,    -3,     4,    23,    24,     5,   -13,   -12,    -1,    10,    -1,    11,    23,    23,    31,    20,    -6,     3,   -30,   -31,    -8,   -33,   -11,     3,    28,     1,    -5,   -22,     1,   -13,    12,    22,    10,   -13,   -22,    -9,   -13,    -5,   -10,     1,    -8,     2,    38,   -19,     3,    -1,   -23,   -24,   -48,   -38,     9,    23,     2,     1,    -4,     3,     8,   -17,     4,   -15,   -20,     0,   -15,   -21,     6,    -5,    -5,    19,    -2,   -10,    -3,   -42,   -14,     7,    -8,    -9,   -19,   -34,    13,    40,     0,     2,    -4,     3,   -12,   -32,   -22,   -11,     0,    -9,    -3,     6,   -15,    -1,     3,    11,     2,   -12,   -24,   -41,   -29,    -8,     6,   -31,   -32,   -45,   -17,    -2,    -9,    -1,    -1,     6,   -30,   -27,     6,     2,   -20,   -20,    13,     1,   -11,    -1,    16,    14,   -24,   -40,   -40,   -12,   -16,     1,    -1,    -7,    -2,    16,     2,   -13,    -9,     0,    -4,    -7,   -45,   -23,    11,    -5,   -15,   -15,   -25,   -20,    15,    17,    12,    17,   -38,   -32,   -42,   -28,    -3,     6,    15,    26,    28,    23,     0,   -20,   -26,    -5,    -3,   -12,   -44,   -30,   -28,   -48,   -31,   -26,   -17,   -11,     0,    -5,     5,     2,   -12,   -24,   -23,    24,    26,    29,    25,     5,    -3,    11,    18,   -14,    10,     4,     0,     6,   -52,   -39,   -13,    -7,    -6,    -3,     4,    15,    15,   -12,   -17,    12,    -7,    -9,     1,     3,    17,    48,    25,     3,    21,    28,    23,    -9,     3,    -4,    -1,   -24,   -43,    -8,    -3,    13,    -6,    10,    22,    31,    10,    -2,   -11,    -8,     3,    -1,    13,    31,    29,    45,    16,     2,    -3,    12,     8,    -2,     0,    10,     8,   -35,    -2,    -8,     9,    -3,     3,    -4,    11,    21,   -11,   -25,   -17,   -10,    17,    11,    -6,    37,    35,    42,    35,    -5,    -9,    15,    11,   -14,     1,     4,     3,   -30,   -24,   -10,     9,    -4,    -7,    20,     6,     9,    -9,   -18,     0,   -18,    21,    -5,    10,    61,    40,    25,    36,     8,     0,    14,    21,    -4,     1,    -3,     4,   -10,    -3,   -23,    -6,     3,     3,   -26,    -6,   -12,    -2,    25,     7,    13,    40,    16,    24,    29,    19,    27,     8,    -2,   -22,   -30,   -18,    18,    -5,    -2,    -4,     1,    -5,   -26,   -23,   -25,    -3,   -32,   -36,     8,   -18,     3,     5,     4,    19,    12,    32,    10,    11,     4,    20,     9,   -23,   -20,     9,     5,     2,     2,    -1,    -3,   -13,   -24,   -44,   -50,   -51,   -30,   -75,   -71,   -59,    -7,    -2,   -14,     3,   -27,   -54,   -51,   -63,   -53,   -40,   -16,   -16,   -17,   -15,   -11,     4,     2,     0,    -2,   -11,   -33,   -62,   -57,   -40,   -77,   -75,   -41,   -28,   -38,   -48,    -4,    -5,     9,   -30,   -23,    -8,   -13,   -28,    -3,    -4,     4,     4,    -2,    -2,     4,     3,     0,    -4,    -7,    -9,    -8,     1,    -2,    -7,   -34,   -19,    -7,   -11,   -16,    -9,    -4,    -3,     6,    -5,    -6,     3,    -3,     0,     0,     3,     4,    -5),
		    22 => (    0,    -2,    -2,    -1,     1,    -1,     0,    -4,     3,     2,     1,     2,    -9,   -12,     9,     8,    -1,    -3,     0,    -5,    -4,    -1,     1,    -1,     3,     0,     0,    -4,    -4,     1,     3,     3,     3,    -2,   -12,   -13,   -28,   -22,   -12,   -18,   -13,   -27,    -9,     0,     0,    -5,   -13,   -48,   -28,   -15,   -16,   -11,     5,     1,     0,     5,     0,    -3,    -4,    -9,   -16,    -7,    -4,   -16,    11,    22,    26,    24,    20,    14,   -13,   -10,    -6,   -14,   -25,   -30,   -29,   -17,   -12,    -4,     3,    22,     3,     0,     3,     2,   -10,   -27,   -27,    22,    18,   -15,    -2,    41,    15,    27,    28,     9,     5,    -9,     0,    -3,   -27,   -20,   -10,    18,     0,   -26,     3,     7,    -3,     1,    -2,    -2,    -1,   -10,    22,    -8,     9,    20,    12,    33,    20,    18,    19,    16,    -1,     5,    10,    16,     7,    -4,    -2,   -19,    -9,   -15,   -11,   -14,   -11,   -11,    -2,     3,     8,     5,    17,    14,    -4,    10,    12,     5,    -2,    -1,     1,     4,     7,     8,    29,    10,    21,   -11,    -8,    -5,     7,   -14,   -14,   -13,   -10,   -10,     0,     0,     5,     2,    -1,     9,    -8,     3,    20,     7,     4,    -4,    11,     1,    21,    38,    23,     2,     5,     4,   -24,   -16,   -12,   -27,   -47,    -2,    -7,    -8,    -3,     0,     5,   -14,     2,    -6,    17,    16,    14,    16,     0,     5,     1,    10,     3,   -19,     0,    -4,    -6,    -8,   -19,   -25,   -15,   -46,   -17,     3,   -13,    -3,   -15,    13,   -19,   -21,    -4,   -13,    -5,     1,    -8,    -1,    22,     6,   -18,    -9,    -6,    -6,    -7,     3,    13,    12,     3,    -1,   -30,   -29,   -17,   -17,    -5,   -13,     2,     1,    -4,   -25,   -25,   -32,   -28,   -22,   -34,   -34,    -3,    -4,    -2,   -16,   -22,   -23,    -1,    -9,    -4,   -13,     1,    -9,   -10,   -32,   -37,   -27,     5,    -5,     1,    -1,    -3,   -34,   -21,    -7,     5,   -15,   -30,   -37,   -24,   -33,   -22,   -45,   -32,   -31,   -12,     9,    11,    13,     6,   -16,   -46,   -16,    -5,    -8,    -4,   -12,    -4,   -15,   -14,   -27,   -20,   -33,   -34,   -62,   -53,   -55,   -54,   -53,   -46,   -32,   -32,   -44,   -22,    -3,   -16,    14,    -4,   -13,   -10,    12,    13,    -1,   -32,    -9,    -1,   -22,   -24,   -21,   -44,   -40,   -39,   -61,   -48,   -31,   -27,   -40,   -12,    -1,    -8,   -16,    -8,   -11,    -7,    13,    -7,    -4,    -9,   -16,   -40,     8,   -23,    -6,    -3,   -20,    -8,   -16,   -30,   -34,   -19,    -2,   -10,   -19,   -18,    14,    37,    27,    17,   -12,    -7,     1,    19,    -6,    -4,   -23,   -12,     0,    18,    17,    17,     7,    -4,   -23,   -20,    23,    -5,    -9,     8,    12,    14,    25,    34,    38,    42,     7,    22,     9,    11,     2,    12,    -5,     1,   -15,     0,     3,    22,     4,    21,    24,     1,   -10,    -1,    20,    18,    32,    19,     2,    11,    29,    27,    20,    -5,    -3,    10,    15,     1,    -6,     6,    -5,   -17,     7,    -5,    -8,    -5,    22,    21,    36,    -4,     3,    18,     3,    27,    10,    18,    11,     3,     8,    -5,    13,     0,    -6,     7,     6,    11,    21,    14,    14,    21,    27,    13,     5,    -8,    38,    32,     8,     4,    -1,    15,    -9,     9,    13,    23,     0,    23,     0,    17,    -9,     0,   -24,     6,    15,    -8,    17,    14,     6,    -1,   -16,     8,    -9,   -39,    24,    -5,    19,    -2,     0,   -11,   -31,   -14,    24,    16,    21,    33,    14,     3,   -19,   -25,     0,     6,     7,    14,    -6,   -14,     5,    15,   -16,    20,     3,    11,     1,    -8,    43,    -2,   -13,    -4,   -41,    -9,   -33,     4,     6,    10,     0,    -3,   -29,   -25,   -24,     3,    29,     8,     9,     7,   -16,     0,    -5,     8,   -14,    -1,   -11,    26,    37,    -2,   -20,    17,    -2,     7,     3,   -29,     2,    29,    -4,   -19,    -6,   -13,    -5,   -13,   -14,   -13,   -15,    14,    -9,     2,   -14,    -8,   -19,    22,   -22,    22,     0,     5,     6,    12,    19,    13,    -4,    -1,    -1,     7,    -2,    16,     0,   -13,    -9,   -10,   -36,   -39,   -20,   -16,     3,   -16,    12,     0,     6,   -24,   -21,   -49,    -2,     4,     5,    12,    35,    17,     4,     5,   -20,   -14,     1,    -9,    -3,   -29,   -17,   -44,   -66,   -13,   -28,     4,     1,   -23,   -19,    11,     4,    -6,   -32,   -53,    -1,     4,    -1,     5,     9,    -8,    -7,   -26,   -21,   -13,    -8,     1,   -12,   -16,   -47,   -29,   -40,   -31,   -32,   -19,   -54,   -34,   -24,     4,   -22,   -18,   -28,   -50,     1,    -2,    -2,   -27,   -12,   -31,   -20,   -59,   -28,   -33,   -43,   -47,   -32,   -54,   -63,   -57,   -55,   -39,   -20,   -63,   -64,   -41,   -17,    -7,   -36,     5,     7,     0,    -5,     4,     4,    -1,    -3,    -1,   -10,   -13,   -24,   -39,   -48,   -28,   -20,   -30,   -35,   -32,   -34,   -46,   -51,   -35,   -44,   -34,   -16,   -12,    -1,    11,    20,    22,    -3,     3,     0,     1,    -2,    -4,    -9,    -8,    -5,    -7,   -10,    -1,    -4,     1,    -7,    -5,   -13,   -18,   -21,   -15,    -7,    -9,     4,   -15,    -3,    -9,     5,    -3,    -4,    -5,    -2,     4,    -1,    -4,     4,    -3,    -5,     0,     2,    -4,    -5,    -2,     0,    -7,     1,     0,    -3,    -3,     2,    -5,   -10,    -5,    -1,     5,     0,     4,     2),
		    23 => (    1,    -1,    -2,    -2,     4,    -4,    -1,     1,    -2,     2,     1,     2,    -2,    -7,     2,    -2,     1,     1,    -3,    -4,     1,    -2,    -2,     5,    -4,     5,     1,     2,     2,    -3,     0,     3,    -2,     0,    -1,     2,    -2,    -3,   -12,   -12,   -14,    -8,   -13,   -13,   -13,   -19,   -17,    -7,    -6,    -6,    -5,    -4,     4,     4,     0,    -1,     2,    -2,     3,     5,    -4,    -5,     0,    -5,   -25,   -20,     3,     0,   -15,   -13,   -17,   -25,   -40,   -27,   -20,   -23,   -14,    -7,    -9,   -21,    -1,     3,    -2,    -2,     3,     1,    -7,     8,    -7,    17,    27,    40,    19,    10,   -15,    -4,    -1,     4,   -14,     6,    14,    -8,   -48,   -29,   -10,   -32,   -20,   -34,   -10,    -9,     5,     1,    -3,     8,     2,     6,    21,    22,     4,    14,    31,    22,     2,    -7,     5,     7,     6,    -2,     0,     2,   -28,   -40,   -55,   -22,   -26,   -47,   -27,    -7,    -6,    -1,     5,     2,    15,     3,     6,    19,    15,     2,     4,     0,    12,    14,     4,    20,     3,     6,     8,   -16,   -19,   -12,   -46,   -42,   -53,   -44,   -22,   -19,   -10,    -4,     5,     5,     7,    14,     5,    26,    25,     6,    17,    24,    26,    -7,    -2,    11,     2,     8,     6,     4,    12,    -6,   -14,   -45,   -47,   -43,   -12,   -12,   -24,    -4,    -1,     3,     0,    20,    32,    32,    11,     6,    -6,    -3,     1,    -6,   -13,    13,     4,    -1,    18,    10,    -7,    -6,   -37,   -46,   -48,   -52,   -26,    -3,   -22,   -11,    -9,    -3,     6,    11,     2,    26,    23,    17,    -2,   -37,   -14,   -62,   -40,   -11,   -10,     9,    15,     2,     2,    22,   -30,   -34,   -48,   -53,   -37,   -12,   -25,    -1,     5,    -7,    -5,   -10,    -9,    -7,   -11,   -47,   -76,   -67,   -42,   -43,   -12,    -7,    16,    19,    11,     6,     0,   -31,   -66,   -47,   -43,   -25,   -19,   -12,   -23,     2,    -2,   -13,     7,     1,   -29,   -49,   -85,   -90,   -55,   -20,    19,     2,     4,    16,    23,    -3,    -2,    10,   -29,   -52,   -66,   -52,   -11,     2,   -20,   -10,   -15,    -7,     4,    -7,    -4,    -7,   -52,   -56,   -50,   -38,    25,    16,    21,    36,    19,    25,    12,     0,   -31,   -31,   -23,   -39,   -33,   -32,   -22,     2,   -26,    -6,   -14,    -3,     4,    -7,   -11,   -18,   -17,    -3,    -8,    25,    23,    35,    15,     5,     1,     5,    -5,     9,   -24,   -31,   -15,   -22,   -19,   -21,   -11,   -14,   -24,    -3,   -11,    -5,     3,    -3,    -8,   -16,     1,     8,    22,    54,    36,    14,     0,   -15,     0,    -4,    25,     3,    -1,   -28,   -12,    -7,    -1,    -2,   -15,    -4,   -26,   -24,   -18,   -11,     1,     2,     2,   -19,     4,   -11,    -9,     0,    10,    -4,    -5,   -14,   -15,     2,     1,   -15,    -7,   -10,   -10,    11,     1,    23,     4,    11,    -1,   -51,    -4,   -14,    -6,    12,     1,   -13,    -3,    -2,    -9,   -39,   -16,   -28,   -16,   -27,   -12,    -2,    -1,   -32,     0,    13,    -4,    -6,    -3,    25,     6,    11,    20,   -28,    -4,    -6,     0,     1,     2,   -16,   -14,   -13,   -29,   -50,   -12,   -30,   -31,   -51,   -73,   -42,   -14,   -22,    -3,    11,     1,    11,     5,    25,    27,    18,    13,   -53,   -43,   -10,    -3,     8,    13,    10,   -16,   -13,    -8,     5,    24,     4,    -9,   -50,   -62,   -46,   -47,   -23,    -1,     8,   -20,   -23,    -5,     7,    12,   -20,   -10,   -54,    -9,   -13,    -5,     9,    -6,    24,    14,    16,    37,   -16,    38,     7,    -8,    -4,   -10,   -22,   -16,   -11,    17,   -13,   -13,    -1,     3,     3,    -2,   -25,   -21,   -27,   -17,   -12,    -4,    -2,   -27,     6,    12,    11,   -10,   -10,    13,    -7,    -9,    14,    25,    21,    -8,    -5,   -23,    -8,    -6,     2,   -11,   -19,     1,    -8,     6,   -16,   -26,   -13,     2,    -3,   -23,     8,   -15,     6,    11,    -6,     8,    12,     0,   -16,   -13,   -14,     2,   -11,     2,    -2,     4,   -17,     3,   -27,   -22,    -8,    10,    -8,   -21,    -5,    -5,     0,     7,     1,     1,     2,     5,     8,     7,    14,     1,    10,    18,     2,   -18,   -18,     4,   -14,    -4,     2,    -7,   -20,    -6,    -7,   -15,    -5,   -14,     0,    -1,     0,     0,    15,    31,     8,    22,     5,     0,     8,     7,     5,    -2,     1,    -2,    -1,   -19,    -8,    -7,     1,    -8,    -3,     7,    10,     8,   -20,    -1,    -4,    -2,     2,    10,    41,    41,     9,     6,    19,     6,     5,     5,     1,   -13,    15,    -7,     2,    -5,   -10,     9,     1,     6,     2,   -15,     3,    17,     2,    -4,     1,     0,    -1,   -10,     7,    -5,    -3,   -29,    14,   -11,   -13,   -11,    10,     0,    -2,    -2,   -11,   -12,   -11,    -4,   -14,   -14,   -24,   -27,   -22,   -14,    -6,     1,    -3,    -3,    -1,     4,    -8,    -6,   -10,    17,    25,    23,    -5,   -10,   -21,   -47,   -19,   -24,   -14,    10,     2,    -2,    20,    -5,   -26,   -37,   -25,     2,    -7,    -4,    -4,     0,    -3,     4,    -9,   -12,   -14,   -11,    -2,   -13,   -21,   -13,   -16,   -27,   -29,   -36,     0,     7,    -7,    -5,     3,   -12,   -18,   -26,     0,     0,    -2,     1,    -1,     1,     2,    -3,     3,    -2,    -4,    -4,    -1,     1,    -6,    -9,   -28,   -17,   -33,    -1,    -7,    -3,     3,    -2,     3,    -7,    -5,   -10,    -5,     5,    -5,     4,     1),
		    24 => (    0,    -1,    -5,     3,     3,    -2,     5,    -2,    -3,     0,    -3,    -2,   -14,   -13,    -7,    -9,    -2,     4,     1,     1,     2,    -5,     1,     4,     3,    -5,     0,    -1,     2,    -1,     1,     4,     1,    -3,   -14,   -16,    -9,   -21,   -28,   -13,   -42,    -7,    14,   -15,   -28,   -17,   -21,    -8,   -16,    -5,    -7,   -17,    -3,     0,    -2,    -2,    -5,     0,    -6,   -45,   -50,   -11,   -17,   -34,   -36,   -24,   -32,   -44,   -44,   -15,    -5,   -32,   -27,   -25,   -16,   -34,   -15,    -7,    -4,     0,     1,    -5,     3,    -1,     4,    -2,    -5,   -38,   -37,     0,   -17,   -36,   -30,   -44,    -4,   -24,   -50,   -30,     1,     1,    18,    12,    13,     1,   -13,    -2,    14,    12,    20,   -12,     1,    -3,    -4,     4,    -2,   -10,     9,   -30,    -4,   -13,   -10,    -2,    -6,     5,   -12,    11,   -19,    -3,     9,    -3,   -17,   -24,    18,    16,    37,    43,    24,     4,   -20,    -6,    -4,     0,    -9,    11,   -16,    -5,   -14,   -21,   -18,   -13,     2,    13,     6,   -11,   -15,   -16,   -33,   -37,   -19,    -8,    12,    -1,    -2,     6,     3,    -1,     2,     3,    -4,    -3,     3,    -7,   -10,     9,   -17,   -27,    -8,    11,     9,   -16,   -20,    -5,   -14,   -11,   -73,   -90,   -39,    -2,    23,     6,    15,     6,   -22,    -9,     2,   -20,    -1,    -4,    -4,   -14,    -6,   -10,   -14,   -12,     6,     3,     2,    -2,     4,     6,    -6,   -46,   -84,   -75,   -22,    14,    11,    21,    40,    28,   -15,   -29,    23,   -17,    -8,   -14,    13,   -10,   -23,   -21,   -14,    -7,    -8,   -24,    -4,   -14,    -8,    13,   -15,   -42,   -74,   -57,   -10,    10,     2,     4,    23,    20,   -12,    -4,    12,   -22,    -1,    -9,    15,   -14,   -14,   -10,    -8,   -14,     3,     4,    -6,   -14,     7,     6,   -29,   -64,   -77,   -46,    -9,    32,    16,    -2,    21,    12,     3,    -3,   -18,    -7,     3,    -1,    12,    19,   -11,   -12,   -20,   -11,     6,     0,    -4,     9,    10,    -3,   -54,   -71,   -48,   -25,    26,    25,     5,    -5,     0,     6,     4,    -7,    -7,   -14,    -2,   -10,    -7,     6,   -11,   -13,    -6,   -12,    -1,   -10,     9,     7,    -3,    -9,   -22,   -45,   -31,    -5,     6,    28,   -10,    -1,     0,     7,    -6,   -14,   -14,   -24,     0,     1,    12,   -15,   -11,   -20,   -11,     4,     4,    -5,    -1,    -2,     9,   -14,   -49,   -27,   -31,    -6,    26,    13,     2,   -13,    -2,     5,   -18,   -22,   -15,   -26,    -4,    -9,    -7,   -15,    -7,    -1,    -4,    -4,    11,    -4,    -3,   -12,     1,   -21,   -23,   -22,   -21,     0,   -11,    -9,    -5,    10,    10,    -4,   -37,    -5,   -16,     0,     0,    -1,   -21,    31,     6,    40,    -6,     8,   -22,    10,     3,     1,   -15,   -23,   -13,   -18,   -13,     1,   -20,     6,    -2,    -8,    -3,   -12,   -14,   -28,    -2,    -2,    -1,     5,    51,    27,     8,    14,   -13,    -3,    -3,    26,    21,     3,   -16,    -7,   -21,   -21,   -20,    11,    -4,    -1,    -3,   -21,    13,    -9,   -49,   -29,   -20,    -7,     3,     5,    17,     1,   -39,    -7,    18,    22,    39,    24,    45,    -2,   -12,     0,   -16,    -5,     3,    -3,     1,     0,     6,     0,    16,   -29,   -28,   -29,   -13,   -14,    -5,    -2,    -3,   -25,   -25,   -12,     9,    26,    36,    19,    29,    14,   -16,    -2,     5,     0,    -4,     5,    31,    21,    11,    19,    12,    -2,   -33,   -21,    12,   -15,    -5,     2,    -2,   -51,     6,     4,    -4,     6,     6,     3,     2,     4,    18,    -3,     9,    15,    10,    16,    21,    15,     8,    12,     8,   -18,   -36,   -21,     0,    -2,     0,     0,    -5,   -33,    -7,    16,    20,     4,    -4,     3,    -8,   -12,   -19,    -6,     1,    15,     1,     0,     8,    21,    -2,   -22,   -12,   -19,    -4,   -36,   -12,    -2,    -2,    -4,     3,   -37,   -30,    -8,   -19,   -15,   -20,   -34,   -37,   -33,    -7,   -15,     7,    -4,   -15,    -7,   -19,    22,     8,   -12,     4,     5,     7,   -28,   -13,     0,     1,     0,    -8,   -30,    -9,   -13,   -15,    -8,   -30,   -57,   -54,   -21,   -15,    -9,     0,   -12,    -2,    -4,    -3,    13,    -4,   -12,    17,    15,    -3,   -32,   -15,    -3,    -4,     1,    -4,   -25,   -29,   -18,   -24,   -34,   -44,   -40,   -43,    20,    -3,   -14,   -18,    -6,    -2,   -14,   -10,     3,   -17,    14,    17,    23,   -14,     3,    -8,    -4,    -3,    -5,    -2,    -7,   -22,   -12,   -24,   -30,   -12,   -11,     0,    16,     7,    -7,    -3,   -17,     7,    -5,    -4,    -7,   -28,    16,     3,     6,   -20,   -12,    -7,    -3,     1,     2,    -1,    -6,   -11,     4,    -3,   -22,    -6,     0,    -2,    -6,    -5,     1,   -16,    -2,    13,    11,   -25,   -13,   -32,    -2,    20,    14,   -24,   -16,    -6,     1,    -4,     3,   -12,     4,    -5,    -5,    -8,     0,     2,    -7,     1,   -13,     1,     4,   -33,    -2,   -12,   -22,     5,    -5,   -26,   -31,    -7,     5,   -14,    -3,    -4,    -3,     3,    -2,     1,    -5,    -2,    -6,    -6,     0,    -3,    11,    12,     8,    14,     6,   -52,   -35,   -14,   -18,   -26,    -6,   -32,   -38,   -33,   -13,    -9,    -1,     1,     3,     4,     3,    -4,    -4,    -2,     1,   -10,   -14,   -17,    -6,   -14,   -12,    -6,     2,    -1,    -4,   -20,   -26,    -6,   -14,   -10,   -22,   -18,     0,     0,    -4,    -4,     1),
		    25 => (   -4,     3,     2,    -4,     1,     0,     2,     4,     0,    -4,    -2,     1,     1,    -5,    -4,     1,    -1,     5,    -1,     1,     4,    -4,    -3,    -2,     4,    -4,    -2,     1,     2,    -3,     5,     5,    -2,     5,    -2,    -1,     1,     3,    -5,   -10,    -4,    -8,    -3,   -10,   -13,   -17,   -15,    -8,     0,    -1,     0,    -2,     3,     1,     5,     2,    -4,     2,     1,    -4,     1,    -1,     1,     0,    -8,     1,   -11,   -12,    -9,    -5,   -15,    -2,   -12,    21,    17,   -18,     7,    -2,    -6,    -5,    -7,   -14,    -3,     2,     1,    -3,    -4,     6,    11,   -15,    -8,   -11,    -5,    -5,    -7,   -15,   -20,   -33,    -9,     7,     5,    15,    18,   -12,     9,    18,     7,   -18,   -15,    -7,    16,     2,     3,    -2,    -7,     9,    -6,     2,    -3,    -4,    -6,    -3,   -15,   -46,   -33,   -36,    -1,    15,   -14,    10,    16,     0,   -11,    -2,   -11,     9,    10,     9,     2,   -28,     0,     1,   -11,     2,    -5,    -2,    -7,    -6,    -7,   -16,   -36,   -42,   -20,   -16,   -13,    -7,     2,    -6,   -10,    -1,     1,   -19,    -8,    19,     8,    29,    -7,   -15,     1,     3,     3,    -5,    -7,   -15,     2,   -12,    -8,   -15,   -21,   -58,    -7,    -9,    20,     2,    -3,   -15,     1,    18,     8,    -5,    23,    20,    24,    23,    -2,    -1,    -1,    -1,     2,   -10,    -8,    -6,     6,     0,   -13,   -44,    -8,   -42,   -18,    -5,    -3,     6,    10,     4,   -11,     0,    -6,    10,    20,    22,    15,    36,     7,     3,    -5,   -15,   -18,    -8,    -3,    -5,    11,   -13,   -17,   -12,    -4,     2,    23,    -4,    -6,    -3,   -13,   -11,     5,     4,   -12,    11,    22,    33,    30,    32,     1,    16,    -4,     0,   -20,   -12,    -3,     8,   -13,   -13,     0,    -4,    12,    -7,    10,   -17,     1,    -4,   -13,     4,    -5,    -9,    -4,    -3,    21,    32,    54,    32,     0,    23,     0,    -7,    -3,    -1,    -9,    -2,     1,    -1,    -8,   -28,    14,   -10,     9,    11,    25,    -1,    -9,   -15,    11,    13,    15,   -17,     6,     9,    32,    22,    19,    20,    -4,     2,    -7,    -4,    -2,    -1,     7,    -3,    -2,    -6,    14,    -3,    -1,    -5,   -14,   -14,   -35,   -30,   -26,     6,   -35,   -17,    -4,     5,    -6,     8,    27,     7,     3,     3,     2,    -4,   -11,    -3,     7,     5,    14,     1,     6,    -6,     5,    16,   -11,   -35,   -65,   -70,   -64,   -70,   -64,   -65,   -42,   -20,   -21,    -1,    16,   -26,    -3,    -6,     2,     0,   -13,    -3,    15,    12,    -6,     4,     9,   -13,     7,     3,     3,   -27,   -40,   -51,   -68,   -54,   -58,   -57,   -58,   -34,     2,     0,    23,   -13,     7,     1,    -9,     1,    -7,   -11,    -4,     2,    -3,   -10,    13,   -14,    -3,    -1,    -9,   -11,   -25,   -53,   -64,   -52,   -45,   -38,   -30,   -25,     4,     5,     0,   -14,     2,    -7,   -11,     0,   -10,   -28,   -23,   -26,    -2,    -6,    -5,    -5,    18,   -10,     5,     7,    -4,    -1,   -28,   -42,   -49,   -37,   -29,   -15,    -9,     0,    -4,    -7,     5,    -7,   -11,    14,   -10,   -22,   -37,   -41,   -17,   -19,   -11,    -6,    -1,     3,     9,     0,     8,     4,   -23,   -36,   -51,   -35,   -26,   -23,    -7,    -8,   -14,    -5,     3,    -3,   -26,    31,     9,   -22,   -38,   -40,   -18,   -28,   -33,    -6,    12,    -3,     4,    -3,    13,    22,   -23,   -30,   -41,   -26,   -18,   -27,   -22,    -9,   -17,   -16,    -1,    -5,     1,    35,    26,    15,     0,    -4,   -27,   -31,   -25,   -24,   -14,     5,    -6,    -9,   -12,   -12,   -22,   -14,   -42,   -21,   -14,   -17,    -7,    -7,   -18,    -6,     1,    -3,     6,     4,    24,    19,    25,    31,    -5,   -22,     1,   -18,   -20,    12,   -17,     0,    -1,    20,   -22,   -15,   -19,   -10,   -11,   -16,    -5,   -26,   -13,   -11,    -5,    -3,     2,     4,    -8,    17,    18,    34,    16,     3,    -3,     3,     6,    13,     3,     6,    21,    -2,    -9,   -25,   -17,   -10,    -6,    -1,    -3,     0,    -8,    -2,     1,    -3,    -1,    -6,   -17,   -14,   -19,    16,    19,     9,    -3,    11,    10,     4,    19,    11,     6,    -9,    -4,   -14,   -15,    -5,    -6,    -7,     0,     1,    -6,     1,     0,     4,   -11,    16,    -3,   -18,     2,     9,     1,    -1,     1,    23,    15,    -3,     2,     5,   -17,     1,    -3,   -14,   -18,     1,     1,    -3,     2,    -9,    -2,    -4,    -2,    -2,    14,    11,    13,    -7,    -1,    29,    26,    24,    11,    27,    16,     5,    10,     0,    -1,    17,     2,    -2,    -8,     0,    -1,    -3,     4,    -6,   -19,     0,    -2,     1,    -9,    -5,     0,   -17,     5,    19,     3,    32,    22,    20,    19,     9,     2,   -11,   -15,     9,   -10,     5,    -2,    -3,     1,    -2,    -2,   -27,   -10,     4,    -3,     2,     3,    -1,   -22,   -21,    -3,   -17,   -11,    15,    -4,   -10,   -10,    -2,   -27,   -23,   -15,   -11,    18,     9,     0,    -9,    -5,    -3,     3,     0,    -1,    -1,    -3,    -2,     0,    -3,   -11,   -11,   -36,   -35,   -15,    -6,    10,    17,    23,    10,   -29,   -35,    -9,     0,   -10,     1,     3,     4,     5,   -13,     3,    -1,     0,     0,     3,     4,     2,    -1,    -7,     1,    -7,     0,    -4,    -2,    -1,     5,     4,    -2,    -6,     0,     1,     3,    -1,    -5,     2,    -4,   -18,     0,     1,    -5,    -5,     0),
		    26 => (    1,    -1,     4,    -2,    -3,    -4,     2,     4,    -2,    -2,     2,    -4,    19,    15,    -2,     2,    -1,    -3,     2,     2,     1,    -1,     2,     1,     3,    -2,     4,    -2,    -4,     5,    -2,     1,    -3,    -2,    13,    20,    22,    14,    43,    39,     7,    18,   -19,     4,    -8,     2,    15,    18,    52,    19,    10,    20,     5,    -1,     2,    -5,    -4,     0,     7,    13,    27,    36,    16,    24,    47,    38,    20,    22,   -37,   -23,    -1,    -3,    -2,    23,    13,    -2,    15,    16,    29,    17,     4,   -21,    -3,     2,     4,     1,   -42,    -8,    -2,    36,    31,    10,     5,     3,    -6,   -27,   -37,    -6,    17,    10,    -6,    16,    15,    11,    -2,   -12,     3,    36,    18,   -28,   -22,     3,    -1,     3,   -38,    -1,     0,    29,    -3,    -8,    20,    27,    -9,   -21,   -59,   -15,     2,   -17,     8,    -6,   -20,     2,    -9,    16,    18,    34,    -3,   -39,    22,    35,     5,    -3,   -31,   -25,    11,   -14,   -37,    20,    13,     5,   -24,   -52,   -20,   -12,     1,     0,   -30,    -5,   -29,   -17,    -2,     1,     6,    23,     5,   -20,    47,    31,     0,    -4,    13,    -8,     6,   -13,   -24,    13,   -10,   -36,   -22,   -26,     4,   -27,   -26,    -3,   -11,    -8,    -4,     5,    -8,   -17,    20,     1,    11,   -15,    13,    19,     0,     1,     1,   -15,     8,    -5,   -13,    -6,   -17,   -27,   -26,    -4,    -6,   -13,    -9,   -15,    -4,    -8,   -22,    -7,    -9,    -4,    -1,     4,     5,    -2,     8,    15,    -4,     5,   -20,   -17,    11,   -16,   -24,   -23,   -17,   -31,    -3,    -9,   -17,   -12,   -22,   -22,   -15,   -20,   -42,    -1,   -37,    -1,    -9,    -8,    12,   -50,   -10,   -34,     4,     0,   -24,     8,     5,   -38,   -11,   -28,   -25,     1,    -4,     5,   -17,   -13,    -6,   -34,   -53,   -47,   -50,   -28,   -30,   -28,   -74,   -25,     6,    -2,   -12,   -36,    -3,    -3,   -30,   -25,   -15,   -29,   -40,   -41,   -25,    10,   -16,    -6,     4,    -2,   -18,   -22,   -37,   -29,   -18,   -13,   -14,   -14,   -23,    18,    22,    35,   -20,   -44,     3,    -2,     2,   -18,   -11,   -13,   -22,    -2,    -5,     6,    15,    10,     6,    25,     7,    -8,    -4,   -13,   -27,   -35,     8,   -20,   -17,     5,     6,    -9,   -24,   -11,     2,    -1,    -5,   -19,   -15,   -29,     0,    12,    23,    33,    31,    10,     3,     6,    -3,    -6,     9,    -5,   -22,   -49,   -37,    -9,    17,    35,    24,    -3,   -41,    -8,     4,     1,    -9,   -16,   -17,    -2,    30,    15,     6,    22,    31,     8,     3,   -12,    -7,     0,    -2,     2,   -18,   -15,   -25,   -14,    10,    35,    23,    11,   -13,     4,     0,     4,    -5,   -32,   -26,    21,    10,    11,    24,    33,    10,    20,    -2,   -19,    -3,    -3,     8,    -7,    -8,    -6,    -7,    14,    27,    22,     7,    11,   -31,   -22,     2,     1,   -12,   -36,   -31,    25,    27,    30,    44,    41,    25,    19,    19,     5,    -9,   -18,    -5,     0,    -3,     8,     4,    -8,    27,    23,   -27,   -13,   -41,   -21,     2,    -2,    -1,   -30,    -5,    19,    16,    33,    53,    47,    35,    32,    31,     2,     5,    -3,    12,    -7,    -9,    24,    14,     6,    20,    27,   -16,   -27,   -38,   -23,    -4,    -5,    -2,   -29,   -29,    12,    13,    22,    18,    18,    38,    13,    32,    41,     3,    -2,    -6,   -11,    -6,    10,     9,    20,    -2,    -5,   -10,   -29,   -45,   -35,     4,    -1,    -5,    -3,   -17,   -12,    -4,    17,   -10,    12,    11,     1,    28,    40,    12,   -24,     1,    -1,   -14,   -23,    -2,    -6,   -11,   -17,   -48,   -33,   -24,   -24,     2,    -2,   -25,     2,     0,   -34,   -23,    -7,   -21,     1,    -6,    15,    13,     5,    -1,    -7,   -10,    13,   -13,   -11,    -9,    -2,    -4,    -4,   -22,     6,   -18,   -29,     4,    -7,    -2,   -34,     7,   -26,   -22,   -19,   -15,     5,    -6,    -3,    -6,   -19,    16,    -4,   -22,   -14,    -2,   -10,    -5,   -10,    22,     0,    17,    33,    -7,     1,    -4,     0,   -12,   -16,   -16,   -12,   -22,    -7,    -5,     7,     4,   -21,    27,    27,     3,   -17,    -4,     1,     4,    16,    -4,    -2,    21,    24,    22,    10,    -4,    -9,     2,    -3,     0,   -12,   -17,   -44,   -45,   -28,    13,   -16,     2,   -13,    21,    26,     8,    12,    20,     3,     5,    10,    -8,    17,    -8,    -1,   -15,   -36,    -5,    -6,     5,     0,     4,    -5,   -20,   -35,   -41,   -31,   -18,   -10,   -11,     2,   -14,     3,    -4,     9,   -14,     0,    20,    27,     1,   -23,   -38,   -30,   -28,   -27,   -42,     2,     5,     2,    -1,    -1,   -12,   -11,    -5,   -27,   -28,   -41,   -46,   -32,   -11,   -21,     3,    13,    18,    20,     5,   -49,   -21,   -49,   -29,   -23,   -15,   -18,     2,     0,     3,    -1,     0,    -4,     1,    -8,    -7,   -25,   -13,   -15,   -23,    -1,    23,    -1,   -19,    -8,   -22,   -19,    -7,   -18,   -36,   -11,   -14,   -12,   -10,    -2,    -1,    -3,     4,     0,     2,    -4,    -1,    -8,   -12,    -5,    -2,    -6,   -15,   -12,    -3,    -5,     0,    -6,    -3,     1,    -2,    -5,    -6,    -8,    -5,    -3,    -5,     2,    -1,     4,    -5,    -1,    -4,     5,    -4,    -4,     4,     1,    -3,    -2,     0,     1,     4,    -1,    -4,    -1,     0,    -5,     0,    -5,    -1,    -7,    -2,    -2,    -1,    -5,     1,     0),
		    27 => (    5,     1,     5,     1,     3,     3,    -2,     4,     2,    -2,    -3,     4,    -3,    -4,    -1,    -2,     1,    -5,    -4,     0,    -4,     4,     1,     0,     1,     1,    -3,     0,    -4,     2,    -1,    -5,    -4,    -4,    -2,     4,     5,    -2,    -1,   -22,   -16,   -19,    -1,    -4,    -7,    -5,     3,    -2,    -2,    -5,    -5,    -4,    -1,    -2,    -3,    -4,    -4,     3,     5,    -6,    -8,     1,     0,    -7,    -5,    -3,    -6,   -13,   -22,   -14,    -5,    -4,    -2,     3,    -2,    -5,     0,    -2,    -7,    -1,     2,    -4,     0,     3,     5,    -5,    -1,   -10,   -10,    -8,    -8,   -12,   -19,   -18,   -13,   -26,   -18,    -9,    -4,    -7,   -13,   -12,    -2,   -13,     0,   -17,   -13,    -8,    -4,     1,     4,     2,    -4,     4,     1,    -1,   -26,     0,    -7,   -25,   -23,   -32,   -43,   -41,   -36,   -43,   -32,   -35,   -26,   -12,   -10,    -6,    -1,   -18,   -28,   -21,   -17,   -13,    -8,     3,    -1,     4,     2,   -15,     5,     7,    -6,   -25,    19,    16,   -22,   -17,   -29,   -25,   -22,   -30,   -39,   -80,   -97,   -64,   -45,   -17,    -2,   -44,   -33,   -32,   -16,    -1,    -2,     2,     5,    43,    34,    27,   -12,   -25,    27,    -3,   -16,    -3,    13,    17,     1,   -30,    -5,     4,    17,    -3,    11,    39,    -1,   -55,   -41,   -39,   -27,    -1,    -3,    31,     0,    33,    32,   -10,     1,     2,     3,    14,    25,    21,    14,     0,    -4,    -6,     8,     9,     3,    23,    16,    21,    32,    35,    -2,   -16,   -31,   -16,   -24,    38,     9,    25,    13,   -21,   -18,     6,    14,     4,     3,     9,     6,     8,    -2,     7,    11,    -4,     7,    10,     7,    16,    12,     6,    12,   -22,   -43,   -10,    -2,    24,   -12,     4,    14,    11,    -1,    18,    19,    25,    24,    16,    25,     1,    -7,    -3,    -7,     4,    -1,    20,     8,    35,     7,    -1,    -4,    -9,   -39,     0,     1,    14,    -1,   -16,    26,    20,     4,     9,    12,    11,     4,    27,     5,    -9,   -34,   -18,     2,    27,    -5,    15,    19,    10,     8,   -10,   -20,   -24,   -25,     6,     1,   -11,    30,    -5,    25,     8,     9,    19,     1,     4,    33,    42,    -5,   -51,   -76,   -13,     8,    14,    -5,    -3,    18,    -8,    -5,    -9,     6,   -36,    -9,     3,     0,    17,     4,     3,     2,    21,   -16,    12,     3,     0,    20,    -5,   -45,  -114,   -75,    -8,    10,    -2,     7,   -34,    -2,     6,    -4,   -42,    -2,   -13,   -11,     5,    -3,    19,     2,    -4,   -17,    -5,     7,    15,    19,    15,    12,    -1,   -71,  -122,   -45,   -14,     4,     0,   -24,   -33,     2,     5,   -33,   -40,   -14,   -10,   -13,    -7,     0,     4,    18,     3,    -5,   -11,    21,    11,     9,    10,    25,   -37,  -102,  -104,    -2,    -4,     6,    -6,   -28,    -5,     0,   -16,   -16,     2,    16,   -10,    -7,    -2,     0,    -4,    17,    -4,   -16,     5,    -1,    19,    -1,    -6,     1,   -67,  -113,   -26,   -13,   -23,    -4,   -10,    -7,    -4,     8,    -8,    -3,     7,    17,    -3,     0,    -4,     5,     1,    15,   -15,   -19,     1,   -11,    -1,    -5,   -26,   -31,   -66,   -38,   -13,   -18,   -12,   -18,    -8,   -14,    -8,     4,    -3,   -10,   -31,   -35,   -16,    -2,   -10,     3,     1,    -1,   -12,   -17,   -12,   -44,   -24,   -18,   -18,   -13,   -10,   -35,   -28,   -16,   -10,     3,     1,    17,     7,    -3,     5,     0,   -32,   -42,   -19,     0,   -21,     5,    -4,    25,   -28,   -33,    -6,   -18,   -21,   -22,    -4,    -6,   -25,   -31,   -19,    -4,   -20,     3,    10,    11,     7,    -2,   -27,   -13,   -22,   -48,   -38,     0,   -13,     5,    12,     2,   -32,     5,    16,    -6,   -37,    19,    19,   -11,    -1,   -13,    -8,     7,    -9,    -7,   -17,   -17,    -5,    -3,   -22,     7,   -22,   -24,   -13,    -4,    -4,     1,    24,    -6,    -9,   -13,   -36,   -29,    -8,    -2,     5,     3,    -9,    23,   -11,    -4,    -4,   -24,   -16,   -20,    -1,   -21,   -51,   -38,   -38,   -31,    -3,   -11,     4,    -1,     4,    -3,   -19,   -34,   -28,   -26,   -40,    -9,   -17,     5,    21,     8,    -2,     3,    -8,    -8,   -21,    -8,     3,    -4,    11,     9,   -18,     2,    -2,   -13,    -1,     1,     2,    -6,   -16,   -23,     7,   -26,   -18,    -6,     3,    -2,   -11,   -10,     5,    -6,     5,   -13,   -11,     8,     8,   -19,    -8,   -13,   -18,    -8,     2,   -40,     2,     1,     3,    -7,   -19,     6,    24,    10,     4,   -16,    10,    17,   -13,   -27,     4,   -13,     1,     2,     2,   -12,    -3,   -21,     2,   -26,   -15,    -7,    -3,   -22,    -2,     1,    -3,    13,    27,    56,    33,    -4,   -10,     2,   -15,    20,   -11,    -8,   -31,   -39,     6,    -9,    -6,   -12,    -3,   -18,     4,   -13,    -8,    -2,   -10,    -1,     2,     3,     4,   -25,    19,     4,   -30,   -22,    -4,     8,    -1,   -26,   -11,    21,    -4,    17,     8,    -1,     5,     2,    -8,     5,    34,    17,   -18,    -5,     1,     3,     0,    -1,     0,    -5,   -15,   -25,   -35,   -15,    21,    28,    -6,   -27,   -22,   -17,     8,     0,    16,     8,   -11,     0,    24,    16,    -5,    -2,    -6,    -9,    -5,    -2,    -5,     0,    -4,     2,    -1,    21,    25,     9,     2,    13,    13,     9,     2,     3,    25,    25,    -5,     0,    25,     7,    19,    15,     5,     4,    30,    -5,    -3,    -4,     2),
		    28 => (   -1,    -4,    -3,    -1,     1,     5,    -4,    -1,     0,    -2,     5,    -3,    -4,    -5,     0,    -3,     4,     3,    -4,    -1,    -2,     4,     0,     0,     0,     0,    -1,     3,     1,    -4,     2,     4,     1,     5,     2,     0,     4,    -5,    -5,   -17,   -18,   -21,   -21,   -39,   -30,   -39,    -6,    -9,    -3,     7,     2,     2,     3,     0,     1,    -5,     4,     0,    -1,    -4,    -6,    -3,   -10,    -1,   -14,   -34,   -55,   -51,   -25,   -19,    -8,   -45,   -46,   -40,   -18,   -32,   -19,   -22,   -27,   -21,    -8,    -9,     4,     1,     3,    -5,   -17,   -13,    -8,   -34,   -56,   -69,   -81,   -89,   -55,   -50,   -12,    25,   -14,    -2,   -14,   -28,   -56,   -54,   -14,     9,    19,    24,    16,    -1,   -11,    -2,    -2,   -19,   -11,   -34,   -41,   -66,   -31,   -29,    -9,   -13,    -2,   -23,   -22,    12,    11,     0,    -6,   -15,   -21,     9,    18,   -20,   -16,   -16,    13,   -21,    24,    -3,     3,    -2,   -29,   -25,   -22,   -56,     0,    -3,     6,    -1,   -19,    -3,    -9,     0,    13,   -14,    -6,    -4,   -30,    -5,    -5,    21,    15,    -8,    37,    31,   -25,     6,    -1,    -1,   -10,   -46,   -17,   -23,    15,     1,    -1,    -3,    -5,     8,     8,   -15,   -14,    -6,     6,    -4,    14,   -13,    10,    17,    19,    27,     9,   -20,   -22,     2,    -4,   -17,   -10,   -40,     3,    10,    -4,    15,     4,    -4,    13,    -3,    -9,   -14,   -24,     3,     3,     0,     5,     0,   -21,    18,    33,    11,   -10,   -17,   -31,     5,   -16,   -21,   -35,    -3,    -4,   -10,     9,    11,    -3,    17,    -4,   -19,   -11,     6,   -13,   -35,   -23,     6,    16,     2,     0,    -4,    22,    13,    25,   -20,    17,    15,    -3,   -15,   -38,    -4,   -30,    -6,    -6,   -12,    17,    -4,   -11,   -10,   -15,    -7,   -22,   -29,   -12,    10,   -26,    19,    -9,   -12,    -6,    21,    28,    -1,    13,   -15,    -4,    -5,   -51,   -46,     9,    -5,    -9,    14,    -2,    16,   -11,    -4,    -6,   -16,    34,     6,    -9,   -14,    -7,     7,     4,     1,     4,    41,    23,   -24,     8,    -7,     1,    -4,   -31,    33,    11,     9,    -6,    -3,    11,    -3,     4,    -2,     8,    17,    32,    36,     3,    -3,    -7,    -6,    11,    10,    -3,    13,    50,    50,    26,   -21,     1,    -2,   -22,    37,    22,    17,   -12,     3,    -2,   -22,   -23,    22,    35,    36,    19,    23,    11,    29,    -9,    30,     8,     0,   -31,    -6,    13,    34,    16,   -23,    -1,     1,   -14,    44,     3,     5,    -8,    11,   -15,     2,     7,    33,    21,    33,    29,    27,    17,    15,    18,    25,    -9,   -33,     5,   -16,   -31,    -4,   -12,     2,    -3,    -4,    -6,    32,    10,     5,     9,   -15,   -24,    -4,    41,    24,    18,    33,    16,     2,    16,    13,    15,    11,   -31,   -40,   -23,   -17,   -27,    32,   -32,     1,    -2,    -2,   -12,     0,   -44,   -30,   -11,    10,     5,    26,    28,    21,    18,    32,    22,    11,    20,    14,    -4,   -17,   -22,   -33,     6,     9,   -36,    36,   -72,   -24,    -5,    -5,    -6,    -6,   -10,    -8,     7,     5,    10,    13,    40,    11,    35,    -3,     9,     6,    33,   -21,   -14,     3,   -27,   -14,    -6,    32,   -40,    16,   -59,   -27,    -3,    -3,    -7,   -26,    26,    11,    41,    -7,   -16,    17,    29,    39,    34,    38,    28,     0,    35,     1,   -24,   -11,   -18,   -11,     7,    50,    16,   -30,   -15,   -36,    -5,    -6,   -11,   -32,    30,    -3,    -9,     6,    -7,     4,    18,    25,    49,    59,    27,    22,    -6,   -16,   -12,   -29,    -9,   -16,   -10,    11,    -7,   -35,   -19,   -14,    -4,    -4,   -37,   -15,   -16,    -2,    13,    -8,    13,     7,     7,   -19,     4,    28,     8,   -16,   -36,   -21,    -1,    -9,     5,    -9,    12,   -16,    -7,   -42,   -56,   -13,    -1,    -1,   -15,    -1,    -4,     3,    14,     5,   -28,    -7,   -13,   -22,   -16,   -16,    -7,   -14,   -10,   -21,     1,    -8,    12,   -14,    19,   -22,   -17,   -32,   -33,     1,   -17,    -3,   -23,     5,   -10,     4,    -3,   -15,   -25,     0,   -28,   -39,   -32,   -22,   -18,   -25,   -25,    20,    22,   -11,     2,    -6,    -4,   -22,   -51,   -31,   -56,    -9,   -10,    -8,   -13,    -3,     8,   -23,    -9,     2,     4,    -5,   -12,   -25,   -17,   -29,   -22,    -6,   -19,   -28,    -8,   -11,    -5,    21,   -20,   -28,   -40,     7,   -25,    -3,    -2,    -1,   -17,     8,     2,     0,   -30,    -2,     7,    14,   -20,   -17,   -19,    -4,   -24,    -3,    -3,     1,     1,    17,    29,   -18,     8,    18,   -19,     8,   -33,    -2,     4,     4,   -15,   -12,   -55,   -42,   -36,   -50,   -29,    -2,    -1,    -8,    -1,    -6,   -21,   -13,   -27,   -35,   -18,    24,    -9,   -32,   -12,     6,   -13,   -19,    -9,    -5,     1,    -2,   -17,   -13,   -12,    -3,    23,    18,    -9,    -3,    33,     5,   -31,   -16,    -2,    12,    19,     0,    10,   -23,   -13,   -22,   -32,   -22,   -34,   -23,   -14,    -2,    -1,     2,     3,   -14,   -15,   -31,   -40,   -39,   -48,   -70,   -55,   -28,   -24,   -24,   -27,   -69,   -36,   -23,   -29,   -55,   -41,   -25,   -15,   -15,    -1,    -4,    -1,    -5,    -1,     2,     2,    -2,     0,    -5,    -4,   -17,   -30,   -33,   -20,    -5,   -10,   -25,   -30,   -36,   -22,   -24,   -15,   -19,     2,    -4,    -2,     1,     0,    -1,     3,    -3),
		    29 => (    4,     0,     2,    -5,    -1,     0,    -4,     4,     0,     4,    -5,     1,     4,     3,    -4,     4,    -1,    -2,    -2,    -3,    -2,    -4,    -1,     3,    -1,     0,    -1,    -5,     0,     1,     5,     0,    -3,     2,     1,     2,     3,    -4,    -1,    -8,   -12,    -8,     1,    -5,   -16,   -21,   -17,   -10,     4,    -8,    -1,    -2,     3,    -3,     2,    -5,     1,     3,    -3,    -6,    -8,     1,    -1,   -10,    -4,    -8,    -9,   -17,    -1,    -1,   -30,   -22,   -18,    -5,    -5,    -4,   -37,   -13,   -24,   -14,    -6,    -3,     0,     3,    -1,     2,     2,    -6,   -13,   -31,   -29,   -26,   -34,   -33,   -60,   -60,   -40,   -46,   -87,   -34,   -43,   -63,   -47,   -32,   -50,   -54,   -36,   -20,   -14,    -6,    -3,     2,     3,    -3,   -14,   -14,   -16,   -52,   -73,   -27,   -33,   -40,   -19,   -12,    -8,    -6,   -15,     7,    -8,   -30,   -10,   -73,   -63,   -19,   -27,   -15,   -11,   -36,   -24,    -4,     1,    -4,    -2,    -7,    -5,   -20,   -25,   -24,   -13,     4,     5,    20,     4,    15,    10,    -5,     5,    12,    23,    24,     8,   -32,   -33,   -31,   -11,   -25,   -17,     3,    -4,     3,    -4,   -21,   -19,   -35,   -13,   -25,     0,    22,    10,   -12,   -22,     4,     6,    13,     8,    -2,    30,    19,    23,    -7,   -11,    13,     4,    -8,   -17,   -30,    -2,    -5,   -23,   -17,   -24,   -28,   -34,   -29,    -1,     8,     5,   -11,     0,   -18,    -3,   -12,    -8,    -2,     0,     8,   -11,   -20,   -23,    -6,     5,    14,   -20,   -11,   -16,   -19,    -9,    -8,    -8,   -25,     7,    -5,    10,    24,    15,    -6,    -6,    -4,   -11,    -6,    -4,    -9,     3,   -13,   -33,   -27,   -30,   -18,     9,    -3,   -23,    -8,    -3,   -18,    10,    28,    29,    12,    13,     0,    11,    27,    -3,    -4,    -8,   -13,   -14,   -15,     7,    20,    19,    -9,    -5,   -10,   -27,   -41,   -23,   -33,   -53,   -20,     2,   -25,   -21,    16,    60,    33,    36,    22,     5,     6,    -8,   -10,     8,   -10,   -11,     9,    44,    35,     4,   -12,   -13,    -9,   -18,   -14,   -16,     8,   -16,    -9,     3,   -48,    -4,     1,    33,    34,    32,     5,   -17,    -4,    -5,     5,    -6,    14,    22,    13,    49,    34,     3,   -25,   -13,    -4,    12,    10,     4,    27,    -6,   -14,     3,   -12,     7,   -11,    24,    20,    27,    -7,    -3,    -6,    -9,    -3,    -2,    10,    50,    35,    21,     4,     8,    -8,     9,    -3,     6,     9,   -13,   -17,   -19,   -13,    -2,   -14,    -8,   -13,    18,    28,    -5,     1,   -12,   -14,    -6,     4,     2,    37,    46,    49,    22,     6,    10,   -11,     1,     8,    12,     6,    -2,    -7,   -15,    -7,     1,   -16,   -20,   -15,     3,     4,    18,     3,     4,     6,    -6,     5,    18,    45,    52,    36,    34,    11,    14,    15,    12,    -1,   -12,   -21,   -15,   -15,     2,     2,     4,     4,   -34,   -13,    -7,    -8,    11,    -5,   -19,    -9,    -8,    -1,    15,    48,    48,    28,    29,     9,    28,    15,    24,     9,   -15,   -32,   -33,   -14,    -3,    -9,     3,    -7,   -32,   -27,    -8,   -16,    20,     7,    14,   -13,    16,    11,    22,    23,    41,    29,     3,    14,    28,    25,    37,     2,    -9,   -18,   -43,   -31,    -8,   -12,    -3,     0,   -30,    -5,   -13,   -27,    21,    26,    -5,     9,     3,    34,    24,    16,    38,    14,     6,    15,    22,    15,    25,    -1,    -7,   -18,   -41,   -16,   -25,    -9,    13,    -3,   -31,   -13,   -31,   -33,    25,    30,    28,    19,    13,     5,    -2,     7,     6,     9,     3,    39,    16,    26,    18,   -11,    -2,   -26,   -48,   -23,   -25,   -24,     0,    -1,   -42,   -10,   -37,   -33,    15,    30,    20,    23,    13,     7,    -7,     2,   -18,     3,    33,    24,    14,     2,     1,     1,    10,    -4,   -13,    -8,   -12,   -10,     1,    -5,   -38,   -15,   -37,   -23,   -17,     6,    22,     5,   -10,     2,    10,   -10,   -18,    -6,    15,     8,    -1,     1,    -5,   -11,   -10,     0,    -4,    13,   -13,     3,     1,     2,   -35,   -15,   -30,    -2,   -13,     3,   -20,    -7,   -14,     3,     8,   -16,   -18,    15,     2,     1,   -21,   -15,    -8,   -10,   -18,    -7,     8,    -1,   -32,     0,    -3,     0,   -25,    19,   -20,   -30,    -9,   -15,   -15,    -6,    -6,     3,     4,   -26,    -7,     4,   -23,   -26,   -29,   -15,   -13,   -29,   -20,   -16,     6,   -22,    -9,    -2,     0,     3,   -17,     6,   -13,   -19,    -4,   -24,   -28,   -25,   -24,    -2,     7,    -3,     3,   -15,   -29,   -22,   -21,   -18,    19,   -19,   -21,   -29,     4,    -6,   -17,    -3,    -4,     3,   -22,   -30,    -9,     7,   -25,   -23,   -10,   -11,   -10,    -9,     3,     0,   -13,   -35,   -28,   -18,   -23,   -21,   -13,   -12,     0,   -12,     1,    -3,    -2,    -3,    -2,     3,    17,   -11,    -5,    -8,   -27,   -40,   -23,     1,   -15,   -13,     0,    -9,   -10,   -34,     3,    -9,    -7,   -21,   -13,   -12,    -1,    18,    -9,     1,    -6,     1,    -4,    -3,    -1,    29,   -13,   -29,   -21,   -24,   -19,   -15,   -18,     0,     4,    -2,     0,    -8,    23,    15,    12,   -27,    -2,     5,    -4,     4,     5,     4,     4,    -3,     5,    -2,    -3,    -3,    -3,    -8,    13,    17,     8,    11,     7,     3,     1,    20,     8,    -6,    -4,   -17,     0,     1,    -8,   -17,    -7,   -17,     0,    -1,     0,    -2),
		    30 => (    4,    -4,    -2,    -1,    -3,    -2,     4,     2,     0,     1,     0,    -4,     2,    -1,    -9,     0,     0,    -1,    -3,    -2,    -5,    -1,    -4,     2,     1,     5,    -5,     4,    -5,    -3,     0,     0,     4,    -1,    -3,   -22,   -19,   -32,   -20,    16,     7,     5,   -13,    20,    28,    21,   -12,    -6,    -4,    -6,    -6,    -3,    -1,     1,    -2,     1,     0,    -1,     3,    29,    26,     1,    -4,    -3,   -19,   -25,   -38,   -48,   -27,   -41,   -36,   -61,   -52,   -57,   -37,   -31,   -28,   -24,   -34,   -20,   -11,   -11,     0,    -3,     2,     3,     1,    18,    -9,   -18,   -17,   -29,   -27,    -9,   -32,     5,    17,    22,   -12,   -41,   -14,   -10,   -37,   -50,   -12,   -22,   -20,   -22,   -29,    -4,   -15,    -1,     4,    -2,   -16,   -34,    -8,   -42,     5,     1,    -5,     3,    10,    -4,     6,     5,   -16,   -18,   -35,    -1,     0,    15,     2,    -1,   -12,   -22,   -41,   -48,   -20,    -3,    -5,    -2,    -8,   -25,    -5,    -9,    16,    10,    -1,   -13,     9,    -8,   -26,   -27,   -10,   -18,   -23,    -5,    11,    12,   -18,   -17,     3,   -29,    -3,   -61,   -37,    -4,    -3,     1,    -6,    -2,    -6,     0,     2,    16,     9,   -43,    -1,   -15,   -30,     4,   -10,    -6,   -10,    -2,     0,     4,   -11,     1,     9,    -1,    13,   -51,   -15,    -2,     4,   -11,    -1,   -16,    -4,    -5,     0,     0,   -22,     1,    -5,    25,    -8,    19,    -2,   -14,     6,    -1,    14,    21,     7,    25,    14,    34,     7,    -1,   -32,     0,    42,   -32,    21,     6,   -13,   -34,   -27,   -13,    -6,    -1,    23,     0,     8,    -4,     3,    28,    26,    31,     7,    25,    26,    25,    25,     2,     3,   -26,   -46,   -15,    -4,    -2,    34,   -25,   -23,   -16,   -19,   -23,    -2,    11,     7,     1,    -1,    -3,    15,    12,    17,    12,   -13,     4,    33,    15,    -4,     1,     8,   -38,   -20,    -6,    -9,    -6,    30,    15,   -30,   -16,    12,    -1,    -4,    -4,     4,    -9,   -12,    -7,     1,    22,    10,    24,     3,    -1,    12,    14,     5,   -20,   -17,   -39,   -50,    -3,    -3,    34,   -26,    -7,   -56,     1,     9,     7,     9,   -16,   -11,   -24,   -22,     4,   -12,   -18,   -11,    -9,   -13,   -15,     2,    28,     6,   -32,   -42,   -39,   -32,    -4,    -1,     6,   -23,    -6,   -11,     6,    19,    14,    -2,     8,    -5,   -31,   -12,    -6,   -31,   -18,    -6,   -12,   -14,   -10,    -1,    19,    23,     0,   -22,   -10,   -18,   -13,    -3,     8,     0,    17,    25,     9,    36,    20,     1,    16,     0,   -18,    -7,   -27,   -12,   -30,    -8,    14,     4,     9,   -27,    11,     1,    -2,   -24,   -11,   -22,   -21,     3,     0,    -2,    -5,    43,    48,    49,    23,    17,    23,    26,     9,     0,   -20,   -24,    -3,   -24,    -2,     2,    13,   -10,   -33,    -1,   -14,    12,   -31,   -43,     0,     1,     0,   -20,   -16,    31,    55,    15,    32,    36,    53,    32,   -10,    26,   -18,   -18,   -10,   -15,     1,    -3,   -11,    -4,   -23,     3,     7,    -2,   -24,   -47,   -23,    -3,    -1,   -12,   -38,    33,    35,    22,    22,    43,    47,    18,    37,    27,   -16,     5,    11,   -14,    -9,    -1,   -15,   -11,   -27,   -32,    18,   -34,   -52,   -66,    35,     3,    -3,   -11,   -48,    13,    14,    -9,    20,    11,    21,    29,    31,     1,   -15,    -7,    -5,    -3,     2,     2,     1,     1,   -32,     9,   -10,   -35,   -39,   -34,    50,    -4,    -4,    -8,   -53,     0,    -7,    -7,     1,    22,    10,    15,     3,    12,    -3,    -4,     2,    -9,   -17,   -14,   -13,   -14,   -13,     1,   -12,   -17,   -31,   -34,   -12,     1,    12,   -14,   -38,   -17,    -6,    -8,    -5,    -8,   -28,   -14,    -5,    22,     5,    -3,     0,   -11,   -21,    -6,     1,   -15,     1,     3,   -16,   -15,   -54,   -29,   -12,     1,    18,   -12,   -45,   -11,    -2,    -8,   -17,   -25,   -30,   -11,     8,    -5,     7,    19,    10,    -3,   -15,    -1,   -14,   -13,    -9,    -9,   -11,   -19,   -49,     0,    -4,    -4,     3,   -39,   -26,   -28,    -7,    15,     5,   -13,   -13,    -9,    -7,    10,    28,    21,    26,    24,     6,   -11,   -33,   -28,   -11,     3,   -11,   -14,   -14,    32,    11,     0,     3,   -53,   -16,   -49,   -16,     0,    10,    30,    -2,    12,    12,    42,    17,    33,    28,     3,    -3,   -15,   -18,     2,    10,    18,    19,   -22,   -14,    18,     9,     2,    -3,   -13,   -53,   -42,   -10,    11,    -7,    -1,   -12,     6,     7,    11,    11,    20,     5,    16,   -15,   -14,   -13,   -12,    13,    -8,   -18,   -22,   -16,   -39,     0,    -2,     1,    -5,   -12,    -7,    16,   -14,   -23,   -29,   -47,   -45,   -29,    12,    34,    32,    29,    26,    -4,   -12,   -47,   -33,   -15,   -24,   -28,   -16,     1,    -3,     4,     2,     4,     0,   -16,   -82,   -65,   -16,    -6,    -6,   -52,   -40,   -27,    -4,   -11,   -15,   -24,    -7,    -4,   -32,   -53,   -39,   -37,   -21,   -10,     2,    -1,     3,    -2,     1,     1,     4,    -2,   -42,   -36,   -52,   -18,   -25,   -41,   -39,   -20,   -23,   -25,   -43,   -35,   -25,   -57,   -56,   -26,   -35,   -39,   -18,   -22,    -7,    -3,     0,    -2,     1,    -5,     1,    -2,     2,     1,    -5,    -3,   -15,   -10,     3,     3,     2,   -14,     0,     1,    -9,    -9,   -13,   -13,    -6,   -18,   -19,   -17,    -2,     3,    -4,     5),
		    31 => (    3,    -4,    -2,    -2,     1,    -4,     2,     3,    -3,    -3,     2,    -4,     2,     5,    -3,     3,    -4,    -4,     4,    -1,    -1,    -5,    -4,    -4,     1,     3,     3,     5,    -2,    -1,     3,     3,     3,    -3,    -2,    -5,    -2,     0,    -7,    -7,    -6,   -19,     9,    11,     1,   -11,    -6,     3,    -2,     2,    -1,     0,     4,     5,     3,    -2,    -4,    -3,    -1,     0,    -4,     2,    -3,     4,   -15,   -24,   -16,   -16,   -32,    12,    -8,    -2,    11,     3,     7,    26,    26,   -44,   -36,   -22,    -8,    -9,     4,    -4,     1,    -1,    21,    16,     0,   -21,   -30,    15,    22,    22,    -3,   -29,   -12,   -17,     2,    21,     3,    -1,    -1,    23,    19,   -11,    -4,   -13,   -20,    -5,    -5,     1,    -2,    -3,    24,    20,    16,    25,     0,     1,    15,     5,    17,    -3,    -2,    13,    -2,    -3,     2,    26,    35,    24,    -3,    -5,     4,    -4,   -14,   -25,   -33,   -23,     3,     4,    12,     7,    26,    31,    23,    24,   -10,   -24,   -10,   -12,    -1,    -4,   -15,    -1,    -7,    -9,     2,    26,    11,    -8,    -8,    15,    -9,   -35,   -25,   -24,     2,    -4,   -21,     8,    29,    26,    29,    20,   -12,   -14,    -2,    -7,   -18,   -11,   -13,   -18,     4,     1,     5,    10,     7,   -17,   -16,     1,    -2,   -15,   -35,    -4,     1,   -12,   -34,   -13,   -47,     4,    26,    28,   -19,   -13,   -17,    -6,     2,     9,     9,     2,     3,   -23,    -3,    10,    10,    -7,    -1,    18,    -6,   -29,   -64,   -37,     1,   -32,   -36,   -46,   -44,   -19,    10,    -1,   -22,   -15,    -2,    -4,    26,    22,    27,    -4,    -6,   -10,     9,     4,   -20,   -10,    13,     3,    -6,   -26,   -89,   -18,     3,   -10,   -29,   -50,   -40,   -20,   -26,   -10,   -23,   -17,    -5,     7,    30,    31,    21,    -8,    -1,   -11,     1,     5,   -14,   -28,     1,   -10,   -22,   -26,   -40,   -22,     0,    -9,   -29,   -14,   -38,   -29,   -29,   -15,   -20,   -36,   -19,    -9,    36,    31,    18,    -3,    -6,     9,   -11,   -15,   -19,   -21,   -28,   -29,   -25,   -17,   -13,    -5,    -4,     6,    -3,   -22,   -24,   -31,   -40,   -38,   -36,   -24,   -28,   -23,     0,    27,     9,    15,   -13,    -6,   -10,   -19,     4,   -17,   -10,   -34,   -34,   -18,   -20,    26,    -1,    -4,   -42,   -13,    -6,   -26,   -24,   -51,   -35,   -29,   -15,   -15,     3,    28,    -6,     1,    20,     4,   -10,    -9,    10,   -25,   -24,   -14,   -24,    -7,     4,    23,     3,     1,   -36,    12,   -11,   -30,   -17,   -30,   -24,   -19,   -16,   -23,     1,    -4,    10,    12,    31,    22,    -2,    -9,    -9,   -45,   -36,   -34,   -33,     4,     4,    -2,    -5,    -1,     9,     4,   -17,   -21,   -25,   -16,   -24,   -14,   -25,   -22,     7,    -5,     2,     8,     7,     6,   -11,   -28,    -9,   -32,   -24,   -18,   -25,   -23,    -9,    -3,     1,     0,     6,   -17,   -33,   -27,   -28,   -32,   -22,    -4,    -5,    -3,    -1,    11,     9,     3,    13,    12,     6,   -13,   -28,   -52,   -44,   -34,   -85,   -42,   -23,   -16,    -4,     0,    10,   -36,   -32,    -3,   -12,   -22,   -13,     7,   -10,   -14,    -7,     4,     3,    -3,    12,    -1,    -6,    -7,   -20,   -36,   -20,   -15,     7,   -27,   -16,   -20,     4,     0,   -14,   -38,   -18,   -12,   -21,   -39,     7,     1,    13,    14,   -12,   -11,    24,    18,    14,     7,    -2,    -1,    -8,    12,    11,    -7,     9,   -14,   -22,   -22,    -3,     3,     3,   -44,   -28,   -28,   -59,   -39,    -1,    16,    19,    -9,   -23,   -13,     7,    29,    24,    -9,     6,   -29,   -15,    -8,    -7,     8,     9,    -2,   -20,     2,    -5,    -1,    -9,   -45,   -51,     3,     2,    -2,    15,    21,    20,    -7,   -14,     7,    12,    11,    11,   -12,   -16,   -34,   -26,     0,    19,    19,    26,    12,   -25,    -6,    -3,     2,   -17,   -46,    -9,    25,    30,    41,     8,    27,    24,     2,    13,    17,    10,     7,     7,   -17,     7,    -8,     9,    13,    25,    22,    25,     3,    -8,     0,    14,     9,    -6,    -2,    -8,    15,    22,    28,    37,    37,    17,     1,    15,    33,     1,   -14,     6,   -11,     6,    -3,    14,    18,    20,     5,     6,    11,   -16,     2,     7,     8,   -13,    -5,    -6,    23,    27,    27,    22,    36,    17,    15,    15,    31,   -31,   -21,    -4,    -8,     5,    14,    26,    19,   -19,    -8,    14,     1,     3,     1,     1,     2,    -7,    -7,   -12,     8,     8,     1,     8,    37,    22,    20,    23,    -2,   -27,   -15,   -23,     9,    -9,    -8,    12,     2,    -8,   -23,   -26,   -19,    32,    -5,     1,    -4,     5,    -6,   -20,     2,   -10,     3,    -7,    13,    11,   -26,    -7,    -3,   -30,   -28,   -28,     6,    -6,   -26,    -9,    14,    -3,   -32,   -32,     3,     5,     5,    -5,     1,     0,    -8,   -22,   -37,   -21,   -50,     4,   -21,    -5,   -22,    17,    -1,   -26,   -32,   -37,   -51,   -59,   -44,   -81,   -30,   -20,   -14,    -7,    -8,    -9,    -1,    -1,    -3,    -1,    -6,   -26,   -54,   -77,   -83,   -58,   -54,     8,     2,   -33,   -32,   -31,   -33,   -21,   -42,   -22,    -7,   -15,   -16,    -4,    -5,    -1,    -1,    -2,     3,    -4,    -1,    -1,     3,    -4,    -7,    -1,     4,     3,    -4,   -32,   -26,     3,    -8,   -23,    -9,   -10,    -2,     0,     0,     4,    -4,    -3,     4,     2,    -5,     3,     5),
		    32 => (    0,     4,     1,    -3,    -2,    -1,     1,     2,     0,    -2,    -1,    -4,   -10,    -8,     5,     0,     0,    -4,    -1,     0,    -3,     3,     4,    -1,     2,     3,     4,     2,     0,    -4,    -2,     4,    -1,    -1,     4,     2,   -19,   -13,   -10,    -5,    -8,    -9,   -30,     1,     5,    -8,    -4,   -24,   -12,    -8,   -13,    -1,     4,    -5,    -2,    -1,     2,    -3,    -1,    -5,    -6,    -2,    -2,   -15,    -6,     5,     7,    -7,     5,    -7,    -4,   -12,   -15,   -19,     6,    -2,   -21,    -8,    -7,     1,    -1,     8,     5,     0,    -3,    -5,    -2,    -9,   -17,    13,     9,     7,   -14,   -14,   -26,   -15,   -29,   -36,   -22,   -11,   -37,   -45,   -31,    -9,   -29,   -31,   -11,    -3,    -1,    -2,     2,    -2,    -5,    -3,    -9,    -7,    19,    23,    31,    23,    24,    17,     1,     7,    11,   -12,   -15,    -7,    -7,   -28,    -9,    -4,   -23,   -21,   -30,   -14,   -11,    -7,   -15,    -1,    -4,    -5,     7,     6,     8,    -2,     7,     6,    11,    19,    12,    11,    -4,   -16,   -24,   -33,    -7,    -4,   -19,   -15,   -13,    -8,   -22,   -16,    -3,     1,   -11,   -10,     3,    -1,   -12,    19,    18,    18,    29,    -1,    -6,     1,    -2,     3,   -12,   -10,   -12,   -13,    -3,     0,    -2,     1,   -18,    -8,    -6,   -20,    -8,   -15,    -8,    -1,     3,     0,     3,    29,    30,    10,    29,    14,    28,    -2,   -13,    -1,    14,    -4,   -21,    -7,    -6,   -19,    -1,    -7,    -9,    -9,   -17,   -44,   -27,   -13,   -17,    -7,   -12,     7,     1,    11,    15,    10,    26,    20,    14,    16,     5,    -4,    13,    -7,    13,    -7,   -31,   -13,   -19,    -7,   -10,   -26,     2,   -16,   -30,   -17,   -26,    -9,     4,    -6,    -3,    -8,     2,    15,     4,     6,    -6,   -10,   -32,   -18,   -12,   -14,     5,     2,    -8,   -22,    -8,    -2,    -1,    -7,     7,    -8,   -27,   -13,     8,    -3,     0,    -4,     2,   -29,   -16,    -1,    12,     1,    -9,   -27,   -23,   -53,   -51,   -23,    -5,     0,    -7,   -10,    -8,    -8,     9,   -18,   -19,    -2,   -12,   -11,   -13,    -2,     5,    -5,   -13,   -18,   -22,   -18,    -6,    -8,   -10,   -27,    -7,   -15,   -48,   -24,   -13,    -6,    -2,   -17,   -11,    -3,    -8,   -18,    -2,    -9,    -1,     3,   -33,    -8,     2,    -2,    -4,     1,   -27,   -48,   -35,   -31,   -27,   -27,   -18,    -8,   -16,   -25,   -14,   -25,   -11,    -5,   -18,     1,   -14,   -11,    15,     5,    29,     9,    -6,    -5,    -4,     0,    -2,    -8,    -8,   -45,   -55,   -48,   -34,   -32,   -21,     2,    -2,    -5,   -10,   -30,   -18,   -20,   -14,     0,    11,    -6,    21,    30,    41,    24,     3,   -10,     5,    -9,    -9,    -6,   -21,   -37,   -54,   -38,   -30,   -17,    15,     7,   -12,   -26,    -3,   -15,   -21,   -31,    -7,    24,     3,     7,    20,    13,     9,     5,    12,    20,     5,   -13,    15,    13,   -16,   -36,   -30,    -6,    -1,     7,    17,    -3,     7,    17,    14,     1,    -8,     4,     6,    39,    30,    15,     3,    19,    26,    25,    18,    30,    -2,    -6,    19,     3,   -13,   -38,    -5,     2,     0,     1,     7,     4,     5,     2,     0,    -9,   -28,     4,    22,    32,     6,    22,    23,    25,     6,    40,    12,    15,     4,    -4,    26,    -6,   -21,    -8,     7,    19,    11,    24,    -2,     0,   -16,   -15,     9,    -6,   -33,    20,    32,    -6,    -3,    14,    -5,    -3,   -27,    24,    -4,    18,     2,     4,     5,    20,   -30,     3,    14,    11,    11,    -5,   -15,   -10,     4,   -18,     2,   -11,     9,    25,    17,   -18,   -23,    -8,   -13,   -12,    11,    30,     4,    42,    -3,   -20,   -12,   -10,   -30,     0,     7,    20,     7,   -12,   -16,    -3,    -9,     1,    -9,    -2,    17,    20,     2,   -16,   -25,   -30,     4,   -18,   -27,     1,    28,    32,    -4,   -18,    -1,    -3,   -21,     0,    11,    11,     9,   -15,   -21,     1,     3,    14,   -11,    -1,     5,    -5,    -5,   -16,   -23,   -24,   -19,   -23,   -33,    -4,     6,     3,     0,     5,     7,     4,   -31,   -19,    -6,   -18,    12,    -5,    -6,     6,     0,     6,    -1,    14,    19,     1,     4,   -12,     0,     4,   -13,     3,   -20,    -5,     8,    -5,    -1,     3,    -2,    14,   -24,   -38,   -19,   -20,   -16,   -15,    -9,    19,     4,    23,    21,    -2,     1,     8,    -1,   -12,     5,     2,   -25,     3,     2,    -3,   -13,     0,     0,     2,    -3,    17,   -23,   -34,   -24,   -17,   -17,     2,    11,     9,    29,    18,     4,     3,     8,    13,   -10,    -9,   -11,    -6,     6,    10,     6,    10,   -16,     1,     1,     2,   -25,   -19,   -38,   -26,   -34,   -14,   -25,   -33,   -29,   -22,   -21,   -22,    -8,   -11,   -30,    -8,     4,    10,     6,   -11,    -1,    10,    16,    -2,     2,     2,    -2,    -3,     2,    -2,    -7,    -7,    -6,    -4,   -16,   -36,   -49,   -36,   -34,   -61,    -5,    -4,   -18,     1,   -10,    14,    15,    11,   -14,    -4,     6,     5,     3,     0,     2,    -4,     3,    -3,    -1,   -17,   -16,   -14,   -13,   -30,    -5,    -8,   -16,   -15,   -21,   -14,   -26,   -33,   -27,   -16,   -15,   -11,   -16,     2,     1,     1,    -3,     1,    -5,     2,     4,    -4,    -4,     1,     3,    -1,    -5,    -1,   -10,    -8,   -10,   -19,   -14,     4,     0,    -8,    -4,    -4,    -7,   -14,   -13,    -1,     5,    -1,    -3,     5),
		    33 => (   -4,    -1,     0,     4,     3,     4,     0,     4,     3,    -2,     4,     0,     0,    -3,    -5,     1,     2,    -5,    -5,     2,     3,     4,    -4,     1,     1,    -3,     1,    -2,     0,     3,    -2,    -4,    -4,    -1,     1,     1,     4,    -5,    -6,    -1,    -4,    -6,    -4,    -5,    -2,    -9,    -3,     4,     0,     0,    -1,     3,    -2,    -2,     3,     0,    -5,     2,     0,     1,     0,     4,    -4,    -1,   -13,   -16,    -7,    -7,   -19,   -17,   -30,     0,   -10,    -6,   -10,    -8,   -17,    -7,    -8,   -10,     0,     3,    -5,    -4,     2,     5,    -1,    -3,     1,     1,     2,    -3,    -1,    -1,     2,     1,    -1,     0,     2,    -5,   -12,   -10,    -6,   -12,    -4,    -3,    -4,   -13,   -15,   -11,    -2,     0,    -3,    -1,     1,    15,    -5,    -4,    -2,    -2,    -4,    -1,     0,     1,    -8,    -8,    -5,    -5,    -1,    -2,   -13,    -8,   -12,    -7,    -2,     0,   -33,   -16,    -9,     2,     1,     0,    -1,     6,    15,    -2,     5,    -3,   -11,   -17,   -14,   -16,   -19,    -7,   -17,    -6,     1,    13,    16,    10,     0,    -9,   -12,   -10,    -8,   -27,    -7,     1,    -1,    -3,    12,    -5,    12,    12,     4,     4,    -2,     3,     7,     3,     9,    -6,    -8,    -9,   -15,   -21,     2,     5,    -6,   -20,   -16,   -11,    -2,    -2,   -19,    -4,     1,     4,    21,     2,    -6,    11,     1,    12,    12,    13,     4,    11,    -1,   -14,   -10,   -19,   -17,    -7,   -15,   -34,   -19,   -14,   -14,   -14,   -11,    -6,   -28,    -6,    -5,     7,    19,    15,    11,    -2,    14,    16,    14,    -8,     4,   -10,   -15,    -2,     5,     7,    -1,     9,     2,     0,   -17,   -10,    -5,    -3,    -5,   -14,   -23,     1,     4,   -21,    43,    10,    13,    -1,    23,     9,     0,    13,    10,   -20,   -14,     2,    15,    -2,   -28,     4,    11,    -3,     0,    10,   -12,     0,   -25,   -26,   -11,     0,     5,   -17,    39,    12,    -5,   -12,    11,     0,   -13,   -24,   -18,   -16,     0,     3,    21,   -20,   -26,    -5,     5,    -6,     5,     8,    -3,    -3,   -22,   -10,    -3,    -3,     1,    -3,   -16,   -13,    -7,   -14,   -24,   -20,   -24,   -29,   -11,     0,     7,   -11,   -19,   -19,    -4,    -2,     5,     1,     5,     8,     8,    -5,   -10,   -22,    -8,     0,     5,     1,   -19,    -8,    -8,   -24,   -29,    -1,    -6,    -9,    -5,     0,   -11,   -36,   -16,    -1,    -2,    11,    12,    -4,    -1,     2,     0,    -7,    -9,     3,     1,    -4,     2,     2,   -12,    -8,    -2,   -12,   -17,     0,     4,     5,   -12,     2,   -10,     8,    -4,    -4,    -8,    12,    -7,    -8,   -17,     0,     4,    -8,   -12,   -10,   -13,   -10,    -2,    13,    -6,   -10,     1,    -3,    -8,   -18,   -10,   -13,    -1,    -4,   -13,     4,    13,     9,     3,   -14,   -22,   -14,   -20,    -7,    -7,    -3,    -9,   -28,   -14,   -10,    -3,     6,    -5,   -11,    10,   -12,   -12,    -6,     1,    -9,    -1,    -1,     3,     6,     8,    -8,     2,    -2,   -13,   -20,   -10,   -10,    10,     0,    -7,     0,    -4,     0,    -3,     0,    -6,    -9,     1,   -12,    -3,   -10,    -3,    19,     3,    -5,    -5,     3,     2,    -8,     1,   -19,    -2,     0,    -6,    -1,    10,     1,    -6,     3,   -20,   -13,    -4,     7,    -4,    16,     2,    -4,    -2,    -6,     1,    15,    -4,     8,     6,    -4,    -8,     1,    -5,   -22,   -20,   -12,    -6,    -1,    10,    -1,   -13,    -5,    -2,    -6,    -7,     2,     1,    13,    13,     9,    -1,   -15,    -1,    12,    24,    -4,     4,    19,    -3,    -7,    -9,   -21,   -21,   -11,    -4,    10,    16,     4,   -10,    -8,    -3,   -11,    -5,    -2,     4,     3,    16,    10,     3,    -7,    -4,    -2,     9,    -9,     8,     2,   -11,    -8,   -14,   -12,   -13,   -12,     7,     6,    22,    17,   -12,    -5,    -9,    -7,    -1,     1,    -4,     5,     6,     7,    10,    -6,   -13,     3,    -2,   -28,    -3,    13,     0,   -14,    -4,    -8,   -12,     3,    -6,     8,    20,    17,   -17,   -14,     0,    -5,     0,     0,     2,     9,    10,     3,    -3,   -17,   -25,    -5,   -13,   -26,   -26,   -17,   -23,    -5,     7,   -10,    -3,     2,    -1,     1,     1,    17,   -13,   -13,    -1,     3,    -7,     0,     2,     7,    19,     5,    -1,   -11,   -26,   -13,   -10,   -28,   -38,   -22,   -34,   -24,   -10,    -7,    18,    23,    10,    -9,    -2,    17,    -5,   -12,    -4,     4,     1,     3,    11,    -5,    -3,    -6,    -5,    -5,   -16,   -27,    -8,    -6,   -19,   -17,   -22,    -4,    15,     6,    11,    -9,     1,     5,     9,     2,   -10,   -14,     4,    -5,    -1,    -1,   -10,     0,    -8,    -8,    -5,     7,   -15,   -19,   -25,    -4,   -29,   -10,    13,    31,    19,     0,   -10,    -6,     2,    -4,   -11,     7,   -19,   -10,    -6,    -2,     0,     0,     8,    -9,   -22,   -24,    -8,     3,    13,     0,    -9,    -8,     6,    31,    44,     7,    14,   -11,    -2,     1,    12,    -1,   -18,   -47,    -3,     0,     1,     1,     1,     3,    -2,   -17,   -18,   -18,   -29,   -21,   -19,   -30,   -16,   -14,    17,    30,    21,    -4,   -11,    -9,    -8,   -11,   -16,   -13,   -25,     4,     4,    -1,    -1,     4,     0,     4,    -1,     5,     1,     1,    -5,     4,     4,   -17,   -17,    -7,   -10,    -9,    -7,   -18,    -1,     2,    -6,    -4,    -9,   -10,    -1,    -1,     1,     1,     3,     0),
		    34 => (   -4,    -3,    -2,     2,     0,     1,    -4,     3,    -1,     4,    -5,    -3,    -1,    -3,     1,     4,     2,     4,    -1,     2,    -2,    -3,    -1,     0,     3,    -4,    -3,     3,    -4,    -5,     5,     5,     2,     0,    -5,   -10,    -9,     3,    -5,     2,     3,   -19,   -15,    -4,    -3,    -8,     1,     3,    -2,    -4,    -7,    -4,     0,    -4,    -3,     0,     4,    -3,    -4,    -4,   -11,     2,    -9,   -16,    -7,    -3,    -8,    -9,    -4,   -12,   -15,    -7,    -4,   -13,    -3,    -1,   -15,    -6,    -6,    -3,     2,     0,     1,     4,     3,    -3,    -1,    -5,    -6,    -5,   -23,   -11,   -18,   -10,    -4,    -7,    -9,   -18,   -28,   -28,   -18,     6,    -1,   -12,    -6,    -1,    -3,    -4,     1,    -5,     0,    -1,     2,    -1,    -1,    -6,    -9,    -3,   -10,    -8,    -3,    -6,    -9,   -10,   -12,   -23,   -33,   -17,    -9,   -11,   -26,   -21,    -4,   -16,   -20,    -5,     5,    -2,    -5,    -6,     2,     5,     3,    -6,    -7,    -2,   -10,    -4,   -12,   -16,    -5,   -20,   -32,   -19,     0,    13,    -7,   -41,   -37,     1,   -13,    -6,    -8,    15,    17,     2,   -15,    -4,    -3,    -1,     4,   -12,    -8,    16,   -13,    -3,   -13,   -12,   -19,   -13,    -6,     0,    30,     2,   -61,   -74,   -24,     4,    28,     1,    17,   -16,     6,    -6,    16,   -26,    -5,   -28,     1,    -4,    -5,    23,    -5,    -4,     3,   -12,   -32,   -19,    13,    11,    11,   -50,   -66,   -51,    -9,    14,     6,    -3,    16,    11,     7,     7,     1,   -14,    -9,   -24,     6,    -4,    -4,     3,     3,    13,    -2,   -10,   -34,     5,    16,    18,   -23,   -27,   -56,   -14,     4,     2,     7,    -3,    15,     5,    11,    -2,    -9,   -21,     3,   -20,     8,    -5,     2,    -9,   -16,    -6,   -17,   -23,   -20,    24,     3,    -1,   -15,   -50,   -38,    -4,     7,    13,     9,     2,     6,     3,     4,   -11,    -2,   -10,    -5,    -3,   -15,    -2,    -1,   -24,   -20,    -5,   -21,   -22,    -5,    25,    -1,   -17,   -33,   -16,   -11,    -8,    -5,     1,    -5,   -24,   -35,     2,   -23,    -2,    -9,    -9,    -3,    -2,   -17,   -10,   -16,   -18,   -11,   -21,    -4,    -8,     7,    12,     1,   -13,    -1,    15,    -8,     1,     0,    19,    -9,   -10,   -20,   -25,   -16,    -7,   -18,   -24,     5,     0,   -29,   -20,   -29,   -15,   -22,   -12,   -14,     2,    10,    -7,     1,     0,     6,    -6,     2,    -7,    -7,     3,    -5,     9,   -10,   -22,   -15,   -14,   -38,   -26,    -4,    -3,   -20,   -19,   -31,   -15,     0,    -8,     0,     2,    29,     8,    -9,     7,    13,    12,    15,    -6,   -18,    11,    13,     6,   -20,   -26,   -24,   -33,   -38,    -4,    -2,    -4,   -13,   -30,   -30,   -11,   -14,    -5,   -13,     3,    11,    -2,    -6,     6,    -4,    17,    14,   -17,     2,    11,    25,     9,   -20,    -7,   -15,   -16,   -18,    -3,    -2,     1,    -7,    -6,     5,   -13,   -20,     3,    -4,     5,    -4,    -7,    -5,    -3,    -1,    24,   -13,    -2,   -11,    21,   -17,     4,    -1,     7,   -15,   -11,    -6,     7,    -4,     4,    -8,     1,    -1,     7,   -14,     0,    10,    13,   -12,   -14,    -6,     7,     1,    -3,   -11,   -21,   -35,   -12,   -19,   -16,   -11,     5,     5,     1,    -7,    -4,     5,     2,   -16,    -3,   -10,   -12,     2,   -10,    10,    -4,   -19,    -6,   -12,   -17,   -11,    -3,    11,   -24,   -28,   -22,   -16,    -3,    -7,     8,    -3,     1,     1,    -8,    -6,     3,   -16,     6,    12,     1,    -5,    -2,   -27,   -29,   -22,    -2,   -10,    -9,    -3,    -5,     0,   -24,     0,    -3,     5,     1,    -7,     1,    -2,    -4,     3,    -5,     2,   -19,   -21,     6,    19,    -9,   -26,   -22,   -27,   -16,   -28,     1,    -1,    -8,    -6,    -4,     0,   -17,    -3,     8,     0,   -11,   -16,     1,    -3,     4,     2,    -6,     1,    -4,    -3,    -9,     4,   -15,   -38,   -23,   -37,   -13,   -10,     8,   -12,   -13,   -18,   -30,   -12,   -22,   -11,   -10,   -12,   -12,    -4,     6,     5,   -11,    -5,     3,     1,     4,   -10,   -16,    -1,   -14,   -47,   -29,    -3,    -1,     1,    -8,     0,    -9,   -16,   -19,   -35,   -19,     2,     2,   -11,   -17,    10,     7,     8,   -28,    -8,     1,    -5,     4,     3,   -12,   -15,    -1,   -18,   -25,     2,     2,     7,    17,     4,    -8,   -25,   -10,   -18,   -10,     7,   -15,   -11,    -1,     5,     2,     5,     1,     1,    -4,    -4,     5,   -10,    -8,    -7,   -21,   -14,   -16,     6,    -8,     5,     0,   -17,   -29,   -18,    -5,    -9,    -6,    21,    14,   -23,    -2,     4,    14,     8,     5,     2,     0,     3,     3,     0,    -5,   -21,   -11,    -3,    -5,     5,     7,    16,     7,   -23,    -2,    -5,    10,     0,   -10,    25,    22,    14,     8,    12,    10,    -3,    22,    -1,     5,    -1,     0,   -12,     3,   -18,    -5,   -22,   -11,   -21,   -18,     4,     3,     9,     6,     2,   -10,   -18,    -1,    19,    22,     6,     3,    18,     7,     8,    -3,    -4,     4,     1,     0,     2,    -4,   -17,    -4,   -12,   -15,   -15,   -20,     3,    -9,     8,    -6,   -25,   -11,    -3,   -11,   -25,   -12,   -13,   -38,   -35,    -1,    -7,     0,     0,    -4,     4,    -2,    -1,     5,     2,    -1,    -8,    -2,    -2,    -8,   -31,   -30,   -21,   -19,   -23,    -3,   -13,   -27,    -8,   -18,   -13,   -11,    -8,    -6,    -5,     2,     3,    -2),
		    35 => (    5,    -2,     4,     3,     0,     1,    -3,     1,     1,     4,    -4,    -2,    -4,    -3,     5,    -1,    -1,     2,     2,     0,    -1,    -3,     1,     2,    -2,     4,     4,     1,    -3,     0,     2,    -2,     3,    -1,    -4,    -1,    -3,    -2,     2,    -8,    -7,    -5,    -5,    -9,   -15,   -14,    -5,   -10,    -2,    -7,    -4,    -3,    -1,    -2,    -5,    -3,     4,    -5,    -4,    -7,    -8,     4,   -13,   -11,   -11,   -21,   -25,   -20,   -28,   -25,   -60,   -40,   -23,   -13,    -9,     7,     1,   -28,   -11,     5,   -12,    -9,     1,     1,     4,     3,    -2,     2,    -4,   -25,   -20,   -17,   -39,   -42,   -33,    -8,   -10,    -3,    -8,   -10,   -18,    10,    28,    12,   -17,    -9,   -10,   -16,   -16,    -3,     2,    -4,    -1,     2,    -8,     7,   -16,    -8,   -26,     1,    -9,    -3,    14,    -8,   -27,    -9,    13,    17,    -5,   -13,     2,   -17,   -19,   -10,   -21,   -31,   -35,   -25,    -7,    -5,    -2,     0,    -5,    -5,   -16,     2,   -15,   -35,   -26,   -14,   -14,    -6,   -26,   -23,   -12,   -24,   -23,   -41,   -45,    -7,     9,   -18,   -19,    -6,   -24,   -31,    10,     6,    -2,    -1,    16,   -23,   -25,    12,   -14,   -19,    -6,   -19,     5,    -8,   -22,   -10,     1,   -12,   -20,   -16,    -7,    -6,    -2,    -3,     1,    -5,     0,   -29,    -4,     1,     3,    -6,    17,   -12,   -29,    12,   -27,   -12,    -5,    -4,    34,     7,   -10,    -2,    -2,     6,   -21,   -23,   -39,   -40,   -12,    -4,     3,     4,   -12,    -7,    -1,    19,    -4,    -1,   -20,     2,   -10,    -6,   -15,    -3,    -2,     3,     8,    12,    -8,    -8,    12,    10,    14,    11,    -1,    17,    17,    17,    25,    26,    24,    17,   -15,    12,    -1,    -2,   -21,   -15,   -11,   -36,     8,    12,    -3,    -4,    -5,   -18,   -10,    -3,    13,    12,    27,    44,    31,    36,    24,    29,    25,    18,    42,    34,   -24,     5,    -2,    -4,    -5,   -16,    -2,    -7,    10,     8,    -9,    -1,     2,    20,   -11,    -2,     5,     8,     4,    16,    36,    32,    31,    39,    27,    13,    46,    33,    16,    24,     4,    -6,    -2,    -5,     7,     0,    -9,   -22,    -9,   -16,    10,    -6,    -9,   -17,   -35,   -30,   -26,   -27,   -20,   -33,   -22,     6,     4,    16,     5,    38,    34,     2,     0,    -5,    -2,     4,    -8,   -13,   -17,    -6,    -1,    12,    16,    23,    12,     0,   -17,   -23,   -39,   -34,   -68,  -111,   -70,   -47,   -47,   -28,   -23,    23,    35,   -11,     0,     0,    -5,     8,    -8,   -24,   -28,    11,     1,    -6,    29,    10,    18,     4,     5,     0,   -19,    -1,   -24,   -47,   -62,   -39,   -54,   -55,   -19,    -8,    24,   -11,     9,     3,    -6,    -8,    12,    -2,    10,     7,    20,    18,    -1,     2,    -4,    -4,    -6,    -1,   -10,     8,    -1,   -38,   -41,   -31,   -27,   -19,   -20,   -25,    -7,    -5,     6,     1,   -20,    19,    33,    15,     6,    25,    16,    19,    -4,     2,     7,    -3,   -16,   -18,   -30,    -8,    11,    -1,   -17,   -16,   -30,   -13,   -21,    10,    -7,   -15,     1,     1,   -18,     3,    12,    34,    -4,    18,    -1,    11,    -1,   -12,   -10,    -4,   -29,   -12,   -17,    -7,     9,     0,    -2,   -14,   -11,   -16,   -10,    10,   -18,   -20,     4,    -4,   -35,     5,     9,     9,     6,   -14,    -7,     9,     4,    -6,   -23,   -23,   -21,    -2,   -11,    -2,   -14,    -1,   -11,   -21,    -7,    -7,   -34,   -37,   -35,   -35,    -9,    -5,   -19,   -36,   -17,   -11,     1,   -10,   -12,   -19,   -39,    16,    19,   -10,   -20,     5,   -15,     3,    -9,     1,    11,   -21,    -4,    18,     4,   -13,   -38,   -24,     1,     0,    -5,   -31,    14,    21,    -7,   -13,    -8,   -27,   -34,   -33,    -2,    14,   -22,   -17,    -8,     6,     4,    17,     2,   -24,     8,    31,    30,    35,   -33,   -26,    -1,     1,    -6,   -21,    17,     0,   -15,    -4,   -15,   -13,   -18,     1,     7,    13,   -42,   -13,     5,     0,     2,    13,     9,   -18,     6,     5,    36,    41,   -28,     0,     0,     4,    -6,   -15,    -7,    11,   -17,   -19,    -6,    -3,     4,     5,     9,     6,   -12,    22,    -6,    -2,    -4,    -3,     6,   -12,   -20,     1,    28,    47,    23,    -4,     0,    -2,   -15,    -3,    -7,    11,    12,   -16,   -25,    -2,     3,     7,    18,     5,    -1,    14,     7,    14,    -1,   -18,     4,    -4,   -17,    32,    55,    54,    54,     4,    -4,    -1,    17,    -4,     0,     1,    -9,   -23,   -22,    14,    22,   -11,     0,   -14,     6,     8,    -9,    -2,    -1,   -18,     1,   -16,    -3,    52,    54,    49,    63,    -4,     5,    -4,    -4,     0,   -25,   -35,   -26,   -17,   -10,   -14,     3,     8,    17,    -7,    17,    -6,    -5,    -8,   -12,   -11,     2,    14,    35,    18,    14,   -38,   -12,     3,     2,     2,    -2,     2,   -35,   -38,   -23,   -33,   -25,   -14,   -18,     3,    36,    19,    -4,   -22,   -15,   -13,     6,    -1,   -19,    16,    20,    27,    28,    -4,    -6,    -4,    -2,     0,    -2,     1,   -20,   -42,   -57,   -54,   -50,   -48,   -43,   -29,   -30,   -45,   -73,   -19,    -3,   -11,    -6,     6,    -1,     9,    -1,   -22,   -11,     3,     4,    -1,     2,     2,     4,     2,     0,   -10,    -4,   -12,   -11,    -6,    -3,    -9,   -11,    -8,   -39,   -21,    -8,   -16,   -22,   -14,   -10,   -17,   -37,   -26,    -4,     4,    -3,     0),
		    36 => (    0,     3,     1,     3,     0,    -2,     3,     1,    -4,    -3,    -3,    -1,     6,     3,     0,    -2,     3,    -4,    -2,     4,     3,     2,     3,    -2,    -3,     1,    -3,    -1,    -4,    -3,     3,    -5,     2,     4,    15,    17,    16,    12,    23,     4,    -1,    10,   -15,     1,     3,    10,    22,    14,    43,    17,    17,    16,     5,     2,    -1,     4,    -3,     1,    13,     8,    22,    19,    21,    27,    15,    -9,   -12,   -16,   -22,   -22,     3,    12,    19,    37,    20,     9,     7,    39,    36,    27,    18,    26,    -5,    -2,    -2,    -1,   -30,     4,   -10,    14,    27,    25,     1,   -12,   -13,   -38,   -51,    -1,    23,    15,   -19,   -13,     7,   -12,   -12,    -2,   -20,     6,   -30,   -15,   -23,    -3,     1,     3,   -40,    -5,    13,    32,    24,   -10,   -26,   -22,   -29,   -50,   -65,   -27,   -35,   -18,    -1,   -14,    -7,    43,    28,     6,   -33,   -38,   -60,   -44,   -17,    12,     1,     0,   -19,   -23,    12,    25,    12,    -8,   -12,   -11,   -18,   -55,   -38,     2,     5,   -19,   -10,     0,    12,    13,    23,    16,   -12,     2,   -29,   -43,     2,     3,    -4,    -3,    19,     6,     7,    24,    23,    -2,    -7,   -29,   -31,   -22,   -14,   -18,   -15,    22,    16,     5,     2,    -3,     1,     2,     9,   -16,   -13,   -34,   -16,    -5,     0,    -3,    -3,    -9,    -8,     4,   -11,     1,   -19,   -34,   -58,   -43,   -14,   -17,    10,    15,   -16,   -23,    -8,   -40,     4,    -5,    18,   -22,   -50,   -46,    -9,   -19,     1,     0,   -20,   -15,    -9,     4,    16,   -18,   -28,   -55,   -54,    -9,    -2,    -5,    -6,     7,    -1,   -18,   -47,     0,   -17,   -21,   -20,   -53,   -46,   -21,   -18,   -25,     1,     0,   -18,   -13,    27,    -8,    -4,    -4,   -30,   -28,   -15,    -3,    -8,     5,    16,     8,   -21,   -36,   -48,   -60,   -74,   -70,   -65,   -59,   -47,   -26,   -27,    -8,     4,     3,   -17,    -9,   -17,   -19,   -24,   -22,   -48,   -13,     6,    -1,     5,     8,     1,    -4,   -20,    -7,   -10,   -42,   -43,   -42,   -53,   -59,   -41,   -34,   -24,   -19,    -2,     1,     5,   -30,   -12,    -5,    -6,   -12,     6,     1,     6,     7,    14,    13,    -6,   -29,   -25,   -11,   -20,    -7,   -12,   -21,     0,   -51,   -52,   -48,   -31,   -26,     5,    -4,    -6,   -20,   -19,    -6,    -3,   -20,    -2,     5,    18,    13,     7,    31,   -11,     4,   -22,    14,    -5,    -1,    -9,   -18,     8,     6,   -21,   -48,   -49,   -25,    -4,     2,    -6,   -25,   -20,   -11,   -19,   -24,     5,     3,     9,    33,     7,    16,     1,     3,    -7,    10,    33,     0,     5,     2,    33,    28,   -28,   -55,   -26,    -1,    -2,     2,    -2,   -31,   -21,     5,   -27,     1,    -9,    12,    19,     6,     0,   -12,    -9,    -1,     1,   -42,     8,    16,    -2,    28,    20,     2,     7,   -19,   -25,     0,     1,     5,     1,   -26,    -3,     7,   -16,    -1,    12,    10,    11,   -22,    -8,   -10,    -1,   -29,   -24,   -30,     8,    22,    11,    34,    13,     6,   -25,   -36,   -43,   -25,     0,     3,     0,   -10,    -8,    10,    -4,    19,    -5,    13,     2,    13,    22,    16,    14,     0,     7,    -1,     1,    -3,    15,    30,    17,    -3,   -34,   -39,   -41,   -33,     0,    -2,    -2,     2,     6,    10,     3,     6,    23,    -1,     8,    13,   -12,     1,    -8,   -13,   -12,    -5,    -2,     1,    12,    27,    -9,    -8,   -32,   -26,     0,   -33,    -1,    -5,     2,     1,    24,    -6,   -15,    -7,    -5,    24,    15,   -13,    -7,   -11,    -3,    26,    -5,    12,    18,    10,     6,    -6,   -48,   -38,   -28,   -24,    -5,   -14,     0,   -11,   -14,     5,    17,   -17,    -7,     0,   -15,     6,    11,    21,    -1,   -38,   -14,    10,    -4,    -4,    16,   -10,    -8,   -19,   -51,   -21,   -11,   -11,   -17,    -5,    -4,   -12,   -10,   -31,    21,     8,    -7,    -7,    -6,   -12,     5,    19,    19,   -11,    -3,    -6,   -28,   -19,   -28,    -8,    -2,    -3,    -7,   -25,   -13,   -16,   -21,     3,     2,    -4,   -15,   -15,   -14,   -18,    -1,    -5,    -3,     0,    -9,    21,   -10,    -5,   -11,   -25,    -9,   -15,   -10,   -18,    -7,     4,   -21,   -17,   -16,   -17,   -16,    -4,    -3,    -1,    -6,   -11,   -21,   -28,   -31,   -16,   -19,   -10,     1,     3,    10,    15,    -1,     6,    -9,   -22,   -10,   -19,   -33,   -29,    -8,   -19,   -39,   -17,     4,    -5,    -1,     3,     3,    -6,   -12,   -17,   -20,   -33,   -23,   -29,     0,    13,    10,    -2,     9,    16,   -20,   -38,    20,    30,    18,    -3,    -3,    -7,    -8,    -4,    -8,    -5,    -5,    -4,     2,     4,    -8,    -3,    -3,   -12,   -21,   -32,   -36,   -36,   -17,    -7,     7,    24,    30,     1,    -3,   -37,   -23,    -7,    -8,     0,    -2,    -3,     5,     4,     3,    -1,     5,     5,     5,    -3,   -11,   -16,   -11,    -4,   -16,     9,    21,     4,    -4,     0,    -5,    -5,    -1,    -7,   -16,    -4,     3,     0,    -5,     4,    -2,     4,     2,     0,    -4,    -4,     0,     0,     2,    -1,    -1,    -1,    -2,    -2,     3,    -4,    -1,    -7,    -7,     1,     1,     4,     0,    -7,     0,    -6,     1,    -3,     4,     1,     2,    -3,     4,     1,     1,     2,     4,    -4,     2,     3,    -6,    -1,    -5,     0,    -5,     0,     1,    -6,    -6,     3,     2,     1,     3,     1,     5,     1,     4,     0),
		    37 => (    0,    -4,    -1,     2,     1,     2,     2,     1,     0,     1,    -1,    -4,     0,    -3,     5,     0,     1,    -2,    -2,    -4,     2,     2,    -4,     1,     3,     4,    -5,    -4,     0,    -5,     2,     3,    -2,     0,     2,    -3,    -3,    -5,    -2,   -17,   -21,   -13,   -10,   -16,   -20,   -16,    -6,     1,    -1,    -1,     4,    -3,     2,     4,    -5,     2,    -4,     2,    -1,   -12,   -12,     1,    -4,   -14,   -24,    -9,    -2,   -21,    -9,    -2,     1,    -2,    -1,    -6,    -6,     3,    -2,     1,     1,    -4,     3,     0,     3,     2,    -4,     4,    -4,    -9,    -7,    -5,   -14,   -36,   -35,   -11,   -19,   -17,   -12,   -15,    -8,   -10,   -10,   -24,   -11,   -17,    -6,    -6,    -9,    -1,    -4,     2,    -5,    -1,    -4,    -1,     3,    -6,   -24,   -18,   -14,   -21,   -38,   -36,   -37,   -42,   -42,   -20,   -37,   -29,   -20,   -19,   -21,    -7,   -11,   -14,   -17,   -16,   -17,    -7,     2,     4,    -2,     4,     3,   -29,   -46,     7,   -14,    13,    42,    13,   -26,   -38,   -21,    16,   -12,    -7,   -45,   -53,   -37,   -56,   -46,   -24,   -24,   -24,    -7,   -22,    -3,    -4,     2,     1,     7,     9,    -4,     1,    -3,   -19,     0,    -8,   -33,   -19,   -22,   -27,   -10,   -19,   -43,    -4,    12,    -4,     0,    26,     2,   -22,   -34,    -4,   -35,   -11,     2,     6,     7,    14,    13,     5,    12,    17,     3,     0,     4,   -25,   -14,    -8,   -13,   -30,   -25,    -4,     0,   -49,   -28,    -7,    -6,   -14,   -31,   -15,   -15,    -8,   -12,     6,   -18,     4,    16,    20,    32,    12,     3,    27,    -3,     5,    11,     3,   -23,   -14,   -14,   -12,    13,   -23,   -10,     1,   -10,     5,     1,   -16,   -28,    -8,     2,     9,     0,     7,    43,     1,     6,    -2,    -4,     5,   -20,    10,    27,    14,    21,    13,   -16,   -15,    -3,   -10,     3,    21,    17,    36,     7,   -23,   -17,    20,     1,    24,    14,    17,    46,    20,    21,   -17,     2,    15,     0,    17,     4,     0,    17,    20,    -4,    -1,    -5,    -1,    -8,    -7,    39,    15,   -29,    -3,   -15,    20,    -3,    15,    38,    32,    40,     7,   -15,    -3,   -12,    -1,     6,    15,    -2,     5,     7,     9,   -16,   -12,   -10,     3,   -19,    12,    13,   -11,   -44,   -37,    -9,    32,     4,     5,     5,    44,    19,     8,    -6,    -6,    -9,    -7,    -5,     4,     4,    -9,     8,     8,     4,   -15,    11,     6,    -4,    17,    22,   -26,   -23,    10,    -9,    24,     5,    16,    18,    40,    16,    11,   -14,   -11,   -22,   -17,    13,    10,    -6,   -28,     9,   -19,     2,    -7,    -8,   -11,    33,    22,     8,    -6,    -3,    26,   -12,   -12,    -7,     9,    41,    41,    -4,    17,   -13,   -23,   -16,    -3,    17,    13,   -18,   -50,    -9,   -11,    -1,    14,     0,    23,    17,    18,    10,    35,    34,   -15,   -18,    -5,    -2,     4,    24,    21,   -17,     3,     6,     1,    -9,     2,    20,     0,   -26,   -31,    -3,   -19,   -18,     6,     5,    35,    13,     6,    22,    16,    13,   -24,   -11,    -9,     0,     1,    10,     6,    28,    10,   -11,    11,    10,    28,     2,    -7,   -49,   -22,   -16,     2,    -7,     2,     3,    14,     1,    30,    42,    38,    16,   -60,   -26,     2,    -5,    -2,   -10,    -2,    16,     8,   -15,     1,    13,    12,   -19,   -26,   -41,   -36,    12,     9,     5,    -7,    -4,    -7,    11,    16,    42,    20,     0,   -58,   -16,   -37,    18,     4,    14,   -44,     0,     3,   -15,     9,    13,     5,   -16,   -35,   -79,   -29,    23,    16,     4,     0,    -3,   -17,     5,    11,    21,    -5,   -30,   -14,    -2,   -13,     1,    16,    -5,   -40,    -9,     5,    17,     6,     2,    -7,   -48,   -87,   -73,   -23,    27,     1,   -12,     5,   -17,    -9,   -13,   -38,   -56,   -28,   -22,   -25,    -1,    -2,    -2,    10,    -4,    -8,     8,    26,    20,    20,     3,   -47,   -66,   -90,   -25,   -10,     2,     1,    -6,   -11,   -16,   -19,   -24,   -28,   -41,   -38,    -4,   -20,     2,     3,    -1,    -4,    -5,    -9,   -21,    16,     6,     8,   -24,   -46,   -55,   -45,     0,   -20,     6,    12,    16,   -15,   -17,   -18,   -26,   -14,   -21,   -35,   -35,   -13,    -3,     1,     0,     1,    -3,    -6,     0,    -2,     5,   -10,   -31,   -29,   -47,   -24,    -7,   -10,    10,     0,     0,     3,     4,     7,     7,   -12,   -19,   -22,   -16,   -14,   -22,     3,    -4,     2,   -10,    -9,     6,     8,    -5,   -13,   -31,   -28,   -41,   -24,     5,    -5,    21,    10,    -2,     3,    25,     1,    -2,   -18,   -21,   -32,    -1,    -9,   -16,    -4,    -3,     3,    -6,    -1,     4,    -4,    -2,   -15,   -25,   -27,   -35,   -16,     6,   -12,     0,    -6,    -6,     8,     4,    15,    -2,    -4,    -8,   -33,    -1,    -1,    -4,     4,    -1,     2,    -9,    -1,    -2,    -5,     3,    -6,   -19,   -22,   -42,   -21,   -24,   -14,    15,    -5,    19,    17,    13,    19,     5,     4,     9,   -40,    -2,   -12,     2,    -4,     3,    -1,    -5,     1,     1,    -6,    -1,     5,    10,     6,    -8,   -42,   -27,   -13,   -39,   -15,    14,    11,    15,    28,     4,     8,     8,    -8,    -9,     4,    -1,    -3,    -1,    -5,    -5,     3,     2,    13,   -16,   -15,     2,    20,    17,     0,    -6,   -26,   -31,   -14,    17,    20,     4,   -22,     3,    24,    15,    20,     4,     3,    -3,     1),
		    38 => (   -2,     0,     0,     2,     4,     3,     3,     1,    -2,    -3,    -1,     1,     2,     2,     0,    -2,     2,     4,    -4,     0,    -4,    -2,    -4,     1,    -1,     3,     3,     3,    -4,     4,     0,     5,    -4,     4,    -3,     5,    -4,     2,     2,    -4,     4,    -5,    -9,   -19,   -23,   -11,   -10,     0,    -9,    -3,    -8,    -5,    -3,    -2,    -5,     3,     1,     2,    -7,    -2,     0,    -5,    -1,     1,    -9,   -10,   -19,   -16,     2,    -5,     1,   -12,    -7,   -13,    -6,    -4,   -17,   -19,   -24,   -11,    -3,    -9,    -1,    -3,     3,     3,    -8,    -3,    -2,   -17,    -7,   -25,   -24,     2,    -3,   -16,   -15,   -18,     2,    16,    16,    13,     5,    -9,   -11,    -6,    -2,     4,    -3,    -2,   -13,    -3,    -3,    -4,     5,   -10,   -28,   -12,    -3,    -2,     3,    -4,    -8,    -4,   -13,   -17,    -5,     6,     9,     3,     6,     5,    19,    14,   -15,    -7,   -29,   -13,    -4,   -11,    -5,    -1,    -7,   -24,   -28,   -10,    -2,    -9,   -15,   -19,   -17,   -20,   -22,   -22,   -17,     9,    -6,    -5,    10,    13,    15,     2,    -1,   -19,   -11,     0,     1,   -15,    -2,     2,   -11,   -14,    -2,     6,   -12,    -6,    -9,   -21,   -31,   -32,   -25,   -16,     3,     5,     0,    -1,    -7,    14,   -10,    16,     4,     1,   -19,    -4,    -3,    -1,     4,   -18,   -13,    -8,     6,    -3,    -2,     2,     7,    -3,     6,    -7,    -6,    13,     4,     9,    -3,   -15,   -10,    -2,    -2,   -15,    -1,    -6,   -13,    11,    18,     7,    -8,   -11,    -7,     2,     2,     3,     2,     4,    -7,    12,    11,     0,     2,    -2,    28,    25,     6,     3,   -13,     1,   -14,    -8,   -16,    -4,    19,    36,    26,    11,     4,   -10,    -3,     4,    -6,    -9,   -10,    -5,   -21,   -20,    -3,   -14,    -6,    -1,    10,    18,     3,   -18,   -20,     1,   -12,    -4,     5,    22,    24,    23,     9,   -33,     2,    -5,     0,    -1,    -9,   -12,   -14,   -12,   -12,     6,   -13,   -25,   -21,   -13,     3,    -5,    -7,   -10,   -26,   -13,    -4,    23,    21,     9,     0,   -33,   -18,   -30,    -1,    -2,    -5,    -2,    -8,   -11,   -16,   -10,   -18,    -5,    -5,   -23,   -11,   -12,     9,    -8,     6,   -15,    -5,     6,   -15,    -4,    23,     0,   -10,   -19,    10,   -20,     3,     3,    -3,   -15,    -6,   -15,   -11,   -23,   -30,    -3,     4,    -1,     5,     4,    -5,    10,    -7,     5,    10,     3,    16,    12,    -1,     0,    -2,   -28,   -16,   -31,     1,    -4,   -16,   -26,    -7,    -9,   -31,   -24,   -16,   -12,   -18,    -6,   -11,     7,     2,     3,    10,    18,    -9,    -7,   -19,   -16,     4,    -2,     2,   -14,    -5,     7,    -2,    -2,    -5,   -32,   -12,   -20,    16,    10,   -15,   -41,   -32,     4,    -2,    16,    11,     5,    13,   -15,   -17,   -35,   -10,     4,     2,     5,     0,     3,    -9,   -11,    -5,    -4,     0,    -4,    -8,    -4,    29,    11,   -18,   -18,    -5,    10,    13,     9,     1,    -5,    -4,   -22,   -40,   -19,   -12,    -5,     2,   -17,   -20,     2,   -16,    -9,     3,    -2,    -7,    -9,    -6,    10,    15,     3,     9,    20,    13,    16,     7,   -17,   -27,   -21,    -2,   -29,   -44,   -28,   -19,    -7,   -14,   -24,   -18,     0,   -29,   -14,     3,    -8,    -1,    -7,    -2,     9,    25,    42,    32,    24,    16,     0,   -22,   -13,   -20,   -13,   -25,    -3,   -21,   -15,   -16,   -29,   -17,   -18,   -11,    -6,     3,    -6,     2,    -4,     1,    -3,    -3,    15,    27,    24,    22,    13,   -12,   -22,   -34,     1,    17,   -16,   -22,    -4,     3,    -6,   -17,   -26,   -25,    -9,    -5,    -9,     0,   -14,    -1,     2,    -4,   -18,     8,    31,    14,    -5,     4,   -15,   -36,   -21,   -12,     7,     2,    -5,   -16,     3,     7,   -23,   -14,   -26,   -21,   -13,    -4,     0,   -14,   -10,    -2,    -4,    -2,   -21,    -7,    27,    -6,     9,     5,   -21,   -25,   -19,   -22,   -11,   -12,    -9,   -11,   -11,   -12,   -24,   -29,   -24,   -23,    -5,    -7,    -3,   -13,    -2,   -13,   -10,    -8,   -18,    -3,    22,     3,     3,    12,   -15,    -7,     3,   -17,   -16,   -14,   -22,   -19,   -13,   -27,   -35,   -33,   -28,    -9,    -6,    -2,     0,   -14,    -1,   -13,   -10,    -4,   -12,     5,    -3,     3,     5,    14,    -8,    -4,     2,   -21,   -19,   -10,   -24,    -5,   -17,   -23,   -18,   -28,   -24,   -11,    -6,   -10,    -3,   -13,    -3,     1,     1,     2,   -17,    -8,   -15,   -18,     5,     0,    10,     4,    -1,    -9,    -4,   -14,     1,     5,   -15,   -32,   -23,   -25,   -16,    -2,    -6,    -5,    -7,   -24,     0,     0,     1,    -6,    -6,   -19,    -7,    16,    24,    21,    30,    11,     6,     6,    -5,   -19,     3,   -13,   -16,   -17,   -13,    -7,     0,    -1,     1,   -11,    -8,    -8,     0,     1,     0,    -7,    -6,    -9,   -21,    -3,    14,    12,     3,    -6,     2,     9,    -8,    13,     3,    -7,   -11,    -7,     1,     1,     2,     3,    -1,     0,    -5,   -12,     1,     0,     0,     1,   -20,    -5,   -16,   -21,   -20,     6,     2,     4,     0,     5,    -9,   -13,   -15,    -3,    -6,    -3,    -3,   -20,    -9,   -13,     2,     1,     5,     5,    -5,    -4,    -2,    -2,    -3,     0,   -10,    -4,    -5,    -5,    -3,    -2,    -2,     1,    -8,    -1,    -3,    -2,    -3,    -5,     1,     3,    -1,    -3,     4,    -4,     3,    -2,     1),
		    39 => (   -2,    -2,     1,    -1,     3,    -4,    -1,    -3,     1,     0,    -3,     3,    -5,    -1,     2,    -4,    -5,    -3,    -3,    -4,    -2,     4,     1,    -4,     0,    -2,    -2,     1,    -5,     4,    -4,    -5,    -3,     2,    -2,    -4,    -3,     3,    -4,    -2,   -18,   -16,    -1,    -9,   -10,    -8,   -15,    -8,    -1,    -5,    -3,    -2,    -4,     1,     4,    -3,     4,     1,     4,    -4,     3,     3,     1,    -3,    -6,   -14,   -12,   -12,    -5,     3,   -13,     1,    -1,    -3,     1,     3,    -5,    -8,   -12,     1,    -2,     3,     1,    -1,    -3,     1,     1,   -11,    -8,    -3,    -6,    -9,   -22,   -32,   -19,   -32,   -14,   -20,   -12,   -18,   -10,    -7,    -9,    -8,   -25,   -19,    -7,     1,   -11,    -6,     3,    -3,     5,     4,     0,    -8,   -17,   -24,   -44,    -7,   -19,   -19,     0,    -6,   -13,   -24,   -30,   -37,   -18,   -19,    -6,   -10,   -12,    -4,    -5,    -1,    -5,   -31,    -4,     1,     4,     3,     4,    -4,     0,    -3,   -15,   -16,   -27,     5,    16,     1,    -3,    12,   -18,   -29,   -15,   -24,   -46,   -20,   -17,   -26,    -6,    -9,    -4,   -11,    -7,     0,    -3,     3,    -2,   -17,   -20,   -38,     5,   -13,    15,    16,    23,     7,     3,    30,     3,   -20,   -33,   -22,   -42,   -16,   -40,   -16,    11,     4,   -23,    -5,    -3,    -5,     5,    -7,   -22,   -19,   -29,   -33,   -24,   -13,     3,    25,    10,     3,     1,     8,    -8,   -33,   -12,   -32,   -14,   -26,   -45,   -16,     7,    -1,   -14,   -10,   -11,    -6,   -11,    -9,   -21,   -19,   -22,   -16,   -21,   -13,    -4,   -10,    -4,   -16,     3,    10,    16,   -11,   -25,   -14,   -28,   -13,   -22,   -25,     2,    -1,    -9,   -13,    -4,     0,     0,    -5,   -27,    -7,    -3,    -9,     7,    23,    10,   -14,   -21,    10,     4,    13,     9,    -7,   -13,    -7,   -15,   -28,   -16,   -31,   -18,   -19,   -26,   -23,    -7,    -4,     1,   -13,   -20,     1,    25,   -10,    16,     0,    10,   -16,    -4,    -4,   -10,    -6,   -13,     8,     3,    -8,    -4,   -26,   -19,    -7,   -47,   -50,   -26,   -18,    -1,   -14,    -1,   -28,   -11,    17,    -6,    -4,    34,    21,   -13,   -27,   -13,   -21,    -9,     8,     8,    16,     7,    19,   -14,     3,    -8,   -17,   -38,   -29,   -22,   -43,    -3,   -16,    -4,   -25,   -15,    10,    -4,    20,    23,   -12,   -13,    -5,   -18,   -33,   -11,    -6,    14,    11,    -5,    12,     2,   -10,    -2,    10,   -20,   -15,    -4,   -29,   -23,   -10,    -4,   -25,   -11,    -1,   -17,    24,     0,    -4,     2,    -5,    10,   -24,   -12,    -6,     3,   -17,    -8,    -1,    10,    -3,    12,    10,    -3,   -22,     1,   -21,   -13,    -7,    -8,    -6,    -7,    24,     1,     8,     4,    -3,    -5,    18,    20,    23,     4,     8,   -11,   -34,   -19,     5,    19,    -3,   -11,    11,     5,    -4,    10,   -30,   -12,     1,    -3,    -2,    -7,    22,    11,    15,    14,   -17,     7,     7,    -4,    10,    21,   -20,    -7,   -25,   -36,   -10,    11,     7,     8,    -4,    -5,    -1,     8,   -31,   -19,   -13,    -3,    -5,   -17,     6,    28,   -20,    13,    -7,    -3,    -9,    -7,    -6,     4,    -9,   -28,   -34,   -23,     2,    25,    21,    -7,    -6,   -20,    -3,    13,     0,   -15,   -28,     4,    -3,   -16,     4,     7,   -11,     3,   -15,     1,    -9,    -3,     1,     9,    11,   -12,   -15,    -6,     9,    -1,    20,    -7,   -11,   -34,   -10,   -12,   -23,   -20,   -23,    -4,     2,   -17,     6,   -12,    13,    12,     8,   -11,    -1,    10,    17,    -3,    -2,    16,    19,    14,   -15,     4,    11,    11,   -34,   -22,   -14,   -10,   -23,   -27,   -18,     3,    -2,   -14,    -1,   -12,    -8,     7,    15,    -3,    14,    11,    12,    28,    15,     3,    -1,    -1,   -29,   -20,     6,     6,   -10,   -10,     7,     2,   -31,   -19,    -8,    -5,    -9,    -7,    -4,     6,    -4,   -25,   -27,     7,   -16,     1,   -18,   -23,   -18,   -17,   -29,   -28,   -29,    -9,    25,     5,    -8,   -10,     7,    37,     3,   -33,     0,     3,    -3,   -17,    -4,     4,    -4,    -7,   -28,   -47,   -48,   -18,   -13,   -25,   -24,   -35,   -35,   -44,   -24,   -14,    18,     3,     0,   -12,     3,    22,   -17,   -41,    -1,    -5,     0,   -18,    12,    -5,    -8,    -9,   -13,   -29,   -37,   -11,    15,    -6,    12,    -5,   -24,   -11,   -23,    -2,     5,    10,    -4,     4,     1,    15,   -28,   -19,    -5,     3,    -4,    -1,    19,     6,     4,    -9,   -12,   -18,   -19,   -13,   -14,     2,     8,     2,    -5,   -18,   -12,    -6,   -11,     9,     3,    -5,    25,    30,   -22,   -15,    -1,     3,     2,   -15,    -1,    -5,     1,    -8,   -11,   -13,   -27,   -17,   -21,     1,     0,     2,   -13,    -7,    -1,    10,    21,    38,     7,    28,    45,     9,    10,     1,    -5,     1,    -2,    15,    -9,   -11,     6,    -4,   -14,   -19,   -17,    -4,     5,    -1,     6,   -28,   -33,   -35,   -27,    -6,    22,    13,     9,    -3,   -17,   -14,     2,    -7,     3,     2,     5,     3,    10,    -1,     2,    11,     5,     6,     2,     0,   -12,    -8,     9,     9,    -9,   -25,   -20,   -25,   -22,     1,     3,    11,    23,    16,    -3,    -1,     2,     0,    -4,    -5,    -3,    -6,    -9,     5,    -2,     3,    -2,    -4,    -1,     8,    10,    11,    -1,   -13,   -14,    11,     7,   -12,   -26,    -2,   -14,     3,     3,     0,    -3),
		    40 => (   -5,    -1,     0,    -4,    -3,     2,     2,    -2,    -5,    -1,     3,    -3,     5,    -1,    -2,    -1,     0,     3,    -3,     1,    -2,     0,     2,     4,     2,     2,    -2,     0,    -3,     1,     2,    -1,     2,     2,     5,    -1,    -1,    -4,    -8,     3,    10,    -2,    -3,     7,    14,    14,     0,     0,     5,     2,    -1,     4,    -5,    -3,    -2,     0,    -2,     1,     5,    13,    10,    -2,     1,     3,   -14,   -28,   -24,   -15,   -26,   -39,   -31,   -38,    -9,   -18,   -15,   -24,   -23,    -5,   -22,   -12,    -8,    -4,    -2,     2,     2,    -3,    -5,     8,     1,    -7,   -18,    -7,   -10,     0,    -3,   -13,   -11,     0,     0,    -6,   -10,   -19,   -35,   -41,    -9,   -11,   -24,   -19,   -14,    -5,   -17,     0,     5,    -1,    -3,    -8,    -2,   -29,   -25,   -12,    -9,    15,    -2,   -11,   -26,    -2,     0,    -7,     7,   -18,   -23,   -14,   -16,   -11,    10,   -23,   -13,   -14,   -23,     0,    -1,     3,   -11,    11,    -3,   -13,    -4,     1,    15,   -11,    -4,   -14,   -14,     9,    -4,   -14,    -6,     7,    -1,   -18,   -26,   -18,    -5,   -17,   -10,   -13,   -20,   -18,     4,     2,    -8,    -8,    17,    14,     5,     3,   -30,   -26,    -2,   -10,   -12,    11,    -9,   -16,     5,     8,   -17,    13,    -3,    17,     6,   -31,   -16,   -35,   -18,    -9,     4,    -1,    -8,   -11,    17,    17,     4,   -12,   -36,     4,    -6,   -14,     0,    -8,    -2,     1,     7,    18,    29,    27,     6,     8,     5,    12,   -23,   -13,   -36,    12,    30,   -16,    20,     1,    12,     9,    -9,     2,    -2,    -1,    -8,    -9,    25,     0,    12,     8,    13,    16,    23,   -17,     2,    12,     6,    18,   -30,   -41,   -33,    -5,    -2,    -6,    22,    -1,   -28,    -2,    -6,   -11,     7,     2,   -15,   -14,     1,    -9,    11,    -1,   -18,     6,    12,    -7,    29,    -9,    -1,    -5,     2,   -43,   -37,     0,    -2,    -2,    22,     0,   -18,   -23,     0,   -11,    -4,    -5,   -17,   -26,     3,     1,    16,    -1,    -6,     7,    -2,   -11,    23,    14,    25,    -5,     0,   -28,   -35,     0,    -4,    47,   -16,    -4,   -21,   -26,    17,    24,     7,     9,    -6,    -5,     5,    -6,     5,   -13,   -15,     5,   -19,    -8,    13,    22,    17,   -17,   -18,   -29,   -28,    -2,     3,     7,    -6,    -7,   -20,   -17,    28,    20,    10,    11,    -2,     6,     3,   -12,   -20,   -17,   -35,   -23,    -8,    -7,    10,    24,     7,     4,    -3,    -7,   -31,     2,     1,     9,    11,    15,    -9,     8,    20,    21,    33,    13,    -5,     5,   -26,   -22,    -9,   -41,   -29,   -34,    10,     2,     5,    17,    21,    16,     4,    17,   -17,    -5,    -1,     4,    -3,     6,     6,    31,    25,    44,    26,    10,     2,     6,    -9,    -4,   -22,   -26,   -40,   -18,    -5,    15,    10,     1,     2,    24,    -6,    -3,   -25,     3,    -2,     1,   -10,   -12,    -2,    20,     1,    18,    39,    16,    -3,    -3,   -11,   -15,   -25,   -27,   -12,   -28,    -6,     0,    14,    25,    18,    34,    24,     5,   -39,   -10,    -2,    -4,    -9,   -18,    16,    -2,    20,    29,    11,     7,     9,   -13,   -21,   -21,   -30,   -26,    -2,    -6,     7,   -18,    -9,    22,    14,     0,    13,   -14,   -43,    27,    -3,    -4,   -12,   -30,     6,   -12,    -3,     3,    17,    22,    -1,   -23,   -38,   -26,    -9,    14,    -1,    -7,   -19,   -15,     7,   -19,    26,    -9,     8,   -21,   -32,    31,     5,     4,    -9,   -30,    -8,   -25,    -6,    17,    40,    23,     8,   -19,   -38,   -19,    13,     6,     0,    -7,     0,    -3,     8,     1,    15,   -16,    -2,    -1,   -19,   -13,     3,    14,   -14,   -12,    -8,   -18,   -13,    -7,    35,    14,     8,   -29,   -13,   -17,   -14,    -7,     2,   -12,    -4,   -20,    26,    -5,    12,    -4,    -2,   -37,    -3,    -3,    -1,    11,   -24,     1,    -5,     4,    -8,    -5,    14,    22,    41,   -15,    -1,   -12,    -9,   -18,   -14,   -11,   -16,    -7,   -22,   -16,   -10,   -30,   -27,   -20,    10,     4,    -1,    -5,   -33,   -15,    -8,     0,   -15,   -17,     8,    -6,    -2,   -14,   -17,   -21,   -16,     0,     9,   -11,   -31,   -22,   -17,   -11,    19,    -9,   -17,   -15,    16,     8,     2,    -4,   -31,    -7,   -29,    -6,     3,     3,    21,    18,    14,   -17,    -7,    -7,    -9,    -4,   -20,   -26,   -20,    -2,   -16,     4,     6,   -10,   -11,     3,    16,    10,     0,     5,    -3,   -35,   -27,   -19,     2,     2,    -3,     9,    11,    14,   -10,     1,   -11,   -11,   -13,   -16,   -32,   -16,   -31,    -8,   -20,   -19,   -21,    -7,   -15,    -2,    -5,    -4,    -5,     3,     3,    14,   -17,   -20,    -4,    20,    14,    14,    15,   -13,    -5,     7,   -18,   -31,   -20,   -21,   -18,   -21,   -28,   -22,    -4,     9,     0,    -3,    -4,     4,    -5,    -3,   -26,   -40,   -34,   -27,   -27,   -25,   -37,   -37,   -44,   -21,   -19,   -50,   -50,   -45,   -55,   -37,   -30,   -23,   -21,   -11,    -7,     2,    -1,     1,     2,     3,    -2,    -1,   -11,   -15,   -37,   -18,   -18,   -31,   -35,   -40,   -27,   -26,   -22,   -28,   -21,   -39,   -38,   -24,   -31,   -27,   -12,   -15,     1,    -2,     2,    -5,    -3,    -2,    -2,    -3,     4,    -4,    -5,     3,     1,    -2,     1,     2,    -4,   -17,    -7,   -10,    -9,    -8,    -4,     2,     1,   -16,   -10,    -9,    -2,     1,     2,     2),
		    41 => (    5,    -1,     1,     5,    -5,     0,    -3,    -1,    -5,     1,     2,     2,    -1,     1,     0,     5,    -2,     4,    -3,    -2,    -4,     5,     4,     3,    -5,    -1,    -2,    -4,     0,    -4,    -1,    -2,     4,    -3,    -3,    -4,     4,     0,    -6,    -5,   -10,   -13,     5,    11,     1,   -10,    -3,     3,     3,     1,     3,    -3,    -2,    -5,    -4,     0,     0,    -4,     4,    -4,    -1,    -4,     2,    -1,    -8,    -9,   -14,   -10,   -11,    26,    32,    43,    37,    21,    22,    43,    31,   -27,   -30,   -20,     2,     4,     0,     4,     4,    -3,    16,    30,    -2,   -14,   -23,    19,    13,    -5,   -41,   -41,     2,     4,     6,    18,    37,    17,    16,    20,    31,    28,   -16,   -19,   -10,    -7,     4,     4,     5,     2,     3,    19,     1,     6,    -9,   -24,   -19,   -10,     5,   -11,   -27,   -31,     6,    28,    28,    11,    21,     7,     8,    18,   -16,   -13,    -8,   -22,   -20,   -16,    -5,    -1,    14,    12,     3,    24,     9,   -26,   -18,   -19,    -9,   -10,   -30,   -15,    -5,    16,    26,     7,    -1,   -10,   -11,    16,   -17,    -4,    -9,   -19,   -18,    -9,    -3,    -2,   -20,     2,     2,     7,   -19,   -23,   -13,   -14,   -21,   -21,    -8,     5,     5,    16,    23,    -6,    -5,   -14,    -5,   -12,   -11,     2,     3,     0,   -14,   -11,    -3,    -7,   -27,    -7,   -13,   -33,   -36,    -5,    13,    11,   -12,     3,     2,   -11,    22,     5,     3,     6,   -43,   -24,    -5,   -16,   -22,    -8,    -2,    -1,   -18,   -18,    -4,    -9,   -25,     1,   -14,   -36,   -19,   -15,     7,    47,    -4,   -13,    -9,    -8,     9,    14,    -3,   -10,    -6,   -24,    -3,   -14,   -13,   -10,    -8,    -4,   -17,    -9,    -1,     0,   -29,    -6,   -13,   -20,    -2,     6,    22,    16,     7,   -16,   -17,    -7,     9,    16,    13,   -35,   -15,   -38,   -19,   -21,    -9,   -12,    -8,    -8,    -6,   -13,     5,    -1,   -31,    -4,   -21,   -32,   -18,    18,   -15,   -16,    -8,    -3,     0,   -14,     0,    -3,     0,     0,   -17,   -17,   -18,   -21,    -7,    -4,    -5,    -9,   -12,    15,    -1,     6,     3,    -3,   -12,   -17,     1,   -10,   -29,     4,    20,    -2,    -1,   -23,     1,    -3,    -6,   -17,   -37,   -20,   -21,   -10,   -14,    -3,   -13,    -6,   -19,     3,    -2,     4,    -2,    -4,    -3,    -9,   -10,   -17,   -21,    15,     0,    18,   -13,   -37,    -2,     1,     5,   -29,   -15,   -30,   -18,    -6,   -10,    -3,    -2,    -4,     3,     3,    -2,     3,     4,     0,   -16,    -9,    -8,   -17,    -7,    22,     5,    -3,    -9,   -64,     3,    10,     1,   -13,   -47,   -29,   -17,   -22,   -14,   -30,   -23,    -2,    -2,    -3,     1,     3,    -1,    -3,   -15,   -19,   -25,   -30,    21,    14,     5,   -24,   -65,   -33,    17,     2,   -11,   -30,   -44,   -35,   -30,   -24,   -23,   -21,    -5,    -8,     9,     2,    -4,     0,     5,     5,   -23,   -27,   -33,   -25,    24,    15,   -18,   -38,   -49,     5,     6,    -4,    -1,   -37,   -47,   -40,   -32,   -18,   -18,   -26,   -18,    -8,    -3,   -12,    -2,     3,     1,   -11,   -17,   -25,   -19,   -13,   -11,    -9,   -58,   -45,   -67,    -5,   -15,   -19,   -30,   -47,   -59,   -39,   -27,   -20,   -15,   -36,     9,   -18,   -23,    -9,     3,     2,    -4,   -17,    -3,     8,    29,    -7,   -19,   -15,    -6,   -37,   -47,   -16,    -3,   -22,   -15,   -26,     3,    20,     8,     2,    -4,   -32,     2,   -42,   -11,   -14,    -3,    -1,    -4,    -4,   -12,    28,    -2,    -8,    11,    -9,    -2,   -41,   -48,   -12,     2,    -5,     8,     0,     4,    14,    24,     3,    -8,    -8,     1,   -14,   -25,    -3,     2,    -4,     5,    -8,   -19,    -7,     2,     1,    11,    11,    -6,   -10,   -26,    -7,     0,     4,    24,     3,    -9,    14,    21,    -6,     3,    12,    -3,   -19,   -22,   -16,     0,    -2,     4,    22,    21,   -51,    -8,   -19,    -4,    42,     8,    -4,     1,    12,    16,    12,    24,    10,    28,    22,    15,     9,    35,    18,     2,   -10,    -8,     5,    15,    14,    -6,    33,    29,    15,    -6,    13,    14,    18,    27,   -16,    -7,    14,    -5,    -2,     5,    -6,    11,     4,    17,    22,     1,    -9,     7,    11,   -14,    -1,    10,     9,   -14,    19,    12,    43,    28,     4,    10,    10,     0,    -3,     3,    -2,   -24,    -1,    -2,    -4,    -3,     0,    11,    17,    15,    21,    24,    22,     9,    -2,     4,    -1,     2,    -6,    -1,    13,    32,   -15,   -26,     9,     2,   -12,     1,    -4,     4,     7,    -1,    -7,   -28,   -69,   -57,   -42,   -11,   -20,   -21,   -20,    12,     3,     0,    -5,     1,    -7,    -6,   -15,   -10,   -13,    -8,    10,     7,    -7,     4,    -1,     7,     1,   -24,   -32,   -20,   -36,   -20,    -1,   -17,   -16,   -30,    -7,     6,     3,     2,     2,     0,    -1,     2,    -1,    -5,     1,     7,     9,    -4,     0,    -5,   -32,     3,     8,   -19,   -60,     0,    -9,   -18,   -22,   -19,   -13,    -1,     2,     3,     3,     5,     0,     1,     3,   -10,   -16,    -6,    -4,   -13,   -15,    -2,     0,   -33,   -32,     4,    14,    16,   -19,    -4,     3,     1,    -6,    -5,     4,     4,     0,    -1,    -3,     2,     3,     3,     4,     1,    -2,    -1,     0,     5,    -4,   -13,   -12,    -4,   -10,     3,   -10,   -15,    -2,    -3,     0,    -1,     4,     2,     5,    -5,    -3,     0,     5),
		    42 => (   -5,    -4,     3,     2,    -3,    -2,     2,    -4,     4,     1,    -2,     2,    -5,    -7,     5,     8,     1,     3,    -1,    -5,    -2,     1,     0,    -2,    -4,    -1,    -2,    -3,     2,    -3,    -2,     5,    -2,    -3,     0,     0,     5,     0,   -12,   -10,    -9,     2,   -11,   -13,     4,     1,    -5,   -34,   -11,    -9,    -8,     1,    -5,    -3,     0,     0,     5,    -1,    -3,   -12,    -7,    -1,    -1,    -6,    -4,    -1,    23,    26,     2,     7,    13,    14,    23,    27,     9,    -3,    -1,    -8,   -12,    -7,     3,     3,    -4,     1,    -4,     3,    -2,   -19,   -22,   -11,    -4,   -13,    11,    13,    30,     1,    -7,    -3,    -9,    -4,     5,    25,   -19,    -3,    -4,    14,    -2,   -13,    -6,    -9,    -2,     3,     0,    -4,    -9,   -16,     0,    -6,    -9,    -3,    21,    42,    18,    -1,    20,    -7,    -9,    -3,    14,     7,     8,    -6,   -24,   -16,    -5,   -18,   -21,   -14,   -33,   -17,    -3,     0,    -6,    -1,    -5,     1,     6,    12,     2,     4,    13,    32,    10,    24,    23,    12,    23,    -7,    -6,    14,     9,    -1,   -21,   -19,   -17,    -6,   -43,   -16,     3,     2,     8,   -13,    -6,    14,    16,    27,    12,     7,    12,     7,    -4,   -10,     7,    15,    20,     8,    21,     0,     9,    20,   -12,   -46,   -47,    -4,   -35,    -6,     3,    -1,    15,    -9,    -5,    11,    15,    21,    10,     4,   -10,    -7,    18,    14,    -2,    16,    15,     7,     0,   -11,    -7,     5,   -22,   -27,     3,    20,   -53,   -22,   -13,    19,    19,    -6,    -2,     4,     9,     4,   -10,    -3,   -12,     8,   -10,   -10,    -8,   -19,     5,   -11,   -15,    -8,   -26,   -12,    -5,    29,    15,    -7,   -37,   -22,     3,   -22,    22,     6,     2,     3,     5,     1,     2,    12,    16,     1,   -13,   -16,   -20,    -8,    -9,    -4,   -26,   -21,    -9,     5,    -8,    18,    -4,   -29,   -13,    -9,    -5,    -9,    25,     0,     8,     2,    -2,    -3,   -12,    -3,     4,     8,    28,    -3,    -7,    -2,    -3,     7,   -19,   -16,   -13,   -10,   -24,   -22,   -10,   -17,    -8,   -18,     0,   -12,    -7,   -15,    -1,     7,     2,    -7,    -5,   -20,     1,     7,    15,   -18,     0,    10,     1,    -8,   -27,    -4,     7,     0,   -14,     5,   -11,    13,   -22,   -28,     3,   -12,   -30,    -9,     1,    -3,     3,   -11,    13,    30,    16,     9,    19,   -17,     4,     3,    -6,    -4,     0,    23,    -8,    14,    25,    18,    -3,    -3,    -1,     1,     0,    -6,   -15,   -19,    -4,    -1,    16,    15,    21,    10,     0,   -10,    -1,    -2,     1,    -9,     2,     9,    21,    27,    17,    18,    19,    10,    -9,   -14,    26,     2,    -2,   -15,    -5,    -3,   -22,   -25,     5,    35,    25,     5,   -13,    -6,   -14,   -17,   -24,   -12,   -10,     1,    33,    25,    16,    27,    31,    37,    31,     6,    20,    19,     4,   -11,    19,     6,   -19,   -11,     0,     8,    26,    11,   -15,     8,    -8,   -36,   -30,   -11,    -8,     5,     4,    27,    31,    23,    15,    24,     3,     4,     2,    17,     1,    -2,    21,   -14,   -20,   -20,    -7,    18,    13,    12,     7,    12,   -18,   -25,   -21,    19,     4,    10,    35,    36,    31,    40,    21,    48,    15,    19,    28,    14,    -1,    -2,    20,    -5,   -23,   -11,   -13,    -6,    18,    29,    26,    18,    11,    -7,     1,    11,   -15,    -1,    27,    44,    24,     9,     7,     7,    -8,   -15,    21,    15,    -1,    -1,     3,   -10,   -12,    -7,    -2,     3,    10,    23,    40,    18,    -3,    -8,   -15,    -7,    -2,    23,    38,    48,    37,    13,     6,    11,    12,   -22,   -10,    24,     3,    -7,   -15,    -2,    -6,    -1,    -4,     5,    11,    28,    21,    12,     9,   -27,    -2,     4,     2,    61,    66,    57,    22,    13,    18,     7,     6,   -23,    -1,    17,     0,   -10,     5,     7,     3,   -20,   -24,     2,    14,     4,    20,    15,    18,    -6,   -16,     9,    47,    42,    45,    31,    16,    -2,   -18,     3,    -6,    -5,   -12,     1,    -3,    -2,    15,     0,    24,    -7,   -25,     2,     0,   -11,   -10,     1,     0,     6,    -5,    33,    52,    47,    36,    37,    10,    -5,    -5,   -11,   -22,    -9,     2,     2,    -2,    -5,    -6,     2,   -11,     1,   -19,   -12,    -1,   -12,   -10,    -1,    21,    -3,    -6,    32,    69,    45,    59,    21,    13,    -5,    -5,    -9,     1,    16,    -1,    -3,     0,     3,    -3,    -3,   -11,    -2,   -10,     1,    13,   -13,   -39,   -25,    -1,     5,    26,    55,    74,    60,    47,    22,    -1,    14,   -17,    -2,    11,    12,   -18,     3,    -4,     3,   -13,   -18,   -54,   -53,   -16,   -12,    -3,   -36,   -29,   -18,   -15,    24,    35,    26,    53,    52,    38,    11,    -2,     0,   -12,    -7,    12,     1,     8,     4,     4,     4,    -2,    -9,   -21,   -35,    23,     7,    -6,   -14,     0,    26,    41,    49,    54,    50,    36,    17,    18,    10,    -6,   -11,   -32,    -3,     4,    12,     8,     0,    -3,     5,    -2,     0,    -9,   -26,   -38,   -35,   -35,   -38,   -42,   -21,   -30,   -27,   -37,   -27,   -27,   -26,   -23,   -32,   -13,   -12,   -39,    -1,    -3,    -2,     4,     3,    -4,     0,     3,     5,    -7,    -4,    -3,    -6,    -7,    -4,    -7,    -8,    -3,    -9,   -10,    -4,    -6,    -6,    -8,    -3,   -21,   -31,    -5,    -7,    -5,     3,    -4,    -3),
		    43 => (   -4,    -3,    -3,     1,    -2,    -2,    -1,     4,     5,     2,    -1,     1,    -1,     0,    -6,    -1,     2,     0,    -4,     2,     2,     1,     3,     3,    -3,     0,    -4,    -1,     2,    -1,    -2,    -1,    -5,    -3,     1,     1,    -4,    -3,    -9,   -11,    -8,   -18,   -14,   -32,   -43,   -48,   -18,    -5,    -1,    -4,     0,    -3,     5,    -1,    -1,     1,    -2,     3,     0,    -4,    -8,     2,   -10,   -17,   -33,   -32,    -7,     0,    -4,    -3,     0,    -1,     8,    -3,   -17,   -13,   -20,   -23,   -24,   -30,   -11,     0,     0,     0,     0,     0,     0,   -12,    -7,     6,    -2,     8,    20,    -7,     0,     8,    28,    -4,    -2,    29,    32,    23,    10,   -18,     3,   -14,   -23,   -53,   -43,   -18,     4,     0,     1,    23,   -35,     8,    10,   -11,   -23,   -26,     9,    17,    25,    -7,     1,     0,    -4,     4,    17,    -9,   -13,   -23,   -19,    -5,    26,   -25,   -52,   -47,   -12,    -1,    -1,     2,    -9,     7,   -10,    -2,     7,    10,    -4,     3,    -4,     3,    -3,    10,     4,     9,    15,    -8,   -30,    -3,    14,    -9,   -14,    26,    -6,   -55,   -19,    -2,    -3,     5,   -22,    -9,   -22,     2,    20,    15,     3,     4,    -5,   -23,   -24,     1,    12,    19,    14,    26,    16,    12,    11,    21,     8,     9,    33,   -50,   -42,   -20,     2,    -3,    -5,     4,     3,     1,     2,     8,    -1,    -3,   -14,    -8,    -4,     7,     9,     2,   -10,    17,    19,     7,   -10,     6,    -6,    41,    19,   -67,   -39,   -22,   -16,    -6,    11,    16,     5,     0,   -10,     5,    -4,   -10,     9,    -4,    19,    18,   -14,   -22,    -5,     7,    12,    25,     4,   -18,    19,    18,     3,   -74,   -48,    -3,     0,   -28,     0,    -9,    14,    -3,   -19,   -27,   -24,    -1,   -26,    -4,    46,    32,    12,     5,    16,     6,    -4,     6,    20,    -2,    30,    21,   -38,   -58,   -51,   -20,     2,   -28,     6,    10,   -14,   -16,   -31,   -33,   -37,   -39,   -45,   -10,    27,    41,    52,    17,   -14,    -8,   -16,   -11,     2,    11,     4,    10,   -38,   -24,   -38,   -20,    -2,   -15,    -5,    21,     3,   -18,   -45,   -41,   -18,   -30,   -57,   -12,     7,    42,    26,    23,     8,     3,    -3,   -15,    -9,   -15,   -20,   -38,   -96,   -48,   -31,    -5,     1,    -8,     3,     2,    -7,    -1,   -18,   -33,   -11,   -53,   -11,   -22,    10,    24,    60,    30,    -6,    12,    13,   -14,     0,    -9,   -58,   -67,   -70,   -35,   -26,    -5,     0,    -4,   -59,   -13,   -16,   -18,    -8,   -17,    -5,   -21,   -25,   -14,     4,    19,    41,    15,    37,     8,    10,     9,     5,   -17,   -40,   -17,   -41,   -42,   -28,    -5,    -6,    15,     2,   -34,   -37,   -25,   -16,   -20,   -17,    -7,   -29,    -8,    -1,    21,    16,    25,    10,    -1,   -22,   -18,   -20,   -27,   -14,     4,   -33,   -38,   -21,    -6,    -2,     8,     0,   -22,    -5,    -6,     7,    -4,     7,   -33,   -32,     8,    31,    32,    24,    31,    -8,   -32,   -37,   -17,   -10,    -4,    18,    18,    14,   -29,     5,   -15,     1,     3,     9,    18,     3,   -10,     0,     3,     0,   -15,    -5,    17,    12,     6,    24,    -9,   -38,   -22,   -10,    -5,   -19,   -17,    23,     4,    14,   -53,   -35,   -17,     1,     7,    13,    15,    10,   -20,    -8,    -8,   -25,   -17,    -3,    24,     3,    13,    -2,   -26,   -33,   -19,   -19,    -6,   -26,    -6,     3,     3,     2,   -42,    -9,   -14,   -11,     4,    16,    22,     0,    -6,     7,    16,   -13,    -7,    18,    30,     0,     1,   -12,   -15,   -10,     2,   -13,     4,     8,    13,   -11,   -12,   -22,   -36,    -7,   -20,    -1,   -15,    13,    37,    18,    26,   -14,    17,    -1,     9,    24,     7,   -21,   -14,   -29,     6,     5,    13,    13,     2,     9,     8,   -18,    -9,   -14,   -29,   -36,   -20,     1,   -15,   -26,     8,    -1,   -18,   -19,    11,    16,     5,    16,     8,   -26,    -8,    -9,    16,    17,     7,    -2,    -6,    -4,     8,   -11,    -2,   -18,   -24,    -6,    -1,    -4,    -6,   -16,     8,     2,   -29,     1,    19,    20,    -7,   -15,   -15,   -13,     4,    -7,     2,    -5,     1,    -2,     2,   -13,   -11,    -1,   -19,   -45,   -29,   -12,    -3,     1,     0,    -7,    10,   -19,   -12,    21,     1,   -18,   -10,    -7,    -8,    -3,     2,     0,    -1,    -5,     6,    -9,    -9,    -5,     4,    -1,   -32,   -39,   -53,    -4,    -1,     0,     2,    10,    30,    -7,     2,    25,     8,    16,     5,    23,    12,   -15,    13,   -18,     0,    17,    -2,    15,    -5,   -12,   -18,   -21,   -26,    27,     5,   -17,     4,     2,    -3,    12,    30,    -6,    -1,     8,     3,   -13,   -16,     2,    42,   -23,    -2,    29,    -7,    -7,   -14,     1,     2,    -3,    -5,   -13,   -13,   -28,   -25,   -10,     4,     4,     0,     4,   -15,   -18,   -15,   -24,     7,    11,     2,    35,    34,    52,    16,    -2,   -17,    14,     1,     6,    18,   -21,   -43,   -51,   -56,   -26,    -5,    -9,     2,    -2,     5,     1,   -16,   -35,   -17,   -19,    -9,    -4,   -10,    16,    10,    19,     4,   -30,   -17,    -3,     5,     8,   -16,   -14,   -30,   -40,   -27,    -1,     1,    -4,    -3,    -4,    -2,     3,     5,    -9,   -14,   -11,    -9,    -9,   -28,   -30,   -33,   -26,   -48,   -20,   -22,   -14,    -7,    -8,   -29,   -33,   -15,    -2,     5,    -2,     1,    -2,    -3),
		    44 => (    3,     3,     5,     4,    -4,    -3,     4,     5,     3,     5,     2,     1,     0,     0,    -4,    -3,     1,     0,    -2,     4,     0,     2,    -3,    -2,     4,     5,     2,     4,    -1,     2,     4,    -4,    -1,    -5,    -5,    -8,    -1,    -4,   -24,    -9,   -34,   -26,    -3,   -16,   -12,    -1,    -4,    -3,   -15,    -2,    -6,   -10,    -5,    -3,    -1,     4,    -3,    -5,    -5,   -25,   -27,   -30,   -12,   -22,   -18,   -17,    -7,   -31,     8,     3,   -15,   -37,   -24,   -19,   -19,    -7,    -9,   -11,   -16,    -3,    -2,    -4,     4,    -3,    -5,    -5,    -1,   -33,   -50,   -27,   -29,   -27,   -32,   -20,    16,   -12,   -30,   -61,   -37,    -4,    -9,    -3,   -26,   -27,    -6,    -8,   -20,   -11,     0,   -11,    -1,     4,    -5,     3,    -5,   -21,   -10,     7,     9,     2,    -6,    -1,   -27,   -45,    -5,     7,   -40,   -52,   -57,   -51,   -28,    -9,    -4,     1,     9,    15,    22,     7,   -14,    -7,    -1,     3,    -6,    -5,    -5,     1,    -9,    -8,   -28,   -44,   -35,     3,    28,   -10,   -20,    -7,   -24,   -96,   -51,     5,    23,     8,     2,     2,     1,    -1,   -13,    -9,    -4,    -1,    -1,   -19,    15,    49,    -6,   -31,   -18,   -14,   -23,     8,    22,     7,   -17,   -18,   -69,   -75,   -31,    22,    16,     6,     1,    16,    21,   -47,    15,   -40,    -1,   -34,    -3,   -16,     6,    41,   -21,   -12,    -9,    -4,     7,    13,    -1,    14,    -6,   -37,   -81,   -76,    -5,    26,    12,    -8,     2,    11,    -9,   -12,    16,   -42,   -14,   -30,     7,   -10,     0,    10,   -16,     8,   -17,     0,   -14,    -3,    14,    12,     4,   -39,   -98,   -30,    13,    13,     7,    -7,    19,   -19,     1,    27,    12,   -26,     3,   -25,     3,   -14,    -6,     7,   -13,   -10,   -11,     4,    -2,     3,    24,    25,    17,   -49,   -51,    13,    25,     9,    13,     7,    11,     8,    27,   -25,   -24,   -17,     4,   -16,   -23,     7,    15,    24,     1,   -13,    -2,     8,    -9,    -7,    -3,    32,   -12,   -54,   -36,     8,    25,    21,     3,    -4,    10,    17,     8,   -46,   -15,    -3,    -5,   -10,   -13,   -31,   -14,    10,    25,    -5,    11,   -10,     6,    -2,    24,   -11,   -37,   -54,   -32,   -12,     4,     5,   -23,    17,     0,    -5,    18,   -23,   -22,   -18,    -3,    -1,   -24,   -30,   -41,   -13,     6,    20,    16,   -16,    -6,    16,    21,    13,   -45,   -25,    -6,    -5,    -7,    16,     0,    23,     5,    18,   -27,   -24,   -47,   -27,     3,    -7,   -26,   -29,   -35,   -19,    -5,    -6,    10,    10,    17,    23,     6,     7,     2,     6,     8,    16,   -13,    16,    14,     9,    -3,   -10,   -47,   -38,   -37,    -1,    -3,    -4,    -6,   -31,   -24,    -3,    -4,     1,    -5,    14,     4,    15,     3,    -7,    16,     4,    -2,     2,    -8,    14,     6,   -11,   -13,    -7,   -22,   -26,   -30,     0,    -1,    -1,    -4,     9,    -1,     0,     1,    -5,    13,     4,    14,    11,     0,     6,    10,     2,    -8,    -4,     1,    26,   -49,   -15,    -8,    -5,   -23,   -36,   -25,    -1,    -2,    -4,   -12,     8,    -1,    -8,   -33,    -3,     3,     3,     1,    -1,    -5,     0,   -13,     2,    -6,    -9,    -8,   -11,   -36,   -19,   -11,   -19,   -28,   -39,   -39,    -8,    -2,     1,   -16,     7,    21,    -3,   -24,   -11,   -16,    -8,    -8,    -7,    -1,     1,    -7,     2,   -13,     7,    -6,   -26,   -40,     7,    -7,    -8,   -30,     3,    -7,   -10,   -18,     3,   -21,    34,    45,   -19,   -12,   -25,   -19,   -23,   -45,    -1,   -16,     3,     5,    -4,     5,   -21,     0,    -9,     3,    19,     9,     9,     0,    17,    -2,    -4,    -1,   -22,   -10,    28,    14,   -21,   -27,   -17,    -9,   -24,   -26,    -6,   -21,     2,    -4,   -13,    -3,     4,    -9,   -10,    -6,     8,     5,     8,    18,    11,    -5,    -9,     5,     1,    -8,   -34,   -31,   -37,   -33,   -20,   -25,     0,   -14,   -15,   -20,    -1,    -7,   -12,     6,    -3,   -12,   -12,   -33,   -29,   -19,   -10,   -31,   -45,    -8,     2,     2,     0,    -8,   -20,   -34,    40,    -3,     6,    26,    33,    -9,    -4,     2,    -3,   -10,    -7,    -5,   -34,   -29,     4,     4,    -4,     4,    13,   -17,   -60,   -20,    -5,    -4,     5,     2,   -22,   -38,    22,    25,    16,    14,     1,    16,     1,     0,    -1,   -13,    -7,     2,   -15,   -26,   -11,     0,     4,    -2,    16,   -19,   -18,     9,     4,     3,     2,    -1,   -21,   -33,   -63,    10,    16,    13,    11,     8,    -1,    10,    -6,     6,     7,    20,   -14,   -13,    -7,    -5,    10,     5,    11,   -12,     4,    12,     4,     2,     3,    -2,    -7,   -49,   -42,    -7,   -21,     0,     7,    11,    -7,     4,     0,    -2,    19,     9,   -22,   -53,   -12,   -10,    14,     7,    15,   -20,    21,   -15,    -4,     4,    -4,    -8,    -3,    -1,   -30,   -26,     1,    -4,   -16,     1,     4,     8,    14,     1,   -19,   -21,   -45,   -27,   -19,    -5,    -8,    13,    28,    -6,   -13,    -3,     0,     2,    -3,    -1,   -25,     2,   -27,   -26,   -43,   -21,   -27,   -28,   -20,   -37,   -52,   -59,   -79,   -17,   -22,   -33,   -16,   -20,   -21,   -16,    11,     1,    -4,    -2,    -2,    -1,    -2,     0,     3,     4,     0,   -14,   -20,   -17,   -13,   -28,   -33,    -4,   -18,   -28,    -2,   -22,   -30,   -16,   -14,     2,    -5,     3,     0,    -2,     5,     3,     2),
		    45 => (   -1,    -4,    -2,     0,    -4,    -5,    -1,    -4,     5,    -5,     2,     4,     3,    -3,    -5,     2,    -5,    -3,     3,     3,     1,    -3,    -2,     0,    -2,    -2,     4,    -3,     0,     0,     2,     0,    -1,    -3,    -4,    -1,     3,     1,    -4,    -9,    -9,    -9,   -13,   -20,   -22,   -17,   -25,   -24,   -24,   -19,    -3,     1,     2,    -1,    -5,     4,    -3,    -3,    -9,   -10,   -11,    -3,    -5,    -4,   -26,    -6,   -14,   -10,   -19,   -25,   -26,   -23,    -7,   -13,   -16,   -17,   -14,   -21,   -19,    12,   -34,    -5,    -1,    -4,     5,    -1,    -5,    21,    46,    -8,   -20,   -22,    -7,    10,    -7,   -31,   -25,   -41,   -34,   -16,    12,     2,     3,    -3,     2,     8,   -32,   -27,     1,    39,    35,     2,     2,     4,   -14,    37,    -2,    -2,   -22,   -19,   -18,    -4,    -2,   -36,   -39,   -27,   -21,   -14,   -27,   -24,    -2,    25,    -2,     0,   -24,     2,    31,    26,     3,   -11,     3,     0,   -26,    41,   -10,    -8,   -13,   -25,   -22,   -11,     2,     1,   -32,   -13,   -11,    -7,   -15,    -5,    -4,    17,     4,    -5,   -13,    -8,   -12,     9,    -2,   -10,    -2,    -1,   -20,    -7,   -13,    -9,   -15,   -26,   -13,    -3,    -5,   -23,    -2,     3,    -5,     1,    -3,   -19,    -1,   -10,   -11,   -20,    32,    24,    15,    32,    35,     2,     1,    -6,     4,   -11,    -8,   -19,   -14,   -18,     4,    -7,    -1,    -3,    12,    14,    15,     7,    17,    22,    -4,   -17,    -1,    12,    11,    13,     9,    -2,    41,     9,   -12,    -4,   -21,    -6,   -11,   -17,   -10,    -8,    -7,     1,     1,    -6,    -7,     1,    13,    -4,    -6,     5,     4,    37,    42,    20,    29,    24,     8,    -6,    15,    20,     5,    -9,   -41,   -29,   -13,   -14,   -20,   -11,    -7,   -13,   -14,    -2,    10,    -1,     8,     0,    -3,     6,   -10,   -22,    13,     5,    12,    20,    53,    42,     9,    10,     0,    -3,   -18,   -21,   -22,    11,   -10,    -1,     4,   -13,   -15,    -2,    17,    -3,    -2,     7,    17,   -23,   -82,   -87,   -47,   -41,   -44,   -15,    -1,    11,     5,    16,     0,     3,     0,    17,     9,    10,    -8,    -9,   -19,   -35,    -7,   -23,   -26,   -17,     2,    -4,     4,    -6,   -43,   -50,   -75,   -69,   -70,   -55,   -44,   -10,    -2,   -10,     3,     0,    -1,    22,    10,    -4,   -26,   -35,   -30,   -23,    -7,   -22,   -30,    -1,    14,    -6,   -11,     8,     1,    -8,   -32,   -58,   -51,   -90,   -58,   -29,    -5,   -17,    -2,    -4,     0,    28,    -3,   -13,    -8,   -12,   -17,    -1,   -10,     0,    20,     4,     8,     9,    -5,     6,    13,    26,    16,    17,    -2,   -33,   -47,   -14,     2,   -19,     6,     0,    -7,    17,   -20,   -29,    -3,   -19,   -24,    -6,    -1,    11,    -4,     2,     4,    18,    15,   -16,     0,     9,    24,    -7,     0,    21,    11,   -14,    -8,   -16,     5,    -2,   -18,     3,   -16,     0,    12,    -4,   -10,   -27,    -8,   -12,   -12,    14,     2,   -20,   -12,    -3,   -11,    -8,    24,    -3,    -6,    18,    32,    -1,    -2,    -3,    -4,   -14,   -37,     2,     5,   -25,    26,     6,     3,   -38,   -32,   -35,   -21,    -7,    -3,   -14,    12,     8,    -1,    -1,    29,    21,     1,   -15,     4,    13,    -7,    -8,    -4,   -15,   -45,   -16,    19,    -5,    22,    43,    17,     2,     4,   -24,   -44,   -20,   -23,   -20,     0,     0,    -4,   -13,    17,     0,   -36,   -28,    -6,    -6,   -14,    -9,    -4,    -2,   -35,    -3,     5,     8,    13,    33,    20,     4,     7,   -11,    -1,   -13,    -1,    -1,    -3,     3,   -13,   -17,   -12,    -8,   -19,   -37,   -23,   -11,   -28,   -25,     3,    -7,    29,   -32,   -11,    -6,    15,    27,    19,    28,    13,    21,    20,    15,     7,    -3,    -7,   -13,     7,    12,    -9,   -15,   -17,   -25,   -15,   -12,   -16,   -19,     4,    -6,    24,   -42,   -28,    -2,    -1,   -18,     7,    10,    15,    11,    10,    -2,     4,     0,    -4,    -2,    -2,   -10,    -7,   -15,    -8,    -8,    -8,    -7,    -5,    -4,    -4,     1,   -14,     1,   -18,    12,   -10,    -3,   -26,   -18,   -12,    10,   -11,    -6,     8,     0,     7,     6,     6,   -11,   -19,    -1,    -3,    -7,    -8,    -7,    -5,    -4,    -2,    -2,   -40,    12,    16,    -2,   -21,     2,   -26,   -12,   -10,    -4,     0,    -8,     6,     4,     1,     1,    -1,   -16,    -1,    11,     4,    -3,    -6,    -5,    -3,     3,     2,    -3,     5,     7,    24,    31,     3,   -16,   -21,   -20,    -2,    -3,   -19,   -25,    -3,   -11,     0,    14,    17,     2,    -1,    11,     7,    -2,   -17,    -8,    -6,    -5,    -3,     1,   -19,     0,    -6,    -7,   -23,   -42,   -36,   -14,   -42,   -51,   -18,    -5,   -14,   -20,   -27,   -17,     3,    15,    12,    -1,    10,     2,     6,   -24,    -9,    -2,     2,     5,     0,     9,   -17,   -11,     1,   -10,   -26,    -7,   -46,   -44,     4,   -12,   -13,    -6,    -1,    -7,    -4,    -4,    -5,   -16,     7,     1,     5,     3,    -5,    -3,     4,     4,     5,    -6,    -8,   -11,   -17,   -10,   -13,   -11,    -7,   -11,    -8,    17,    36,    34,    28,    14,    -2,    20,     2,    -9,     1,    -4,    -4,     4,     3,     0,    -1,    -4,     4,     4,    -1,    -7,    -3,     1,    -3,     1,     3,    -1,    -1,     1,    -3,    -1,     0,     1,    -9,    -9,    -8,    -8,   -26,    -5,    -1,    -1,     3,    -4),
		    46 => (   -3,     2,    -4,    -1,    -5,    -3,     0,    -3,    -5,     0,     4,    -1,     1,     3,    -4,     3,     1,     1,    -3,     4,    -2,    -4,    -4,    -4,     4,     0,     3,     3,    -2,     3,    -1,    -3,    -1,    -1,    13,    19,    26,    28,    14,     9,     3,     9,     9,     3,     1,    -3,     6,     7,    34,    11,     6,    10,    -2,     2,    -2,     1,     0,    -2,     4,     3,     6,     2,    21,    28,    29,    15,    -9,    -8,    -8,    -1,    -4,    -3,    -5,   -13,    -4,    17,    16,     5,     6,    17,    16,     5,    -4,     0,     2,    -2,   -23,   -16,     1,     4,    13,    21,     9,    15,     2,   -21,   -24,    -8,    -3,    -3,    -2,    -5,    -5,     7,     1,    16,    -1,    18,    22,    -1,    -9,    -2,    -1,    -5,   -12,    -6,     2,     6,     5,     3,     4,     5,   -15,   -13,     0,   -13,    -7,    13,    10,     0,    -5,     0,    -3,     9,    -1,     8,     6,     2,    11,    14,    -4,     3,     4,    -9,     5,    -9,    -3,     5,     4,   -12,   -20,     3,    -2,   -12,     8,    -8,   -16,     5,     5,     3,     9,     0,     3,    11,    11,     3,    25,    15,     2,     0,     1,    -2,    -5,    -3,    -9,     4,     1,    -9,     4,    -4,     3,   -14,   -14,   -20,   -25,    -3,     5,     9,    13,    19,    13,     9,     0,   -15,     8,    10,    -2,     0,     4,    -8,    -2,    -6,   -13,   -14,     6,     4,     1,    -7,   -23,   -11,     9,     1,   -11,    -6,   -13,    -3,    -1,    -4,    -6,    -5,    10,    -9,     3,     6,     3,     3,    -3,   -17,    -6,     0,    -7,   -16,     7,     6,    -3,   -22,   -15,    -5,    -5,   -15,     7,    11,   -11,   -12,   -20,    -8,   -30,   -25,   -17,   -19,    -7,   -21,     2,     4,    -3,    -5,    -9,   -19,     1,     0,    14,     2,    -9,   -16,   -16,   -17,    -5,     7,     1,    -5,   -15,   -27,   -28,   -23,   -36,   -27,    -9,   -14,     3,    -5,    -1,    -1,     0,    -9,    -4,   -14,     0,    -7,    12,   -16,   -15,   -24,   -12,   -17,    -2,     9,    -2,   -21,   -24,   -13,   -23,   -17,   -24,   -26,    -9,    -9,    -7,   -12,     0,     1,    -3,    -3,    -2,     6,    15,    -1,     3,   -13,   -26,   -16,    -6,     0,    11,    -2,   -24,   -27,   -21,     0,     3,     0,    -6,    -7,     4,   -15,   -10,    -1,     3,    -2,    -1,    -2,   -14,     8,     3,    -8,    -4,   -11,   -24,   -10,    -9,     7,    -6,   -15,   -15,    11,     8,    -3,     6,    10,     8,     6,     7,   -19,   -23,    -5,    -3,     2,    -6,    -4,    -8,    13,    -5,     4,    11,   -19,   -23,   -13,     6,     6,   -18,    -6,     0,    -2,     7,     9,    -4,    -4,     0,    10,    14,   -14,   -13,     2,    -4,    -4,     3,    -3,    -6,    20,    -6,     5,     5,   -16,   -16,    17,    10,    -5,   -16,    -1,     4,    18,    17,    16,    -2,   -16,    -4,    11,    12,    -5,    -9,   -11,     1,     4,    -7,    -6,    -3,    11,    -4,    -1,    -1,    -6,   -17,    -4,    -9,   -21,    -8,     8,    16,    13,    16,    20,    -4,    -8,    -6,    15,    17,   -10,   -12,   -22,    -5,     3,    -5,   -10,    -3,     6,    -5,   -18,     5,   -10,   -10,    -7,   -18,    -5,     5,     4,     7,    16,     1,   -12,    -2,    -5,    -2,     1,     0,    -5,   -10,   -19,    -1,     3,    -9,    -2,    -1,   -15,     0,   -20,     6,    -2,    -6,   -28,   -25,    -3,     9,     2,    -2,     2,    -3,    -9,    13,    10,    -3,    -5,    -1,     2,    -7,   -20,    -1,    -2,    -9,    -1,    -5,   -13,   -21,   -11,    11,     8,    -6,   -15,    -8,     7,     0,     5,    -2,   -11,    -8,    -8,    14,    -1,     0,   -13,    -9,    -1,   -21,   -15,    -2,    -4,     1,     0,    -2,   -14,    -2,    -4,    -4,     2,   -12,     6,    -1,    -8,     5,   -12,    -1,   -10,    -2,    -8,    10,    -4,    -5,    -3,    -5,    -8,    -9,     0,     3,    -1,     2,   -11,     4,    -8,   -10,    -5,    -1,   -10,    10,    -3,   -15,   -11,     3,    -5,   -18,    -7,    -4,     3,    13,     7,   -10,   -15,    -5,     6,    -8,    -1,    -5,     5,    -1,    -7,     1,   -10,   -12,     3,    -5,     7,    -4,    -1,   -14,   -17,    -6,   -10,    -6,    -9,    -2,     5,     9,    -7,   -18,    -8,   -12,     3,    -4,     1,     0,    -2,     2,    -3,     0,    -2,     7,    -2,     1,    -7,    -1,   -11,    -5,    -8,   -13,    -1,     2,    -4,   -15,    -8,   -12,    -6,   -21,   -12,    -8,   -10,     6,    -3,    -3,     2,    -1,    -8,     3,     0,    -9,    -8,     6,     7,     4,     7,    13,   -12,    -7,   -12,     9,    -5,   -14,   -21,   -13,   -19,    -8,    -5,   -10,     2,    -7,     3,    -4,    -1,    -5,     1,    -6,     0,    -7,   -12,    -9,   -12,    -9,    -1,    -1,   -10,    -9,   -14,     1,     2,    -4,   -21,   -21,    -4,    -4,    -5,    -2,    -4,    -3,     4,     1,     1,     0,    -4,     3,    -2,    -9,    -6,    -4,     2,     1,    -1,     0,    -1,     0,    -1,    -5,    -7,     1,    -1,   -14,    -4,    -7,   -16,    -4,    -4,     3,     1,    -3,     3,    -2,    -1,    -1,    -4,    -3,    -6,     0,     2,     2,     0,     4,    -5,     2,     0,    -4,    -3,    -3,    -2,    -4,   -11,    -2,     2,     4,     3,     3,     2,     4,     4,     2,     4,     0,     2,     2,     1,     1,    -2,     1,    -5,     3,     2,    -4,    -4,    -1,     3,     3,     3,    -2,    -4,     1,     1,    -5,     2,     3,     3),
		    47 => (   -1,    -1,     2,    -5,     3,     1,    -3,     4,     1,     0,     0,     3,    -2,     2,    -4,    -1,     2,     1,     0,    -5,    -1,    -4,    -3,     3,    -3,    -1,     5,    -3,    -4,     0,     1,    -4,     4,     4,     4,     0,    -4,     4,    -4,   -27,   -19,   -23,    -7,    -4,   -10,    -8,     3,     2,     4,     2,     3,    -4,     0,    -4,     1,    -2,     4,    -5,    -1,    -3,    -2,    -5,    -2,    -1,     1,    -4,    -6,   -19,   -28,   -18,   -14,   -12,    -5,     2,     0,    -5,    -6,     1,    -6,    -1,    -5,     0,    -5,     4,     1,    -1,     5,   -10,   -10,    -5,    -8,   -17,   -14,    -9,     0,    -7,   -14,    -8,     1,   -21,   -22,   -13,    -9,    -3,    -8,    -2,   -18,    -4,    -6,     2,    -3,    -3,     3,    -3,     5,    -4,    -3,   -16,   -18,   -17,   -24,   -11,   -15,   -24,   -28,   -22,   -14,   -18,   -16,   -19,   -11,    -2,   -11,    -7,   -26,   -15,   -10,    -9,    -5,    -1,    -3,     4,    -3,   -14,   -10,   -26,   -32,   -21,    -6,    -6,   -25,    -4,     6,    -1,   -18,   -41,   -43,   -29,   -40,   -50,   -46,   -29,   -26,   -25,   -21,    -7,    -1,     5,    -4,     0,     3,     6,   -13,   -28,   -36,   -45,   -38,   -57,   -48,   -13,    17,    18,     6,   -15,   -28,     9,    14,     1,    10,    38,    10,    20,   -23,    -8,   -23,    -6,    -4,    21,    13,    20,     9,    -7,    20,    -1,   -18,   -50,   -45,   -43,   -33,    -8,    -6,   -26,    -1,     0,    10,   -16,   -31,   -16,   -13,    -8,    -6,     3,   -13,   -10,   -13,    24,   -10,    -2,    -4,     1,    20,    21,   -16,   -39,   -38,   -38,   -19,   -31,   -33,   -37,   -23,   -17,     7,   -17,   -20,   -32,   -12,    19,     9,     1,   -37,   -13,    -9,    22,   -12,   -11,    -1,     7,    33,    -3,     5,   -12,   -29,   -12,   -18,   -31,    -4,    -6,    -3,     2,     4,   -17,   -13,    28,    19,    39,    24,     8,   -24,     2,    -6,    13,     5,    -6,   -30,   -10,    14,     1,   -17,    -9,     0,    -3,     2,    15,     6,     0,    -8,    21,    13,    12,    -3,    19,    17,    -2,   -17,    -5,   -27,     8,    -2,     6,     4,     2,    -1,     5,    -9,    23,    -7,     0,    -3,    34,    23,    16,    17,     0,   -14,   -11,     3,    11,     7,    11,     7,    12,    -7,   -15,    -5,    31,     0,    -1,     9,    21,    17,    17,   -17,    19,    22,     1,     5,    22,    30,     6,   -16,   -17,    14,    22,     5,    -7,    -2,    -8,    16,    -2,    27,    20,    37,    37,     2,     7,    17,    22,    17,     7,     8,   -24,    -8,     3,    15,     5,     1,   -16,   -18,   -18,    11,    -6,    -5,    -3,    22,    13,    17,   -28,    27,    26,    15,    -7,    -7,    18,    31,    23,     6,    39,     2,   -27,    10,    13,    20,    -5,   -39,   -52,   -14,   -15,    -8,   -15,    19,     6,    13,    12,     8,     4,     2,    -9,   -22,    -4,     3,    -4,     1,    33,   -22,    11,    -5,    15,     0,    21,    20,   -20,   -63,   -54,   -30,    -4,    -2,    10,     0,    23,    18,    -3,    -6,   -31,   -26,    -6,    -2,     0,     2,    -5,    -3,    16,    37,     3,     6,     8,    -2,    -1,   -19,   -77,   -89,   -18,   -10,     0,    -4,     2,   -20,     7,    19,    13,     6,   -20,   -34,   -43,     2,   -18,     4,    -1,    19,    -1,    22,    -2,    -6,    -6,    -1,   -21,   -51,   -63,   -51,    -2,    -9,     5,   -16,    -6,   -11,   -16,    22,    15,     7,   -16,   -26,   -30,     4,   -26,    10,     3,    18,   -29,     1,    -7,     0,    15,    -4,   -43,   -64,   -29,   -17,     2,     7,     3,   -27,     0,   -10,   -10,    22,    11,     2,   -24,   -26,     1,     5,     0,    -1,    22,     4,   -32,    -7,    -2,    16,     5,   -15,   -47,   -54,   -19,   -10,    23,     1,    -6,    -3,    12,   -14,    10,    -5,   -13,   -10,   -25,   -23,     6,    -4,     2,    -2,     5,    -2,   -13,    -6,    -7,    -6,   -16,   -21,   -37,   -26,    -5,     6,     1,     5,   -11,   -20,     9,    -7,    -2,   -11,    -4,    -9,   -19,   -17,    -3,     0,    -2,     4,     5,    -1,   -23,   -27,   -18,   -30,   -43,   -23,   -19,     4,     9,    -4,     2,    -2,   -14,   -16,    -3,     9,     8,     1,     7,    -8,   -23,    31,     0,    -5,     3,     1,    -2,    -5,   -33,   -14,   -17,   -22,   -31,   -21,     2,    -7,     1,     7,    12,    -6,    10,    -9,   -17,     9,   -15,    23,    -9,     0,   -24,     5,     4,    -3,    -1,    -4,    -1,    -6,   -23,     0,     4,   -28,   -14,    -5,   -15,    12,     4,     5,    -1,     0,   -16,    -4,     2,    -9,     0,    11,   -19,    -4,   -23,    10,    -1,    -5,     4,    -1,     0,     0,     6,    13,     1,   -17,     2,    -3,    18,     0,    14,     8,   -25,    12,    -3,    -7,     0,   -14,   -27,    12,     5,    -8,   -29,     5,   -15,     3,     1,     1,     0,    -2,     2,    -7,    10,     9,     6,    -4,    -1,    11,    23,    16,     3,    27,    10,    18,    -1,    -7,     6,    -7,     6,     0,   -29,    10,    -6,     4,    -3,     0,     3,    -1,    -7,    -4,   -13,     3,   -15,     0,    -1,   -21,    -1,    30,    20,    -6,   -12,     2,     7,   -12,   -20,     2,    11,     7,     6,    -6,    -3,    -4,     2,    -4,    -4,     0,     1,     6,    12,    -6,     7,    19,    17,    -6,     1,     6,    16,    -7,   -12,     8,    21,   -25,    -5,    -1,    29,    29,    27,    -5,    -1,    -4,     3),
		    48 => (   -4,    -4,    -1,    -1,     1,     4,     2,    -4,    -3,    -2,    -1,     4,    -3,    -2,    -1,    -5,     3,    -5,     1,    -4,     3,     1,    -3,     2,     1,     2,     3,     4,     4,     0,    -1,     5,    -4,    -2,    -1,    -4,     0,    -4,     1,    -3,    -1,    -3,    -7,    -4,   -13,    -6,    -8,     0,     4,     0,    -5,    -3,     4,    -2,     2,    -2,     4,     4,     0,     2,     0,     0,    -2,    -5,   -16,   -18,   -27,   -21,     4,     2,     3,   -14,   -14,    -1,    -7,     3,   -20,   -17,   -16,    -8,   -11,    -4,     4,    -2,    -5,    -4,    -5,     1,    -8,   -14,   -22,   -19,   -13,   -14,   -16,     5,    15,    11,     4,   -10,    -1,    -6,    18,     6,     2,    -4,    -4,    33,     3,     4,    -8,     5,     4,    -3,     4,   -12,   -20,   -30,   -22,   -23,   -10,     4,    -8,    -5,   -13,   -19,     0,   -16,    -5,    -8,   -14,    17,    40,    45,    11,   -29,   -30,   -11,    13,    -4,     0,     1,   -11,    -7,   -26,   -14,   -12,    -4,    -4,   -13,    -9,     4,     1,   -16,    -1,   -39,   -29,   -20,   -27,     6,    24,    32,    15,   -12,   -20,    -8,     3,    -4,    -3,     0,   -10,   -34,    -5,   -13,    -4,     3,   -19,    -7,    -6,    -5,    -9,    -7,   -11,   -19,    -8,    -6,     3,    -8,    -7,    -2,    -4,   -10,   -24,   -15,     1,     6,     0,    -8,    -6,   -20,    -1,    -1,     0,    -5,    -2,   -12,   -13,   -18,   -24,     1,     2,     7,     4,   -13,    -1,    28,     3,     1,     8,    -6,   -24,   -12,     8,    13,     0,   -18,    -7,     9,     7,     7,     6,    -2,    -4,   -14,   -19,   -30,   -27,   -24,    -7,     7,   -11,    11,    -5,   -13,     4,    26,    22,    -3,   -17,     4,    10,    24,     0,   -11,   -16,    -9,     9,     0,     7,    10,    -5,     5,    -3,   -19,   -29,   -44,   -20,   -11,   -11,    -5,    -1,    -5,     2,    11,    -4,    -7,    -6,   -10,    -6,    -2,     4,   -11,   -20,   -20,     2,    12,     1,    -2,   -10,    12,    -6,    -8,   -25,   -30,   -14,    -5,    11,     8,    -6,    16,    20,     2,    -5,    -6,    -8,   -25,    -1,   -10,    -2,     1,   -12,    15,   -11,     1,     7,    -7,     3,    11,    12,    -6,    -5,     1,    -9,   -30,    -7,    20,    -5,     3,    10,    -5,   -18,   -17,   -24,   -15,    -2,    -9,     1,     4,   -13,   -12,    -8,    -3,   -11,   -13,   -24,    -6,     9,    25,     4,   -18,   -25,   -25,    -3,    11,   -11,    -8,     3,     0,   -12,     1,     3,    -8,   -14,   -12,     0,     0,   -15,   -14,   -24,    -8,    -7,    -3,     0,    11,     6,    24,    12,     7,   -22,   -19,     3,    -8,   -37,   -12,   -12,    -9,    -2,    -5,   -18,   -15,     3,    -4,    -4,    -5,   -10,   -20,   -14,   -18,   -34,   -22,     7,   -16,    -6,     9,     6,    11,    -9,   -15,     5,   -20,   -25,   -28,   -25,    -9,   -19,   -13,   -25,    -9,   -30,   -12,    -6,    -2,    -8,     8,    -1,    -2,   -26,   -23,   -20,   -16,   -30,    -5,    -8,    15,    12,    13,     9,     0,   -27,   -31,   -24,    -5,   -16,   -11,    -9,    -5,   -22,   -20,    -5,    -6,    -9,    12,    -2,   -11,   -16,   -21,    -4,   -18,   -13,    -5,   -12,     9,   -16,    -6,    -6,    -1,   -24,   -11,   -18,     8,   -18,   -15,   -11,   -12,   -26,   -21,    -3,    -7,   -15,    13,    -3,   -15,   -23,   -21,   -40,   -41,    -7,     1,    11,    15,   -18,   -12,   -24,     2,     2,   -16,    10,    12,    23,    -5,   -15,    -2,    -3,   -12,    -9,    -5,    -7,    -6,    -6,   -13,   -29,   -26,   -27,   -16,    -3,     9,    26,    -9,     1,    10,   -10,    16,     5,     4,    -5,     1,    10,    -7,   -12,    -8,    -7,    -7,     2,     4,    -5,    -8,    -4,   -11,   -26,   -22,   -20,   -10,   -10,     1,    24,   -15,    -2,    12,   -21,    21,    21,     5,    -8,    -8,     3,     7,   -16,    -6,   -19,    -7,     4,     5,    -8,    -5,   -15,   -11,   -33,   -27,   -14,    -2,    14,    20,    16,   -11,   -14,     4,   -31,    24,   -13,    14,     5,    -1,    -3,     3,    -8,    -9,   -22,     0,    -9,    -2,    -5,    -4,   -15,   -18,   -37,   -33,   -18,    -8,    12,    15,     5,   -19,    -8,    -3,     1,     0,     0,    13,    -3,     5,     8,     5,   -28,    -6,   -19,     4,    -6,     1,    -9,    -4,    -7,   -18,   -47,   -37,   -34,   -26,     2,     2,    -6,     7,   -11,     4,    -9,   -24,   -10,    -2,     3,    21,     4,   -19,   -16,    -1,   -14,    -6,     3,     4,   -11,   -13,    -4,   -12,   -19,   -16,   -29,   -20,    -6,   -19,    -1,    -6,    -2,     5,    -3,     9,   -13,    -3,    22,     6,    19,    -4,     2,    -5,   -11,     1,    -1,     2,    -2,     0,    -5,   -11,   -28,   -29,   -30,   -13,    -4,   -10,   -20,   -30,   -20,   -10,    20,   -16,     5,     3,    27,    -5,   -10,    -9,   -18,    -8,    -3,    -3,    -4,     0,   -13,    -3,   -12,   -14,   -11,   -28,   -26,   -24,   -17,   -21,   -16,   -18,    -4,    23,    28,    15,    17,     8,     8,   -10,    -4,    -4,    -4,    -2,    -1,     3,     0,    -4,     2,   -18,    -1,   -10,   -16,    -7,    -4,   -15,   -30,   -17,   -15,   -21,   -34,   -27,   -18,    -9,    -5,   -31,   -35,   -12,   -16,    -5,    -4,    -2,     3,    -5,    -3,    -3,     2,     1,    -4,    -2,    -4,    -4,    -6,    -7,    -6,    -9,     3,     1,   -11,    -7,   -14,   -15,     0,     1,    -2,    -5,    -1,    -4,     4,     3,     5,    -2),
		    49 => (   -3,    -3,     1,     1,     2,     1,     3,    -4,    -2,     2,     0,     3,     1,    -1,    -1,    -2,     1,     3,     2,     2,     4,    -5,    -1,     3,    -4,     4,    -1,     3,     3,     1,     2,     2,     0,     0,     3,    -1,    -5,    -4,    -6,   -13,   -13,   -11,    -1,   -36,   -33,   -29,   -11,    -5,     3,    -6,     0,    -5,     5,    -1,    -2,    -4,    -5,     3,    -3,    -8,    -6,     1,    -5,   -15,   -14,    -8,    -9,   -22,   -10,   -11,   -28,   -12,   -26,    -7,    -2,    -7,   -19,    -4,    -5,   -12,    -3,     4,     1,     0,    -3,     5,    -2,   -41,   -12,   -12,    -5,   -21,   -25,   -32,   -30,   -29,   -57,   -40,   -47,   -45,   -42,   -20,     6,   -22,   -23,   -17,   -10,    -4,    -8,    -8,    -4,     3,     1,     3,   -12,   -13,   -13,   -30,   -41,   -29,   -23,   -40,   -30,   -55,   -65,   -15,   -37,   -26,   -16,     4,    13,   -67,   -35,   -45,   -25,    -6,    -5,   -28,   -25,    -6,    -3,     3,    -8,   -13,    -3,   -15,   -31,   -26,   -28,   -26,   -16,     4,   -10,    14,   -16,    -6,   -24,   -22,   -21,   -19,   -11,   -13,   -42,   -36,   -23,   -21,   -19,     2,    -4,    -7,   -10,   -37,   -43,   -89,   -45,    -6,     1,    36,     8,    15,    -5,    28,    -4,     4,     6,    13,    18,     0,    12,    10,   -27,   -27,   -42,   -38,   -24,   -16,     5,   -22,   -30,   -39,   -68,   -85,    -6,   -26,   -10,     5,    14,    16,    27,     6,    -8,    21,    -3,    12,     7,     1,    -4,     1,   -14,   -38,   -39,   -32,   -25,    -9,   -37,   -27,   -24,   -23,   -42,    -1,    -4,   -26,     4,   -11,    -7,    -1,     0,   -18,    -1,   -13,    -2,    -5,    11,   -11,    -1,    14,   -15,   -16,   -24,   -37,   -34,   -16,    -7,   -14,    -3,   -13,   -40,    -3,    -5,     0,   -10,   -18,    -1,     8,    -2,    -7,   -13,    24,    -9,   -11,   -13,     5,     0,    13,     0,    -7,   -14,   -36,   -37,   -13,    -4,   -27,   -40,    -3,     9,     4,   -16,   -14,    -8,     9,    -7,     9,     8,   -14,   -19,   -19,    -8,    11,    -7,     8,    15,     5,    11,    -7,   -19,    47,   -38,   -26,     3,   -61,    19,    -7,    21,    -6,   -11,    -8,    11,    -6,    23,     4,     4,     6,   -16,    -8,     3,    25,     6,     7,    16,    17,    35,   -17,     4,    48,   -30,   -29,    -5,   -15,    10,    10,    37,     9,     5,    13,     2,    25,    -1,    12,   -26,   -31,     5,     1,     9,    25,    30,    34,    12,    22,    25,    36,   -39,   -75,   -44,    -8,     3,   -29,   -22,     4,    49,    38,    13,    29,    27,    16,    18,     2,     7,     8,    16,    12,    29,     0,    13,    20,    27,    20,    54,    11,   -64,   -40,   -28,     0,   -11,   -23,   -14,     9,    38,    31,     8,    13,    32,     9,    22,   -11,   -13,     8,    -7,     1,    20,     4,    14,    25,    -3,    11,    60,    -4,   -90,   -60,    -5,    -3,    -4,    -4,   -49,    11,    35,     3,   -16,    14,    38,    20,     2,   -22,   -17,     6,   -12,    20,    19,    32,    23,    21,   -11,   -21,    -2,   -21,   -80,   -46,    19,    -9,     4,    -4,   -44,   -27,     7,   -22,    -3,    -3,    -5,   -20,    24,   -20,   -10,   -11,   -10,    -2,    -5,     3,    -4,   -12,    -8,   -37,   -10,   -19,   -67,   -36,    -7,   -25,     3,     0,   -51,    -2,   -18,   -20,   -18,     4,    -3,   -11,   -11,   -30,    -7,   -14,   -15,     8,     4,    10,   -16,   -21,   -21,   -20,   -19,   -16,   -54,    -2,    -9,   -17,    22,    -1,   -47,     6,   -18,   -29,   -13,    -5,     3,    -5,     5,    -7,   -18,   -33,     0,    -7,    -5,    -2,     8,    -3,   -25,     5,    -3,   -42,   -92,    -9,   -24,   -15,     3,    -6,   -25,    33,   -15,   -34,   -29,   -32,   -21,   -25,   -22,   -17,   -26,   -56,   -10,    -3,   -15,   -13,    -7,    11,    -3,   -15,    16,   -22,   -42,    -4,   -20,    -7,     5,     0,   -45,    24,   -13,    27,   -16,   -67,   -51,   -31,   -38,    -7,   -32,   -35,     7,   -13,     5,     5,   -14,    10,   -28,   -19,   -10,    -7,     6,    17,   -11,    -4,    -2,     1,   -45,    30,     8,    28,   -15,   -27,   -29,   -26,   -39,   -31,   -31,    -2,   -39,   -16,     5,   -15,   -25,   -15,   -32,    -9,   -15,   -33,   -16,    13,   -78,    -3,     4,    -5,   -41,    26,   -23,   -10,     7,    20,    21,    -2,     9,   -15,    -7,     0,     2,     8,   -11,   -17,   -24,   -36,   -13,    -5,    -6,   -35,     3,   -11,   -47,   -10,     2,     2,   -33,    22,    -7,   -16,   -13,     5,    -1,   -16,     2,   -19,   -14,    -1,    -1,   -22,   -18,   -14,   -13,    -8,    -2,    15,    16,    -9,    -1,    -2,    -7,     4,     0,     3,   -32,   -33,    -5,    16,   -22,    12,    -8,    -4,     7,    18,    -8,   -14,   -31,    -4,     5,   -20,     3,     9,   -14,     3,    23,    28,    -1,   -11,   -16,    -1,    -4,     3,    23,   -22,    29,    12,   -37,   -44,   -15,    -9,   -29,   -23,     8,    -4,    30,    -1,    14,    23,    22,    15,    33,    40,     8,    -6,   -12,    -1,   -18,     5,    -1,     1,     0,    17,    21,     0,     7,     1,     7,     7,   -19,    -5,    22,     6,    31,     6,    14,    34,    44,    12,    32,    31,    18,    19,    18,     5,     5,    -3,    -4,    -1,    -2,    -1,   -23,   -28,    11,     7,    14,    10,    -5,     9,     3,   -14,    21,    17,    12,   -40,   -13,    21,     2,   -24,     8,   -23,     3,    -3,     0,     2),
		    50 => (   -1,    -3,     2,     3,     4,    -2,     0,     1,     3,     3,    -1,     3,    -3,     5,    -5,     2,     0,    -3,    -3,    -3,    -4,    -4,     5,    -5,     3,     5,     1,    -3,    -1,    -4,     4,     4,     5,     3,     2,     4,     4,    -3,    -1,     2,     3,     5,    -3,     3,    -3,    -4,     0,     3,    -3,    -4,     5,    -3,    -4,    -2,     4,     1,     1,    -2,    -1,     8,    13,    -8,    -7,    -5,   -10,   -12,   -17,   -29,   -33,   -33,   -17,   -24,   -19,   -19,    -8,     4,     4,    -1,   -21,    -5,     2,     2,    -5,     1,     4,    -5,     2,     3,    -1,     7,   -12,    -8,   -33,   -33,   -11,     1,     0,    12,    -2,   -26,   -33,   -15,    -9,    -2,    -7,    -3,    -9,    -5,    -2,    -4,    -4,     4,    -3,    -3,    -1,     4,    -9,   -28,    18,    -3,    20,    21,    11,    15,    -7,    -2,    -3,   -21,    -4,    10,    11,     2,   -23,   -33,    -8,    -2,    -5,    -2,    -9,    -1,     1,     3,     1,     9,     4,   -17,     0,    -9,   -29,    -5,     6,    14,     5,    14,     8,    -2,    12,     4,     8,    -6,    -7,    -8,    -1,    -5,   -15,   -21,   -17,   -21,     2,     2,   -14,    -7,    10,    -8,     0,   -12,   -13,    -5,     6,     7,     1,    -1,     3,     6,    20,     9,    11,    -7,    -5,   -22,    -9,    32,    20,   -25,   -26,    -6,     3,    -7,   -13,    -7,   -11,    14,    11,     7,    -5,    10,    21,     5,     5,     0,    10,     2,     1,    14,    -2,    -8,   -23,   -19,   -12,    12,    15,   -18,   -20,     9,     6,     0,     4,   -13,   -12,    -1,    -3,     2,    18,    20,    -5,    -3,    27,    14,    17,   -10,     3,   -14,    -2,   -13,    -3,   -10,     7,     2,     5,   -20,   -28,   -12,    -3,     0,     0,    -8,   -22,    20,   -19,    -1,    -3,     8,    -2,    -1,    -8,    -2,     3,     3,   -15,   -22,    23,    22,    24,    10,    17,    -1,    27,   -31,   -26,    -4,     4,    -3,     1,    -9,   -32,     4,     0,    -3,    10,     5,    15,    -3,   -29,   -12,    -4,    -5,   -17,    10,    15,    -7,   -19,   -10,    28,     6,    25,   -20,   -18,    -4,     0,    11,   -15,   -18,   -25,    -2,     4,    -3,     2,     4,    13,   -27,   -29,   -29,   -24,   -29,    -9,    -3,     0,   -22,   -15,   -21,   -13,     4,    17,   -11,    -3,    -5,     5,     2,     2,   -12,    -1,   -19,     6,    -8,     1,    -6,   -19,    -7,   -21,   -19,   -19,   -25,   -17,   -10,   -20,     4,    -5,   -10,    -4,   -29,     3,    -9,   -20,    -9,     0,    10,     3,     5,    23,    -2,     1,    -1,    24,     6,   -17,   -43,   -41,   -59,   -48,   -32,   -24,   -22,    -4,   -17,     1,    -3,     4,   -19,    -2,    -5,   -10,    -9,    -3,     1,    -3,   -13,   -12,    27,    13,    22,     9,     7,   -16,   -58,   -41,   -49,   -19,   -29,   -41,   -32,    -9,     3,   -13,     3,   -10,    13,    25,    -2,   -20,     1,     5,     3,    -1,   -32,     8,    24,    26,    -8,     4,    14,    13,   -35,   -65,   -38,   -12,   -18,   -26,   -25,   -17,    -2,    -6,     8,     3,    -8,     7,     0,    -2,   -16,     5,     0,    -4,   -38,    20,    23,     3,    32,   -15,    -6,     5,   -18,   -15,   -33,    -2,   -20,   -47,   -39,   -33,   -27,     9,    25,     4,    -1,    -4,   -11,   -14,    -3,    -3,     2,   -10,    -7,    13,    19,    11,     3,    -8,   -12,    13,    25,    12,     9,   -12,   -52,   -65,   -36,   -46,   -22,    -8,    -5,    -7,     4,   -15,   -16,   -26,     3,     0,     1,    -5,    12,   -17,    18,    30,    19,     6,     6,    -9,    -7,     2,   -19,   -29,   -42,   -51,   -22,   -10,    -4,    24,    13,    11,     6,     6,   -13,   -18,    -8,     0,     0,     3,     5,     2,    16,    -4,     5,     5,    -9,    -7,    -5,    11,    -8,    -8,   -20,    -1,    16,   -21,     1,    12,    18,    20,     1,     2,   -14,    -2,    -6,    -1,     3,    -3,     6,    27,    33,   -13,    -2,   -12,   -24,   -19,     5,    10,    -5,    -2,     0,     7,    10,     4,    -3,     9,    13,   -11,    -4,     5,   -17,    -5,    -4,     3,    -8,     0,    24,    36,     7,    21,     6,   -21,    -7,   -15,    -3,   -15,    -7,    17,    16,   -12,    -2,    -1,    -2,    -1,    15,    21,    -6,    -7,    -5,     0,    11,     0,    -1,    -4,    -6,     6,    17,    18,    26,    19,    -5,     5,    -8,    -2,     0,     7,     6,     7,     8,    -1,    -9,     3,    -5,     9,     6,   -16,     1,    -1,     7,     0,    -5,    -4,   -24,   -24,     5,   -10,   -17,     1,    -1,     7,     2,    17,     1,    -6,    13,     0,    18,     3,     0,   -22,   -21,    -9,    -9,   -37,     1,    -8,     1,     3,    -5,    -2,    -7,   -13,     1,    10,     9,    -4,    19,    24,     5,     9,    17,   -14,     9,    -5,    19,    12,    19,   -21,   -24,   -24,   -11,     9,     9,     1,    -4,    -4,    -3,     2,    -2,    -2,    -8,    -6,    -6,    -9,    -1,    -6,   -24,   -18,   -17,   -25,   -39,   -44,   -45,   -57,   -37,   -29,   -35,   -19,    -2,   -10,    -4,     4,     3,     4,    -5,    -4,    -3,    -5,   -10,   -12,    -9,     3,   -13,   -10,   -13,    -6,   -26,   -22,   -40,   -28,   -23,   -33,   -34,   -26,   -31,   -18,   -21,     4,    -5,    -3,    -4,     2,     0,     3,    -3,    -5,    -4,    -3,     3,    -4,    -2,    -2,    -1,    -6,     3,    -2,    -2,     0,    -6,    -5,    -5,    -5,   -20,   -17,   -22,    -4,     5,     4,    -5),
		    51 => (   -5,    -5,    -2,    -3,    -2,     5,     2,    -1,     2,     3,     2,     1,     2,    -4,     0,     0,     0,    -2,     0,     1,     4,     1,     3,    -2,     4,    -3,    -5,    -1,    -4,     0,     4,    -3,    -3,     1,     4,    -5,    -5,    -5,    -4,    -2,     1,    -4,     7,     4,    -4,    -3,    -7,     3,     0,    -2,     3,     1,     3,    -1,    -3,    -2,     1,    -2,    -1,     1,     1,    -3,    -4,    -3,    -8,   -15,   -30,   -27,   -19,     6,   -21,    -7,    28,     7,   -28,   -28,    -8,   -17,   -15,    -9,    -4,     4,     0,    -4,    -1,    -2,    45,    26,     1,   -20,   -12,    -4,   -12,   -15,   -26,   -39,   -22,    -4,   -17,   -24,    -9,   -13,    -6,    36,    30,   -27,    -5,   -15,    -6,    -4,     5,    -4,     1,     2,    40,    42,    -3,   -22,   -13,   -10,   -11,   -28,   -35,   -13,    -4,    22,    20,     0,   -23,   -36,    19,     8,    11,   -11,    -5,    -9,     0,    -6,   -17,   -16,    -3,     0,    39,    21,     7,    -3,    -2,   -17,   -44,   -50,   -11,     3,   -13,    10,     3,     3,    13,   -28,   -14,    -8,   -23,   -15,   -10,    -3,    -5,    -4,   -15,   -16,     0,    -2,   -15,     4,     2,    -8,   -17,    -3,   -42,   -54,   -27,     0,     7,    26,     9,   -16,     4,   -33,   -10,   -31,   -29,    -8,    -4,     3,     0,     1,   -12,   -13,     2,    -5,   -18,     4,    -3,   -22,   -26,    -9,   -59,   -36,     1,     9,    18,    27,     7,    -8,   -19,   -25,   -11,   -56,   -24,   -14,     1,    -4,    -2,    -8,   -32,   -15,     2,    -6,   -16,     7,    -9,   -15,   -24,   -21,   -57,   -27,     2,     0,     5,    19,    31,    19,   -24,   -21,   -14,   -55,   -16,   -13,    12,     0,    -5,    -3,   -20,    -7,     3,    -7,   -19,    -8,    -7,     2,   -13,   -11,   -29,    -1,    10,    -6,   -26,     0,    34,    27,   -21,   -39,     1,     4,   -22,    -2,     9,    -3,   -17,   -10,   -17,   -27,     0,    -7,    -8,    -7,   -15,    -5,   -28,   -13,   -11,   -27,    24,    -2,   -10,    13,    18,    -3,   -11,   -30,   -23,    -1,    -8,   -39,     4,    15,   -22,   -11,     5,    23,     1,     4,    -3,    -7,    -7,   -15,   -35,   -19,   -32,   -22,    -6,    13,   -11,     3,    27,    -7,     0,   -19,   -30,   -11,    15,    -4,    12,    15,   -20,   -13,   -10,    40,     5,     0,   -37,    15,     1,    -2,   -12,   -12,   -10,    23,     7,    -4,     6,     3,    16,   -12,    -4,   -33,   -37,   -19,    31,     3,     5,    19,   -22,     3,     3,    30,     2,    -3,   -36,     2,     2,    -5,    -4,     8,    25,    15,   -38,     7,     8,   -17,   -10,   -13,    -6,   -20,   -24,     9,    35,   -13,   -16,   -30,   -24,    21,    16,    -5,    -1,     0,    -3,     4,    -4,   -19,     1,    12,    -9,   -13,   -34,   -22,     8,    -2,    -5,   -16,     4,     2,     0,     3,     9,   -14,   -27,    -4,    -3,    -7,    25,     5,    -4,     0,     4,    13,    -1,   -23,   -19,    -1,    -8,   -14,   -13,    30,    18,    24,     9,   -25,     1,    -3,    18,    -8,    22,   -10,   -24,    -7,   -24,   -14,     2,   -13,     1,    -3,     4,   -15,    -2,   -13,    -8,     1,    -8,   -19,   -11,    15,     8,    -1,     7,   -19,   -18,    -4,     7,   -19,     3,   -11,   -17,   -18,     0,   -21,     0,    -7,    -2,     5,     1,    -7,    -6,   -23,   -17,   -24,    -8,   -14,   -15,   -10,     5,     4,     4,   -10,   -14,   -20,     5,   -21,   -26,   -16,    10,    11,   -13,   -21,    -6,     5,    -3,     1,    -5,    -4,   -13,    -1,   -17,    -9,   -24,   -15,   -50,   -10,   -17,    29,    14,    -2,     4,    -6,    14,   -33,     9,    -5,   -27,   -25,   -24,     2,    -1,    21,    -4,    -3,     4,    -4,    -5,    -2,    -6,   -15,     9,   -26,   -26,   -10,    -5,    13,    25,    13,    -1,   -18,   -11,   -42,   -13,   -14,   -36,   -22,   -10,    12,    16,    23,     5,     4,     0,   -13,   -13,    -7,   -15,   -31,    -8,   -10,    -8,    -6,    22,     8,    11,     8,     3,    -7,   -11,   -18,     1,   -30,   -46,   -17,    -1,    -4,    22,    -3,     8,     7,     3,   -12,   -13,    -5,   -21,   -46,    -3,    -1,   -13,     0,     2,     4,    -5,     2,    -8,   -29,    21,    -7,     9,   -10,   -34,   -31,   -14,     8,    -9,    -2,    11,     5,     4,     4,    -9,    -6,    -8,   -37,     3,    -2,    -6,   -17,   -12,    -3,     3,    -7,    -8,   -11,    11,     5,    18,    -3,   -29,   -12,   -24,    20,    16,    -1,     3,     0,    -6,   -13,    -4,     4,    19,   -13,     5,    29,     2,    16,    -5,     1,    -1,     2,     6,    28,    24,     7,    16,   -11,    -5,   -16,   -18,    -5,    37,     4,    -4,    -3,    -4,    -6,    -5,    -5,    24,     4,    -4,     4,    21,    29,    -4,   -25,   -24,   -34,   -43,   -17,   -32,   -21,   -19,   -11,   -30,    -3,   -18,    25,    21,     4,     3,    -1,    -4,     0,    -3,    -3,    -1,    -4,    -7,   -14,   -64,   -52,   -36,   -31,    -8,   -40,   -38,   -42,   -35,   -37,   -60,   -23,   -18,   -17,    -1,    -2,    -4,     2,     4,    -4,    -2,    -2,   -14,   -30,   -22,   -19,   -19,   -16,   -13,   -18,   -30,   -32,   -33,   -32,   -24,   -24,    -6,   -13,    -2,   -15,    -1,    -2,    -3,     2,    -1,     1,    -4,    -1,     4,     0,    -4,     3,     0,     1,    -4,     5,    -3,    -3,    -1,    -4,    -7,    -5,    -1,     1,     3,    -3,     0,     2,     1,     1,    -3,    -5,    -3,    -5),
		    52 => (    1,     3,    -3,    -4,     2,     1,    -5,     4,    -2,     0,     3,     5,    -7,    -6,     4,     9,     2,     4,     4,    -2,     1,    -4,     3,    -4,     1,     5,     2,    -1,     2,    -2,     4,    -5,     5,     5,    -5,    -3,    -2,     3,     4,    -3,     3,     4,    -9,    -7,     5,     7,    -3,   -21,   -10,    -1,     1,     3,     3,     3,     2,     5,    -2,    -1,    -7,    -8,    -7,     5,    -6,    -9,    20,    30,    36,    18,    15,   -10,     0,   -14,   -36,   -27,    -1,    10,     1,    10,   -10,     8,    15,     9,    -4,     1,    -4,    -3,    -8,   -30,   -24,   -27,    -8,   -15,    10,    10,    -4,    -5,   -11,     7,    14,    -6,    -2,    -4,    -6,    24,    -7,    -6,    -8,   -36,   -19,     9,    -9,     0,     0,    -3,    -5,    -8,    22,    -6,    -4,     4,     1,     5,    -9,     1,    14,     6,    -2,    10,   -16,     8,   -18,    -6,    12,   -19,   -10,   -33,   -36,    15,   -26,   -12,    -3,    -4,     0,   -12,     4,   -29,   -32,   -43,   -20,    -3,    21,     3,   -15,    12,     7,     6,   -13,     6,    -4,    -1,    -1,     7,    -2,    17,   -29,    29,   -21,    -3,    -3,     1,     1,    30,    24,   -25,   -20,   -11,     9,    20,    20,     2,     3,    23,     5,     0,    -9,     5,     2,    -4,    -8,   -21,    -8,    -5,     2,   -23,   -23,    -3,     1,     0,    -8,    38,    29,    20,    -7,     5,    -6,     1,    -5,     9,     6,    12,     3,    15,    18,    17,     6,    14,    -8,   -15,    25,     3,   -20,   -23,   -19,   -16,   -14,    28,    -5,    28,    18,    15,   -20,    -8,    -9,    15,     1,    -4,    -8,   -15,    -6,     4,    14,    21,    -4,    24,   -17,     0,    23,    21,   -55,   -34,   -24,   -17,     5,    -9,     8,     6,    -8,     6,   -13,   -15,    -7,    19,   -20,     2,    11,   -27,    -8,     4,    12,     6,    -5,    23,     1,   -14,   -14,    21,   -45,   -29,   -14,    -7,     1,    -1,     3,    16,   -31,    34,    17,    -2,    -7,     1,   -18,   -23,    -1,    13,    -8,    -8,    -7,   -11,    -3,     6,    12,    -3,   -10,    21,    -9,   -10,     4,    -6,     1,   -14,    -4,    21,     4,     7,    16,     1,    -8,   -20,   -43,    -1,   -14,   -25,   -30,   -25,     1,    -9,   -23,    -5,   -12,    -2,   -11,    10,    -4,     1,   -22,    -4,    -3,     0,   -28,    -2,     6,   -31,   -12,   -23,   -28,   -21,   -25,   -23,    -9,   -38,   -47,   -12,     0,    -5,   -26,    -5,   -17,    -8,    -5,   -14,    -7,    12,    -2,   -12,    -1,     3,     2,    -3,    -5,   -12,   -43,   -38,   -64,   -38,   -29,   -37,   -48,   -27,   -22,   -11,    -9,   -21,   -18,   -22,   -19,   -21,     8,   -17,    -4,    12,    21,   -11,     4,   -15,   -19,    -7,   -25,   -45,   -50,   -51,   -79,   -50,   -26,   -27,    -8,   -15,     0,   -11,   -28,   -10,   -10,    -9,   -22,   -35,    -4,   -39,    -4,     2,    26,    14,     4,   -13,    -3,   -11,   -48,   -26,   -23,   -34,     6,    -3,   -12,    13,    -1,    16,     5,   -24,     4,    -4,   -29,   -34,   -34,   -20,   -37,   -19,     9,   -11,    30,    42,     0,    -1,   -19,   -31,   -54,   -19,   -22,   -16,    -8,     9,    10,    10,   -18,     7,     9,   -10,   -15,    -6,   -14,   -31,   -21,    -8,    14,   -12,    12,    29,    38,    26,    -4,    -3,     2,   -22,   -19,   -24,    -2,    -7,    -1,     2,    12,     5,   -17,    28,    18,     1,    -4,    -7,    -4,   -27,   -16,    -9,    -8,   -10,   -21,    49,    29,    24,    -3,    -4,    -7,   -42,   -15,   -11,    13,    19,    -8,   -13,     4,    -2,     9,    -3,    -4,    -6,    -4,    13,   -15,   -20,   -25,    16,    19,    19,    36,    60,    -4,    31,    -3,    -9,     9,   -21,   -25,    -9,    19,    12,   -13,   -19,     9,     6,     2,    38,    33,    10,    16,    -3,    -7,   -16,     3,    20,     9,    18,    -5,    17,    16,    32,     2,    -4,    19,    -2,    -2,   -13,    45,    15,    11,    14,    32,    27,    19,    51,    18,    14,    29,    -3,    -5,    -5,    31,    29,    11,     8,     6,    24,    11,     1,     4,    10,    10,    24,     8,     6,    23,    15,    -6,    13,    10,    12,     2,    38,    30,    24,    15,    20,     9,    15,    17,    14,    23,    50,    24,    24,    23,    -7,     2,    -2,    -1,     0,    -3,    25,    35,    19,     4,    20,     5,     8,     5,     3,    13,    10,   -10,   -22,    -1,   -21,     8,    22,    37,    44,    35,    -3,   -33,   -11,    -4,    -4,     4,   -23,   -12,     7,    26,    14,    10,    23,    10,    33,    25,    18,     6,    -7,   -21,   -14,   -15,    -1,    18,    26,    47,    33,    26,     4,   -17,     1,     2,     0,   -25,   -17,    -6,   -14,     1,    14,    35,   -10,     3,     2,    23,   -11,    14,     7,   -25,    -8,    -1,     1,   -28,   -15,    -2,    26,    53,    29,    17,     1,     4,    -1,   -16,    -2,   -21,   -51,    23,    -8,   -26,   -51,   -67,   -20,   -10,    -4,    22,    17,   -17,     6,   -34,   -44,    -4,     7,   -37,   -16,     9,    27,    19,    -2,     3,    -4,    -3,    -1,   -17,   -31,   -35,   -23,   -22,   -33,   -57,   -46,   -27,   -29,   -30,   -18,   -45,   -41,   -33,    -3,   -14,   -19,   -12,     1,    -5,     0,    -5,     3,    -5,     4,    -4,     3,    -3,     0,    -6,     1,     4,    -1,   -15,   -25,    -2,   -11,    -2,    -1,     1,    -5,    -3,     2,    -9,   -17,    -9,    -2,    -2,     1,     0,     0),
		    53 => (   -1,    -2,     1,    -3,    -1,    -3,     5,    -5,     3,     1,     1,    -4,    -5,    -4,    -2,    -1,    -3,    -2,    -2,    -2,     5,    -4,    -4,    -2,     3,    -2,     0,     0,    -3,    -1,     3,     1,    -3,    -1,     3,    -2,     5,    -5,     1,    -1,    -4,    -4,    -9,    -3,   -11,    -5,     0,    -3,     0,     1,     4,     2,     4,     5,     1,    -5,     3,     5,     2,    -4,     1,     3,     3,     0,   -20,   -24,    17,    20,    14,    -9,   -19,   -20,   -29,   -30,   -21,   -10,    -4,   -14,   -16,   -22,    -7,    -5,    -1,     0,    -3,     1,    -1,   -12,    -5,    -1,    -7,     9,     4,    -6,    15,    17,    11,    13,     3,   -12,     7,    16,    19,    -8,    -8,   -11,    -5,   -37,   -17,    -4,    -1,     1,    -4,     9,     2,     0,    -6,     4,     5,    13,     6,    -5,    -9,   -16,   -22,   -25,     0,   -10,   -12,   -30,   -14,     1,   -19,   -16,    20,   -40,   -34,   -18,    -5,    -1,     0,     2,     4,    -8,    -4,    14,    20,    33,     3,   -23,   -33,   -15,   -11,   -14,     0,    -6,    -4,    -4,    -6,     5,    -5,   -14,   -19,   -15,   -15,    -4,   -14,    -5,     0,     7,    -1,     9,     3,     0,     4,    -4,   -26,   -19,    15,    -4,     2,    -9,   -14,    -9,    -4,     0,     1,   -20,   -16,    -7,    -7,    -5,    -6,   -31,   -18,    -7,     4,     9,    14,   -20,   -45,   -19,     1,   -14,   -23,    -9,    -9,     4,    -8,    -1,     3,     3,    -5,    11,    -2,   -21,     5,   -13,    -3,   -17,   -11,   -25,   -18,    -8,     0,    -5,    12,   -28,   -37,     0,   -13,   -20,   -12,     7,     7,    -5,     1,   -15,     4,   -12,     3,     2,    17,     4,     9,    26,    16,   -35,   -59,   -19,   -26,     1,    -3,   -23,   -19,   -22,     4,     2,    13,    -3,    -7,    -8,    12,    19,    28,    14,    13,    -9,   -14,   -10,   -15,   -10,    17,    11,    11,   -28,   -70,   -28,   -29,    -5,     0,   -24,   -11,    16,     7,     6,    30,     3,    41,    19,    22,    18,    -1,    -1,    -4,   -13,   -35,    -2,    15,    16,    11,    -5,    13,    -8,   -65,    -6,   -21,     2,    -2,   -25,   -11,    37,    34,    32,     7,    20,    12,    27,    10,   -19,   -41,   -40,   -34,    11,     8,    11,    17,    21,    33,     6,     8,    -2,   -39,   -36,    -8,    -5,    -2,   -25,   -22,    38,    21,    15,     0,     9,   -24,   -23,   -32,   -71,   -52,   -12,    18,    31,    11,     4,    15,    -2,    -7,   -17,   -11,   -24,     0,     3,     1,     3,     2,   -17,   -47,    16,   -24,   -16,   -12,   -15,   -33,   -66,   -68,   -43,    -9,    11,    23,     5,     6,    -3,   -14,   -18,   -12,    -7,   -36,   -27,    22,   -13,   -11,    -4,    -8,     7,    -7,   -12,   -32,   -38,   -55,   -51,   -50,   -26,   -11,   -20,    11,    18,    10,     7,    -6,     5,   -26,   -16,   -21,   -15,   -38,    -7,    32,    -8,   -18,   -12,    -2,    16,     7,     4,   -11,   -20,   -42,   -56,   -41,    -2,    10,    -9,    13,    27,    44,     0,    14,    -5,    -6,    -2,    -9,     2,   -18,   -10,    25,   -10,    22,     4,     0,     4,    12,    24,     5,   -15,   -23,   -15,   -33,   -22,   -24,   -45,    -5,     4,    -9,   -22,    14,    10,   -14,     3,     3,    28,    -6,   -21,    14,   -26,     9,     1,    -1,     2,     6,     6,     2,    -2,    -9,   -21,   -43,   -55,   -69,   -76,   -92,   -75,   -48,   -29,    18,    -5,   -23,    17,    14,    28,     9,   -19,    -8,   -34,    -4,    -2,    -9,     4,    28,     7,    35,     3,   -16,     0,    -7,   -36,   -33,   -50,   -72,   -55,   -34,   -32,    -2,    22,    17,    18,     6,    -4,    12,    -8,   -44,   -13,     2,   -11,    -1,   -15,   -18,   -15,     9,    15,    -1,     1,   -12,    10,    -5,   -16,   -12,     0,     1,   -10,    -9,     1,   -11,     0,     4,     1,    21,     0,   -14,     8,    -6,   -11,     3,    -3,   -18,    -3,     9,    17,    19,    13,     4,    23,    20,    28,    12,     0,    -9,   -27,   -10,   -19,   -15,     4,    19,    -4,     7,   -16,   -21,   -15,    -4,    -5,    -3,    11,    -8,     1,    -8,    10,     5,    20,    22,     7,     1,     0,     4,    -9,     1,   -19,   -18,   -27,    -7,     9,    13,     0,   -10,   -15,   -23,   -10,    -9,     0,    -5,     3,   -13,     3,     3,    -6,   -12,   -16,    -2,    -4,     5,     3,     6,     6,     9,    -5,    -3,     2,    -3,    17,    -2,     4,   -27,   -25,   -22,   -11,    -7,     4,     1,     2,    14,    20,    23,    15,    -6,    -9,    -6,    -5,   -25,   -10,   -18,    -7,    -8,    14,     3,    13,    14,     0,     6,    11,   -28,   -22,    19,    12,     1,     1,    -2,    -2,    -1,    16,    20,     0,   -18,    -9,     3,    13,     1,     4,    11,     3,     2,    -9,    18,    17,   -10,   -28,    -7,    -9,   -20,   -32,   -21,   -12,    -6,     0,    -1,     4,     1,   -21,   -17,     7,    12,     7,   -12,   -10,   -36,   -31,   -24,   -45,   -30,    -2,    -1,   -24,   -24,   -24,   -14,   -16,   -15,   -28,    -1,     0,     3,     1,    -3,     0,     1,   -16,   -38,   -35,   -25,   -29,   -38,   -34,   -48,   -41,   -35,   -18,   -13,   -14,   -20,   -50,   -45,   -39,    -2,   -16,    -4,    -1,     3,     2,     0,     2,    -2,    -3,    -3,    -5,    -3,    -7,    -7,    -9,    -8,   -24,   -18,   -22,     0,   -17,   -16,   -21,   -16,   -16,   -16,   -23,   -10,    -5,    -3,    -1,    -3,    -2,     5,     2),
		    54 => (   -2,    -2,    -3,     3,     1,    -3,     3,    -1,    -2,    -5,     2,     0,    -6,    -6,    -6,    -5,     4,    -5,    -5,    -1,    -5,    -5,     2,    -4,    -5,    -3,     2,     4,    -1,     5,     3,     4,     4,    -2,   -21,   -17,    -5,     1,   -10,    -1,    -8,     6,    19,    -4,    -5,    -3,    -5,    -3,   -10,    -7,    -7,    -4,    -5,     5,     0,     0,    -4,    -1,    -2,    -8,   -29,    -2,   -13,   -21,   -31,   -10,    -7,    -5,    -9,   -20,   -16,   -28,   -37,   -15,    -9,    -4,   -24,   -20,    -2,    -6,    -4,   -15,    -1,     1,     0,     0,    -9,   -14,   -23,    -8,   -17,   -22,   -10,    -4,   -11,    -6,     3,   -11,   -19,    -3,     3,    14,   -18,   -13,   -18,    -7,   -11,     0,    -3,   -10,     2,     1,     3,     1,    -8,    -5,    -9,   -14,   -24,    13,    30,    16,   -12,   -37,   -47,   -29,   -25,   -23,   -40,   -49,   -51,   -33,   -15,   -11,     4,    42,    31,    19,   -37,    -7,    -4,    -4,   -11,     4,   -13,    -1,   -13,    10,    43,    12,   -27,   -47,   -32,   -18,    47,    27,    20,    -9,   -48,   -59,   -21,   -19,    -4,    13,     8,   -13,    -6,    -5,     1,     2,    -4,   -18,    18,    24,    -9,    18,    19,   -19,   -54,   -63,   -11,     7,     8,    22,    20,     6,   -46,   -87,   -79,    -9,    27,    28,    17,   -40,    10,   -28,    -1,   -16,     1,   -18,    12,    19,    10,    14,    -4,   -10,   -30,   -20,   -29,    -2,    22,    22,    15,    13,   -66,   -92,   -42,    12,    38,    42,     4,   -49,     3,   -35,   -11,   -16,    -2,   -22,    -2,    22,    14,    17,    -6,    -7,   -22,   -30,   -38,     3,    16,    35,   -12,   -45,   -81,   -42,    -7,    21,    12,    -6,    -3,   -18,    10,   -25,    -3,    -6,    -8,   -24,     7,     1,    14,    33,     0,   -15,   -20,   -38,   -14,    -1,    28,    15,    -7,   -43,   -40,   -17,    14,    16,    -6,     7,    -6,   -12,    11,   -22,     2,    -9,   -23,   -26,    -9,     1,     6,     4,   -25,     8,    -8,   -31,    12,    -2,    24,     7,    -7,   -26,   -26,    -1,    10,    -2,     3,   -16,     4,    12,    -4,   -19,    -4,     2,   -22,   -13,   -19,     9,    -6,    -8,     4,    14,    -2,     7,     8,   -24,     2,     2,   -14,   -26,   -19,    -6,     0,     3,     7,    -1,   -18,    -2,   -15,   -35,     1,    -1,   -15,   -53,   -16,    12,    -9,     2,     6,     5,    14,   -20,     7,     6,    -3,   -14,   -16,   -14,   -25,     4,    10,     5,     4,   -22,    -4,   -15,   -39,   -29,    -2,     5,   -17,   -36,   -24,    -4,     0,    10,    -1,    11,    31,     1,   -23,    14,   -22,   -16,    10,     0,    -6,    12,     2,     3,     1,    -6,   -24,   -32,   -37,    -2,     3,    -2,   -15,   -33,   -10,     0,    18,     1,     1,    11,    16,     3,     1,    17,     9,   -10,    -1,    16,    -8,     1,     5,    12,    13,   -13,    -1,   -22,   -10,     2,    -4,    -2,     0,   -31,    -3,     5,    10,    26,    20,    16,    14,    10,    12,    -1,     8,    -4,   -16,     4,     3,     4,   -10,   -12,     4,     0,   -13,   -15,    -6,     7,     4,    -2,    -4,   -25,   -14,     8,    23,    28,    14,     0,   -13,    -6,    -2,    -4,     2,    20,    10,     3,    -5,     1,    10,    -9,   -21,   -19,    -6,   -12,   -28,    -9,    -2,     2,    -8,   -14,    -8,     2,     8,     2,    15,   -11,    -1,   -11,     1,    -3,    19,     7,     5,    -7,   -11,   -13,   -12,    -7,    -3,   -13,   -27,   -25,   -15,   -12,   -14,    -3,    -1,    21,    18,    -7,   -16,   -19,   -13,     6,   -33,   -31,   -17,     3,    17,    -4,   -10,   -12,    -9,   -21,   -35,   -15,   -18,   -21,   -11,   -18,    -7,   -12,    -5,   -11,   -13,    31,     9,   -45,   -31,   -16,    -8,    -5,   -44,   -26,   -16,   -24,     1,    -5,   -11,    -8,    10,   -15,   -27,   -30,   -26,   -27,    -2,   -15,    -9,    -9,     0,     0,     0,   -13,    -1,   -14,   -14,   -17,   -27,     6,   -21,    -3,     1,   -23,    21,     2,   -13,    -1,    19,   -19,   -44,     2,   -11,    -8,    14,   -21,    -5,     4,     1,    -1,   -10,   -40,   -22,     2,   -22,   -29,     6,     9,    -2,     5,    -7,   -38,    -1,   -12,    -4,   -11,     5,    -6,   -32,    -4,   -11,     5,     3,   -26,   -13,     1,     1,    -2,     3,   -23,   -23,     4,    -5,     9,    17,   -16,    -6,    -2,   -11,   -21,    -8,   -13,     4,   -14,     4,    21,    -6,     2,    12,    -5,    15,     3,     3,     4,    -5,     0,     0,   -13,   -17,   -34,   -10,     7,     8,     1,    28,    13,     7,   -22,   -16,   -24,   -23,   -17,     2,     8,    15,    -3,   -12,     1,     9,    14,     0,     2,    -1,    -4,     2,     0,   -29,   -26,    11,     8,     7,     4,     3,    25,    18,   -16,    -5,    -4,   -37,     1,     8,     9,    20,     3,    19,    10,    -2,    26,     2,    -2,     3,    -1,    -5,    -4,   -19,   -42,     8,     0,    -2,    -2,    14,    15,   -37,   -54,   -17,     2,   -32,     7,   -19,   -32,     1,     2,    16,     2,    -4,    -9,    -1,     3,     3,    -2,     4,   -22,    -7,   -23,   -27,   -11,   -17,   -20,   -30,   -22,   -26,   -34,    -8,     2,    -7,     7,   -26,   -33,   -35,   -39,   -29,    -2,    -4,     2,     1,     5,    -2,     1,     2,     2,    -2,    -4,   -10,   -13,   -14,    -9,   -24,   -19,   -15,   -18,   -32,    -4,   -15,   -26,   -22,   -19,   -26,   -17,   -20,    -4,     0,    -1,     1,     1),
		    55 => (   -4,     0,     3,    -2,    -1,     4,     1,     4,    -3,    -4,     3,    -2,     1,    -7,     3,     3,     4,    -4,     1,     0,     5,     2,     5,    -1,     0,    -3,     1,     2,    -2,    -1,    -4,     0,    -1,     0,    -1,    -6,     1,     0,    -3,   -16,    -9,    -6,   -20,   -25,   -22,   -26,   -18,   -21,   -29,   -28,   -10,    -2,    -1,     3,    -2,     0,    -3,    -3,   -16,   -16,    -7,    -8,   -15,   -14,   -25,   -39,   -36,   -41,   -50,   -64,   -32,    10,    13,    19,    10,    -8,    -2,   -22,   -23,    -5,   -21,   -15,     4,    -2,     3,     3,    -8,     0,    -7,   -24,   -46,   -29,   -60,    13,    23,    -3,     7,     0,   -16,   -28,   -24,    -1,    14,    29,    -4,    24,     1,   -21,   -11,    13,    39,     0,    -3,   -11,   -20,     0,   -26,    -4,    -2,     5,     1,    -5,     9,    -2,     9,   -13,    -6,   -16,   -26,   -16,    17,   -23,   -21,    -4,   -13,   -11,    39,    26,     6,   -13,    -2,     3,   -20,     0,   -20,    -7,   -16,     3,   -15,     1,     0,    34,    27,    -9,    11,    22,    -3,   -19,   -45,    -9,    -3,     0,     4,    19,    -1,    24,     9,    -3,     5,     0,    -2,   -28,   -29,   -14,     1,    13,    12,    -3,     0,    24,    34,     4,     4,   -12,   -18,   -22,   -23,    -4,    -9,    -8,     8,    32,    31,    39,    -4,     5,     3,   -16,     4,   -47,   -43,   -19,    14,    31,    28,    23,    25,    10,    -4,     4,    14,    -1,    18,     6,   -26,    -7,     7,     0,     3,    -1,     8,     9,   -10,    17,    -5,   -13,   -37,   -61,   -31,    20,    -1,   -22,    -5,     8,     9,    -2,    -2,     3,    18,    19,    -3,    13,   -21,   -41,   -11,   -11,     4,    -1,    44,    17,   -32,     9,     0,    -4,   -28,   -44,   -17,    18,    10,   -26,     6,   -13,     3,    33,    20,    30,    43,    26,     3,   -12,   -43,   -47,   -47,   -24,     8,    -1,    24,    27,   -17,   -12,    -1,    -2,   -35,   -74,    27,    29,    18,     9,   -13,   -10,    15,    27,    48,    34,    32,    36,     1,   -45,   -23,   -32,   -31,   -19,   -62,   -52,    20,    28,    26,   -16,     3,    -7,    -3,   -16,     7,    16,    12,    -5,    -8,   -11,    -1,    11,    22,    23,     9,    26,    12,    -4,   -15,   -39,   -22,   -18,   -63,   -71,    -3,    -4,    12,     5,    -3,    -4,    -6,   -11,    20,     8,    -1,     3,     0,    -2,     0,   -22,     4,     4,    -4,     5,   -14,   -17,     0,    -9,   -26,    -8,   -46,   -30,   -70,   -30,    27,   -30,     0,    -2,   -13,    -3,    -1,    16,   -12,     1,    -4,    -3,    -1,    10,     3,     4,    -5,     7,    -8,   -23,    -2,    12,     3,     4,   -10,   -37,   -57,   -43,     1,   -20,     5,    -5,    -5,     3,   -29,    -5,    -9,    -6,   -14,    -3,    -3,   -12,    -1,   -17,     4,   -13,    14,    -3,   -12,     4,    13,    -5,     0,    33,     2,   -28,   -17,   -11,     1,     2,   -15,   -10,     4,     0,    -3,    -4,   -36,   -24,     6,    -3,     3,   -12,    -3,     1,    -7,    -4,     3,   -12,   -18,   -37,    -2,    32,    14,   -28,   -27,   -30,     1,    -9,   -35,    30,     3,    11,   -41,   -61,   -29,   -32,   -15,    27,    -4,    -5,    -7,   -19,    -7,   -19,     0,    10,   -11,   -12,    -3,    14,   -10,   -61,   -36,   -34,    -2,    -7,   -53,    53,    11,     1,   -12,   -55,   -38,   -29,   -13,    -3,   -20,   -13,   -14,   -12,     7,    18,     6,    22,     0,    -1,     5,    11,   -34,   -61,   -49,   -50,    -7,     4,   -36,    52,    51,    29,    -3,   -31,   -43,   -61,    -9,   -26,   -16,   -25,    -1,    -3,    12,    15,    -4,   -12,    10,    16,    17,    28,    -3,    -9,   -54,   -17,     0,   -14,    28,     3,    41,    38,    11,   -20,    -9,   -34,   -14,   -18,    -4,    -4,     0,    14,   -11,     9,    28,    -1,    32,     2,    20,    29,    32,    18,   -33,   -36,    -5,   -14,    22,    -5,    18,    21,     4,     0,     2,    -6,   -21,     0,    -4,    15,    -5,   -10,    15,    22,     3,   -19,    15,    -5,    39,    17,    17,    30,   -29,    -1,    -3,    -5,   -26,   -48,    -3,    18,   -11,   -17,    19,    18,    -1,    -8,   -10,    -2,     9,    24,    22,    11,    22,    21,     6,    23,    -4,    26,    10,    43,    15,    -6,    -6,    -2,   -39,   -16,   -30,   -28,   -16,     3,     5,    11,    12,    -5,     0,     7,    -6,     1,     7,     0,     6,    20,   -13,     0,    -1,    44,    46,    55,    35,     1,     2,     3,     7,     9,   -14,    -9,     4,    -6,   -24,     2,    -7,    -4,   -10,     8,     9,    -4,     8,     7,    17,    18,    -7,     8,   -12,    32,    31,    38,    26,    -2,     5,    -3,   -25,    -7,   -20,   -12,   -16,    10,    13,    35,    24,    21,    -6,   -15,   -26,     6,    -7,    24,    20,    26,     9,   -14,     8,     0,    36,   -24,   -14,     1,     5,     1,     0,    19,   -38,   -47,   -16,    -7,     7,   -17,   -24,   -23,     1,   -13,   -29,     0,    27,    37,    34,    24,     5,    26,    42,    36,    36,   -13,    -5,    -3,     5,     4,    -5,   -11,   -17,   -36,   -47,   -43,   -16,    -4,    10,     8,     0,    -8,   -39,    13,    -7,    11,    10,    40,    11,    -1,   -10,   -20,   -11,     4,     4,     3,    -2,     5,     4,    -1,    -9,    -8,    -3,    -9,   -10,   -11,     5,     5,     6,     3,   -49,   -37,   -11,   -17,   -11,   -23,   -28,   -32,   -18,    -3,     3,     4,     2,     1),
		    56 => (    0,    -2,     0,    -2,     3,    -2,     4,    -1,    -3,     1,     0,    -5,     8,    11,    -3,     5,    -4,     4,     2,     1,     5,     2,     2,     1,     0,     1,     2,    -2,     4,     1,     0,    -5,    -5,    -4,    11,    12,    23,    14,    11,     8,     4,    17,    -2,    -7,    -5,    -4,     1,     5,    29,    14,     9,     2,    -1,    -2,     0,    -1,     0,    -2,    -2,    -1,    15,     0,     8,    26,    22,    20,    12,    -8,   -11,   -13,   -11,    -5,     0,    -3,    -3,    13,    16,    21,    16,    27,    10,    10,    -3,    -3,    -3,    -4,   -22,   -23,    -5,    17,    15,    12,     8,    14,    -4,   -18,   -23,   -46,   -21,   -11,    -3,   -19,     9,    28,    16,    11,     6,    26,    18,     3,    -2,     1,     5,     0,   -27,   -29,    20,    27,    17,     3,   -10,     9,     3,   -25,   -32,   -47,   -31,    -3,    -7,   -13,   -31,     2,     2,    -9,   -20,     2,    20,    17,    31,    34,    -4,     5,   -14,   -26,    41,    23,     9,     5,     7,     3,    -1,   -12,   -18,   -34,   -13,    11,    -6,     5,   -13,   -14,   -15,    -6,   -11,     6,    13,    15,    34,    23,    -2,     0,     8,    -6,    31,     9,    16,     6,    34,    14,   -15,   -32,   -34,   -37,    -8,   -10,   -28,   -12,    -1,   -27,   -16,    -2,    -5,    -1,     4,   -19,     8,    40,     1,    -1,     2,    -9,    33,    13,    -6,    18,    15,    19,   -10,   -29,   -39,   -21,     0,   -27,   -33,    -2,    -2,    -4,    -5,   -16,   -18,   -21,   -21,    -8,    14,    35,     0,     2,     2,   -11,    24,     8,    -6,    14,     3,    -2,   -22,   -39,   -43,     1,     3,   -30,    -5,    13,     7,    12,    14,     5,   -17,    -6,    -5,   -11,    15,   -21,    -3,    -3,    -5,   -21,    15,     6,    -8,    12,    -4,   -19,   -41,   -46,   -41,   -14,    -6,   -12,     9,    23,     3,    10,    17,     2,    -7,     3,    -4,   -21,    -7,    -7,    -2,    -3,    -8,   -20,    24,    16,     9,    29,     3,   -20,   -32,   -39,   -31,    -7,    -4,     4,     4,    20,   -17,    -9,   -11,     8,     1,     3,   -10,    -8,     0,    -4,     0,     2,     4,    -6,    19,    18,    13,     7,    -2,   -15,   -25,   -30,   -18,    -3,     4,    -3,    -9,   -35,   -23,    -6,   -15,     0,     9,    12,     3,     2,    -8,   -11,    -5,     1,    -5,   -10,    12,    29,    -1,     7,    -2,   -16,   -24,   -34,   -10,    35,     6,     4,     5,   -13,   -12,   -19,    -8,    10,    20,    16,    13,    -3,    -4,   -21,     4,     5,    -3,    -9,     5,     6,    -5,     1,     8,   -13,   -15,   -37,     1,    19,    -7,   -18,    -3,     2,   -14,   -13,    -8,     9,     8,    15,    13,    -1,    -3,    -5,    -3,    -1,     2,   -14,     3,     6,    -6,     7,     0,    -3,   -20,   -13,    17,    22,   -32,   -23,    -1,     3,    -5,    -5,   -18,    -6,     2,    11,     9,    -2,    -7,    -8,    -4,     0,     2,    -8,    12,     5,    -8,    -3,    -2,    -2,   -18,    -1,     0,    11,   -13,    -5,     2,    -6,    -2,   -19,   -19,     0,     9,    19,     7,    -4,     4,   -31,     3,     3,    -9,    -4,    17,     2,   -14,   -11,   -12,    -9,   -10,    -6,    12,     1,     7,    25,     2,     3,    12,   -21,   -12,    -2,    12,    10,    -4,     5,     0,   -14,     2,     3,    -1,    13,     0,     4,    -7,   -12,    -9,     1,     8,     2,    -8,    13,     1,     5,    27,     1,    10,    -4,   -18,    -2,    -2,    11,     0,     0,    -5,   -13,     3,     1,    -3,     4,    -9,     5,   -19,   -16,   -17,    -3,     0,    12,   -11,     5,   -11,    11,     6,     4,    20,     7,    -3,    -8,     8,    13,    -1,    -4,    -1,   -11,    -4,    -4,    -4,    16,     2,    -3,   -20,   -25,   -21,    -2,     2,    -2,    -6,     0,     6,    14,     2,     4,    19,    20,    13,     6,    -1,   -16,    -9,     5,   -22,    -2,     1,    -6,    -3,   -12,   -10,   -14,    -6,   -28,   -25,   -10,     4,    -9,    -9,     7,     5,    15,     9,    20,    18,   -13,     0,   -12,   -29,   -14,   -11,    10,    -8,     0,    -4,     4,    -3,   -12,    -4,   -14,    -1,   -14,   -12,     4,     0,    -1,     1,    16,     7,     9,     6,   -12,   -16,    -9,     1,    -7,   -17,   -14,   -13,   -10,    -5,     2,    -2,    -4,    -1,   -14,     0,    -8,   -20,   -11,     3,    -1,    -9,   -14,    -1,    12,    -9,     6,    -5,   -10,   -27,     2,    -2,   -14,   -21,   -23,   -25,    -9,     0,     4,     1,     4,     1,    -7,   -10,     0,    -7,   -14,    -9,   -10,    -5,   -14,    -1,   -21,   -13,     7,   -14,   -28,   -13,   -11,    -9,    -2,   -14,   -15,   -19,    -1,    -6,    -3,    -2,    -4,    -5,    -5,    -3,    -6,     2,    -1,    -7,    -3,   -15,    -7,    -3,    -5,   -10,    -4,    -2,    -5,   -10,   -22,   -13,    -6,    -3,    -4,    -2,     2,     2,    -4,    -3,     1,    -5,     4,    -5,    -6,   -12,    -8,    -5,    -8,     1,    -6,    -8,    -6,     1,     0,    -2,     2,     1,    -5,   -18,    -7,     0,     6,    -4,    -2,    -2,    -1,    -5,     4,     2,     4,    -5,     0,    -2,    -1,    -5,     3,    -5,     0,    -1,    -1,     2,    -1,     3,    -5,    -3,     1,   -10,    -5,    -3,     1,    -1,     0,     0,    -2,    -5,    -3,     4,    -5,     0,     0,    -2,    -4,    -5,    -2,    -6,    -4,    -2,    -5,     0,    -4,    -1,    -3,    -3,     3,     3,    -5,     0,     2,    -2,     4,    -4,     1),
		    57 => (   -2,    -4,     4,    -3,    -4,     3,    -4,    -4,    -3,     1,    -2,    -1,     2,    -3,    -3,    -4,     5,    -1,     0,    -2,     1,    -1,    -2,     0,     3,     3,     0,     5,     1,     1,     1,    -2,     3,    -4,     4,     2,    -3,    -2,    -2,   -19,   -22,   -19,   -13,   -42,   -50,   -53,   -11,     2,    -5,     0,    -3,     0,    -3,     1,    -4,     0,    -3,    -3,    -2,    -5,     3,     3,    -9,   -10,   -30,   -31,   -45,   -41,   -25,   -15,   -12,   -27,   -21,   -12,   -15,    -1,   -25,   -22,   -19,   -17,   -16,    -7,     2,     2,    -1,    -2,    -3,   -12,   -10,   -33,   -53,   -53,   -47,   -31,   -47,   -69,   -69,   -49,   -45,   -42,   -29,   -20,   -18,   -33,   -16,   -26,   -75,   -49,   -23,   -12,     1,    -4,     2,     2,    -3,   -20,   -22,   -38,   -51,   -71,   -78,   -93,  -100,   -16,    -4,    -8,   -13,   -23,   -53,   -73,   -60,   -40,   -30,   -27,   -46,   -62,   -62,   -35,    -8,     3,     5,     4,     2,   -27,   -38,   -15,   -30,   -20,    -5,    13,   -12,    12,    20,    18,     0,    -6,   -12,   -37,   -50,   -64,   -66,   -41,   -42,   -91,   -67,   -59,    -5,     2,     1,    -2,   -14,   -12,    -9,    13,    10,     9,     2,     9,    27,    26,     2,     5,   -22,   -10,    10,   -14,    -4,   -27,   -34,   -17,   -28,   -31,   -40,   -42,   -26,   -19,     3,    17,   -14,     4,    -4,    36,    22,    24,    19,    22,    28,    -1,    10,    16,    15,     3,    13,    18,    24,    12,    -8,    -5,    -6,   -12,   -30,   -64,   -40,   -25,   -18,    11,    -3,    18,     0,    30,     2,     9,     5,   -11,    15,    18,   -22,   -27,   -18,    11,    18,    11,    18,    14,    14,    12,    -7,    -1,   -29,   -37,   -38,   -17,    -4,    12,    14,    13,    18,     2,    -7,    -3,    -2,    -7,     4,    14,    -5,   -10,   -24,     2,     4,    24,    21,     6,     0,    20,     7,    16,   -29,    -6,    36,    50,    -3,    23,    -3,   -12,    11,   -25,     3,   -14,     5,     7,     1,    10,   -17,   -24,    -4,     3,    19,    19,    25,    15,    14,    -5,    17,    -6,    -4,    19,    32,    43,    -2,    -1,     0,   -11,    15,    13,   -18,   -11,    -3,    15,     6,   -18,    -7,    19,    -6,    -1,    17,     9,    21,    13,   -14,     4,    22,    18,    -8,   -31,    -2,    28,    -3,    13,    19,     2,    20,    29,     2,   -19,    19,    -7,   -21,    -7,    -7,    -7,    -6,    22,    17,    20,     9,     2,    -3,     6,     1,    11,     4,    16,    29,    45,     0,     7,    27,     0,    20,    24,    -7,   -10,     8,     1,    -1,    -3,   -13,     1,   -13,     7,     3,     3,    -2,     4,   -10,    -5,    23,     8,    22,    24,    -5,   -13,    -1,    11,    10,     4,     1,    18,   -18,    12,    10,    -5,    -1,    -5,     3,   -12,    -9,     1,   -11,    13,    -1,    11,    -7,   -10,     6,   -10,    -6,   -48,   -44,    -7,     4,     0,    -5,    -2,   -10,   -15,     1,     6,     5,    11,    13,     6,    -6,     2,    12,    18,   -10,     2,     9,    10,    -4,    -1,   -14,   -29,   -41,   -49,    -5,   -33,     2,     0,    -7,   -23,     5,    13,   -13,   -16,    -9,     8,    10,     1,    10,    27,    17,    39,     9,     5,     2,   -11,   -18,   -11,    -4,    -9,   -18,   -45,   -34,   -33,    -4,    -5,   -18,   -34,     9,     5,    -3,   -18,   -16,   -34,    -9,   -13,    19,    23,    17,    16,    -3,   -11,   -15,   -13,    -9,    -7,     0,    -2,    21,   -26,   -14,   -35,     7,     3,    10,   -57,     2,    -6,   -22,   -17,   -16,   -18,   -14,    -2,     4,     6,    10,   -11,   -31,     2,    -1,   -14,    23,    22,     6,    23,     7,   -41,     5,   -23,     5,     6,    -3,   -22,   -16,    -3,   -11,   -26,    -1,   -14,   -19,    -4,    11,    16,    -5,   -33,    -3,     1,    -4,    -4,     8,    27,    -9,   -21,    16,   -43,   -38,   -13,    -2,    -2,   -11,   -12,   -45,   -34,   -26,   -18,   -34,   -12,   -32,   -30,   -14,     8,     4,   -17,    -4,     2,   -36,    -3,     4,     7,   -17,   -42,   -17,   -37,   -32,     3,    -3,     1,   -17,   -31,   -42,    -5,   -10,   -10,   -13,   -30,    -8,   -11,    -9,     8,   -11,    -6,     5,     0,   -28,   -13,   -16,    21,   -16,   -37,   -53,   -14,   -10,     0,    -7,    -7,   -23,   -29,    -2,     5,     0,   -11,    12,    -1,   -12,    -5,     5,   -13,    -1,     2,    23,    -3,    -6,     7,    21,    -2,   -23,   -95,   -51,    -5,   -16,     0,     2,    -5,   -18,   -34,     6,     8,     8,     6,    21,    11,     0,     9,    27,    16,    32,     5,    17,    15,     1,     0,    15,    -4,   -23,   -83,   -45,   -23,   -38,    -2,    -4,     3,    14,   -11,    32,    32,    32,    29,    28,     2,    15,    22,    25,    51,    44,     3,    29,    21,     4,    17,    16,    10,    -6,   -58,   -31,   -33,   -25,     3,     0,    -3,    -4,    13,    14,    19,    16,    18,    16,    21,    37,    35,    27,    23,     9,   -13,    44,    17,    12,    13,    -1,    23,    26,    -8,    -8,   -26,   -18,     3,    -1,     3,     4,   -17,   -14,   -24,     2,    18,    18,    28,    29,    30,    28,   -24,   -43,    -4,    18,     3,     8,    27,    15,    22,    28,    10,   -12,    -3,    -4,    -1,    -2,     3,    -3,    -1,    10,    11,    -7,   -12,    -1,    13,    22,     4,    -2,   -33,    -7,     8,   -13,    15,     9,    11,     7,    23,    11,    30,     2,     0,    -4,     1),
		    58 => (    2,    -2,    -1,     1,     3,    -4,    -3,     5,    -2,     2,    -4,    -5,    -2,    -4,     1,     2,     1,    -4,     4,    -2,     3,     0,     5,    -1,     0,     0,     0,     5,     1,     1,    -3,    -4,    -4,     3,     1,     1,    -2,     2,     5,    -7,   -14,    -8,   -10,    -6,   -15,   -15,   -16,    -7,     3,     3,    -3,     5,     1,     4,    -2,     3,    -3,    -4,    -3,    -1,    -2,    -4,    -8,   -11,   -30,   -30,   -42,   -21,    -3,    -3,   -17,   -17,   -25,     6,     3,   -14,   -14,   -14,   -13,    -5,    -5,    -4,    -1,    -3,    -1,    -1,    -8,   -11,    -7,   -16,   -32,   -60,     6,    15,    14,    -3,   -16,   -20,   -14,    17,   -18,   -24,     4,   -15,   -12,   -14,    14,    27,     1,   -10,   -15,     4,    -2,   -15,   -13,   -37,   -31,   -35,   -19,    20,    45,    38,    30,    15,    -5,    -3,    13,    15,    12,    31,    -6,   -20,   -26,   -32,   -15,   -27,   -35,     3,    18,    -7,     2,     4,   -26,   -31,   -25,   -37,    -3,    50,    18,    22,    13,    26,    28,    12,     3,     8,    14,    28,    -2,    30,    -2,     5,    12,    -9,   -12,    -9,   -26,   -10,     2,    -5,   -40,   -33,   -35,   -18,   -12,    23,   -10,     2,    20,     4,    -3,     8,    -4,     9,    -2,    -7,     8,     8,    19,     1,    -3,    14,   -10,   -17,    -8,    -6,     2,   -27,   -33,   -39,   -33,   -25,    -1,     3,    -4,    -2,    -4,    21,     0,     6,   -19,    14,     7,    -4,    -6,     5,   -12,    -5,   -10,    37,    22,   -37,   -25,    12,     9,   -19,   -29,     4,    -4,    -3,    -5,    20,     8,     4,     5,     1,    -4,     4,    -2,    -4,    -6,    -2,    14,    33,   -13,    28,    22,    35,    38,   -22,    32,    36,     3,    -9,   -37,     9,    20,   -11,     1,    18,     9,     0,   -13,     0,    -3,     0,    11,    -6,    -7,    10,     4,    -4,    23,    21,    22,    16,     7,   -10,    32,   -41,    -3,    -3,   -45,   -30,    41,    12,   -15,    14,    14,     7,    20,     7,     8,    -5,    19,   -33,   -25,     3,    -5,     1,     6,    24,    11,    23,    17,   -33,    13,   -16,     3,    -5,   -21,    -1,    38,    33,     8,    22,     7,     2,     8,     0,   -10,   -10,     7,   -29,   -26,   -19,     2,    -1,    10,    15,    17,    21,    25,     8,    38,    -8,    -2,     3,   -31,     8,    37,    65,     2,     3,    23,    10,    -1,   -13,   -21,   -20,    -3,   -15,     1,    -2,   -16,   -10,    13,    14,    34,     4,    15,   -15,    19,   -35,     5,    -3,   -19,    -2,    13,    36,    12,     6,    16,     2,    -2,    -5,    -5,    -8,    -5,     6,     1,   -26,   -13,   -10,    17,     7,    29,     2,   -19,   -21,    15,     5,     1,    -8,    -8,   -24,   -35,     5,    23,   -31,    17,   -41,   -28,    -8,   -16,   -18,     1,     4,   -11,   -28,     1,   -24,   -33,    10,    -2,   -10,   -27,    -4,   -17,   -11,     3,     3,   -14,    12,   -59,   -14,   -19,   -23,    10,   -24,    -8,    -8,   -28,     3,    10,   -16,   -12,     3,   -22,    -9,   -16,   -26,    -8,   -33,   -42,   -10,   -45,   -27,     3,    -5,    -8,    16,   -56,   -24,   -29,   -46,   -25,    -2,   -29,   -20,    -3,    15,    -2,    -9,   -21,   -39,   -19,    -2,   -21,   -30,   -16,   -10,   -16,   -16,   -51,   -27,     1,    -5,   -12,   -27,   -15,   -28,   -32,   -30,    -4,   -20,   -19,   -32,    -8,   -10,   -16,   -30,   -14,   -12,   -14,    -7,     3,    -7,    -8,    -5,    -5,   -49,   -24,   -38,    -6,    -7,   -18,   -51,     0,   -28,     1,     9,     4,    -4,   -10,   -13,     5,    -2,   -18,   -54,    -2,     5,     1,     9,    -5,    -9,     2,    -1,     2,   -46,   -20,   -25,     3,     2,   -38,   -47,   -11,   -28,   -18,     8,    30,     8,     5,   -11,   -20,   -18,   -32,   -22,    -6,    23,     2,    10,    11,   -16,     7,    23,    30,   -60,   -45,   -30,     2,     1,   -14,   -39,   -30,     6,    15,     4,    26,   -10,    27,    -1,    14,     1,   -20,    -7,    24,    16,     4,     1,    20,    21,    19,    49,    11,   -73,   -46,     2,   -12,   -20,   -18,   -21,   -25,     5,    33,     4,    21,    33,    15,    13,     8,    18,    15,    39,    -2,    27,   -28,    12,     2,     3,    37,    32,   -13,   -56,   -35,     0,   -13,   -17,    -9,   -17,    15,    33,    20,    30,    27,    26,    37,    36,    17,    27,    46,    47,     7,     6,    11,   -10,     0,     1,    31,    18,   -18,    -3,   -35,    -3,    -4,     3,    -5,    -9,    32,    -3,    12,    -7,    14,    15,     4,     5,    30,    30,    30,    33,    30,    25,    30,    42,    10,   -12,    43,    22,   -11,    -4,   -35,     0,     4,     1,   -14,   -21,   -13,   -14,    -8,   -11,    12,    21,    10,     4,    28,     9,    13,    20,    43,    -5,    -2,    -6,     4,   -21,     6,     7,   -20,   -48,   -25,    -4,     4,    -1,   -15,     2,   -59,   -47,    -3,    -4,   -20,   -35,   -19,   -20,   -12,   -10,    13,    16,    -5,   -11,     9,    -5,   -34,   -31,   -32,   -17,   -19,   -12,    -7,     1,     1,     2,     1,   -13,   -27,   -47,   -44,   -10,     8,     3,   -23,   -12,    11,     7,   -38,   -81,   -37,   -22,   -19,   -60,   -51,   -24,   -28,   -10,    -2,     2,     0,    -3,     0,     1,    -2,     3,   -12,   -10,   -13,    -8,   -16,   -15,    -3,    -5,   -20,   -33,   -39,   -31,   -16,   -25,   -13,   -14,     0,     0,   -10,     0,    -1,    -4,     1,    -1),
		    59 => (    4,    -3,     4,    -1,    -4,     4,    -3,    -3,     5,     0,     4,    -3,     2,     2,    -2,    -4,    -3,    -5,    -3,    -2,     5,    -2,    -5,     5,     5,     4,     3,    -3,     2,     4,     1,    -4,    -4,     4,     1,     0,    -5,    -2,     1,    -6,    -8,   -11,     4,    -6,    -3,    -8,    -1,     4,     2,     4,     2,    -4,    -3,    -4,    -5,     4,    -2,    -4,     2,     4,    -5,     3,    -4,    -3,    -8,    -5,    -2,    -8,    -4,    -4,   -15,    -5,     4,    -4,     2,    -4,    -4,     3,    -2,     1,    -3,    -3,    -1,     3,    -1,    -2,     3,    -4,    -7,   -10,    -8,    -1,   -13,   -20,    -6,   -16,    -5,   -21,   -14,   -16,    -4,     3,     8,     1,   -20,   -15,    -6,    -6,     1,    -6,     1,     5,     4,    -1,     3,    -1,    -2,    -5,   -20,    -7,    -6,    -1,   -10,     1,   -28,   -38,   -32,   -26,   -22,   -21,   -11,   -28,   -31,     0,    -4,     0,    -3,   -21,   -17,    -5,    -4,    -1,     0,    -2,    -5,     2,    -4,   -13,   -40,   -15,   -19,     2,     6,     0,     7,    -1,    -9,   -31,   -39,   -22,    -4,    -6,     0,    -2,     2,   -20,   -10,     3,    -2,     3,    -6,    -3,   -14,   -22,   -19,   -30,    -7,    13,     3,    23,    23,    19,    -2,   -11,    15,    -6,   -50,   -46,   -22,     1,     2,    -3,     0,     1,    -3,   -14,    -5,     0,    -6,     3,   -10,   -24,   -37,   -28,    -2,   -17,     6,    21,     2,    10,   -11,   -31,   -24,   -25,   -54,   -69,   -24,     5,    -1,     1,    -9,     0,    -5,   -11,   -10,    -5,   -10,    13,     4,   -25,    22,    -6,    18,     2,    -2,     4,    -7,     3,    -6,   -23,   -26,   -14,     7,   -17,   -37,    -7,    -6,    -9,   -11,    -3,    -2,    -1,    -3,   -18,   -16,     7,    -2,   -16,    16,    15,     7,    13,    21,   -11,   -12,     5,     4,   -20,   -31,    14,    13,   -13,   -24,   -19,   -23,   -10,   -18,   -24,   -11,   -11,    -2,    -6,    -8,     7,    -5,   -25,    22,    12,     9,     4,     2,   -42,   -37,     7,    25,    -5,    14,    -1,    -1,   -12,   -22,   -24,   -27,   -18,   -16,   -19,    -3,   -18,    -3,   -27,   -11,    13,   -12,   -28,    10,    23,    17,     5,    -8,    -4,    15,    51,    -2,    -5,    -4,    18,    -7,    -3,   -36,   -41,   -26,   -24,    -9,   -17,     1,   -16,     4,   -10,   -11,    17,    -9,     9,     9,    -4,    -2,    20,     9,     4,    17,    34,   -13,   -28,    -6,    15,     0,    -1,   -14,   -22,   -36,   -27,   -16,   -13,   -15,   -18,     3,   -11,    -9,   -14,   -17,     1,    43,     6,   -20,     3,     7,    -9,     0,    -6,    -9,    -6,    -2,    -4,   -16,     9,   -16,   -21,   -20,   -20,    -9,   -11,   -13,    -1,    -4,    -2,    -8,   -10,   -12,   -11,    28,     3,   -11,    -9,    22,    -1,   -16,   -10,     7,     8,    -6,     1,     1,     0,   -15,   -27,   -29,   -29,   -13,   -21,    -1,    -2,    -5,    -1,    -8,   -11,    14,   -19,   -18,     4,    -6,   -14,    11,     4,   -10,   -29,   -13,     7,     8,    -1,    -7,    -7,   -45,   -40,   -28,   -26,    -8,    -5,     0,   -13,    -4,     0,   -14,    -2,    -1,   -12,   -43,    -4,     8,   -16,     5,    47,    17,     7,     3,   -20,   -17,   -17,    -6,   -17,   -59,   -22,   -12,    -9,    -8,    -6,     1,   -21,    -2,    -2,   -18,     2,    -1,   -16,   -34,   -40,    -4,   -30,   -11,    13,    23,    15,     3,     2,   -23,   -25,   -16,   -13,   -38,   -24,    -9,   -14,   -22,    17,   -15,   -10,    -5,     0,   -16,    -1,     1,     0,   -10,   -25,   -32,   -31,   -32,   -13,    17,    -9,    -8,   -11,    -6,    -1,   -23,    -8,   -16,   -27,     1,    -9,   -26,    -3,   -13,   -10,    -5,    -1,   -13,    -3,     0,    -8,    -4,    -1,    -7,    -5,   -26,   -41,   -39,   -37,   -28,    15,     8,     3,   -15,   -15,   -25,   -28,   -14,     0,   -18,    18,   -13,   -11,    -2,    -6,    -1,    -8,    -2,    -1,    -2,   -20,    -1,   -20,   -22,   -36,   -47,   -29,    -2,     4,    -4,    -6,   -13,   -14,   -11,    -9,   -11,   -12,     4,    12,   -16,     1,     3,    -5,     2,    -7,    -4,    14,    -6,    -7,    -3,     3,     5,    -5,   -12,    -5,     5,   -16,    -3,     1,    -1,   -26,   -10,   -17,    -9,    -4,     9,    19,   -22,    -5,    -1,    -3,    -7,    13,     0,     5,     9,     8,     9,    15,    -7,     5,    15,     7,     6,    10,    -3,    10,    -6,   -24,   -16,   -27,    -6,     0,     7,    -5,    -1,    -3,     4,     3,   -11,     6,    -4,    -4,    10,    -2,     8,    -7,     5,    -6,     0,    -2,    -3,    15,     1,     9,    14,   -10,   -11,   -13,    -3,    10,     6,     5,   -11,     0,    -1,    -1,    -2,    -2,    -5,     3,     0,   -14,     2,   -10,    12,   -12,   -34,   -26,    -8,     7,    12,     9,    10,    12,    10,     2,    -3,     7,     5,     7,    -3,     1,    -1,    -2,     9,    -2,    -3,     2,     2,    -8,    -6,     7,   -16,   -21,   -13,     5,   -25,   -20,     4,    19,     6,   -21,   -25,   -22,   -19,    -9,    -7,     7,     2,     4,     2,    -3,     3,     9,     1,     0,     1,     2,     5,    13,   -10,   -22,    20,     2,    20,    11,     7,    45,    17,   -21,     4,     2,    -4,     7,     7,     3,     0,    -5,    -5,    -3,     0,    -3,    -3,    -5,     9,    12,     6,   -15,    -7,     5,    -2,   -15,   -19,    36,    34,    -3,    -8,    17,     7,   -14,   -11,    -3,    -2,    -1,     4,     1),
		    60 => (    1,     0,     3,     3,     4,     0,     4,     4,    -1,     1,     2,     5,     0,    -1,    -4,     3,    -1,    -4,    -4,    -4,     3,     3,     0,    -4,     0,     1,    -1,     5,     0,    -2,     4,     1,     0,     2,    -2,   -11,    -9,   -12,   -22,   -10,     3,     6,   -29,    28,    34,    35,     1,    -5,    -7,    -6,     3,    -1,     3,     3,     0,     0,    -1,    -4,     4,    29,    36,   -10,   -16,     5,    -7,   -20,   -32,   -27,   -34,   -66,   -34,   -16,    -2,   -25,   -17,   -18,   -19,   -16,   -46,   -18,   -22,    -4,     2,     4,     3,    -3,     4,    31,    10,   -30,   -35,   -30,   -29,   -24,   -16,   -37,   -52,   -24,   -28,   -31,    12,    13,     0,   -24,   -24,   -35,   -50,   -25,   -19,   -21,   -37,     4,     0,     0,    -3,    -9,   -12,   -61,   -22,   -26,     3,    27,    -3,     5,   -29,     0,   -11,    11,    27,    13,    -2,     1,   -22,   -22,    -9,   -13,   -41,   -70,   -29,     2,    -1,    -5,   -16,   -10,   -14,   -31,    14,    -6,     6,    39,    24,    21,     5,     3,    17,    15,    16,    17,    15,     1,    -2,    -4,   -17,   -12,   -39,   -61,   -14,    -7,     2,     1,   -22,    -2,   -40,    11,    24,    24,    21,    15,    26,    12,     3,     2,    14,   -14,     6,    -5,   -20,     7,    -4,   -24,    -1,   -46,   -26,   -70,   -20,    -7,    -1,   -10,   -19,   -22,   -23,    -1,    22,    21,   -11,    11,    -7,     4,     7,     8,   -22,   -25,   -11,    -6,    -8,   -22,    -7,   -20,    -5,    -1,   -24,   -13,   -36,     6,    45,   -28,    -2,   -31,   -29,     2,     3,   -23,     4,     8,   -11,   -22,     2,    -6,   -37,    -3,    -8,    18,    -3,   -11,   -12,     5,     0,    17,   -29,   -67,   -35,    -8,    -6,    -8,    17,    -1,    -7,     8,   -23,   -12,    -5,    10,    -9,     8,    19,     7,     8,    17,    12,    16,     8,    11,     8,    -7,    -1,    17,    -7,   -41,   -11,    -8,    -7,    -6,    21,     8,     3,   -14,    -6,   -14,     4,    14,    -4,    -6,    -1,    15,    46,    34,    31,    37,    -6,    14,     9,   -13,     7,    18,    -1,   -24,   -30,     0,    -3,    49,   -30,    -4,    -9,   -29,   -10,   -15,   -19,    -9,   -14,    -3,    12,    54,    20,    25,    60,    46,    40,    24,    19,    10,     9,    12,    29,   -29,   -30,    -3,    -4,     1,   -30,   -10,    16,   -29,   -26,   -31,   -25,    -5,   -11,     3,    29,    41,    28,    34,    24,    22,    23,    15,   -11,     1,    -2,     8,    15,   -14,   -24,   -16,     1,     4,     0,   -13,    21,    -4,     2,   -17,    -5,   -20,   -15,     9,    11,     3,    -2,     5,     1,    -9,    -5,    -8,   -10,     7,     5,    24,     8,    13,   -42,   -15,    -4,     0,    -5,   -39,   -14,    -7,   -18,    -5,    -1,   -12,   -12,     1,   -12,    -8,   -38,   -44,   -44,   -19,    11,    -8,    17,    36,    36,    20,    34,    29,   -36,    -4,    -3,     3,   -25,   -36,    -7,   -17,   -23,    10,    -1,   -27,   -24,   -18,   -28,   -27,   -59,   -34,   -23,    -7,   -14,    -2,    21,    15,     4,    15,    25,    31,   -39,   -34,    -5,     1,   -14,   -17,    14,    -9,   -25,     6,    -5,   -14,     1,   -13,   -23,   -32,   -34,    -4,   -28,   -24,    -9,    15,    13,    -8,   -13,   -22,    -4,   -11,   -55,   -12,     1,    -3,   -19,     1,     6,     4,   -15,    10,    -5,     6,    12,    18,     8,    20,   -13,   -13,   -21,    -5,    -5,    13,    -4,   -32,    -8,   -11,    -6,   -35,   -35,    10,    -3,    -1,   -16,   -12,    19,    17,    13,    -8,     5,    20,    22,     9,     3,   -13,   -26,    -9,    -9,     7,     6,     5,   -24,   -19,   -11,    12,   -30,   -33,   -27,   -19,     4,     8,    -5,   -10,     1,    27,    17,    30,    22,     6,     0,     5,    23,   -10,   -15,     0,    -2,     3,     3,    25,   -12,   -18,    -5,    12,    -1,   -54,    -7,    -5,     1,     8,   -23,   -18,    29,    19,    14,    24,    13,    35,     0,    11,    34,    10,     2,    12,     0,     9,    -2,     5,   -22,   -27,   -13,    -8,   -19,   -63,     5,     2,     3,    -4,   -24,   -14,     2,    -4,    25,    35,    29,    21,    14,     4,    20,     2,    -6,    13,     8,     0,     8,     7,   -10,   -19,    -3,     4,   -32,   -31,    62,     0,    -3,    -2,   -13,   -14,   -42,   -23,    -5,    34,    26,     4,    36,    17,    -4,   -12,     9,    23,    14,    10,    -9,    -8,   -24,   -25,   -10,    -2,   -22,   -13,    38,     7,     2,     4,   -12,   -28,    -9,   -27,   -22,    -3,    24,    19,    14,   -17,    18,    -6,     5,    11,     9,    25,    -6,   -27,   -43,   -29,   -36,   -11,   -24,   -33,   -32,    -5,     5,    -3,    -9,   -15,     8,    16,   -27,   -16,   -15,    -8,   -14,   -45,   -29,   -27,   -26,    15,    -5,    -1,   -16,   -39,   -22,   -40,   -34,   -25,   -21,   -11,    -3,     0,     3,     3,    -4,    -9,   -39,   -24,   -43,   -65,   -36,   -38,   -41,   -24,   -38,   -22,   -26,   -33,   -72,   -62,   -62,   -70,   -49,   -56,   -40,   -18,    -4,    -1,     4,     4,    -1,     0,    -2,     1,   -13,   -39,   -55,   -26,   -21,   -38,   -27,   -30,   -20,   -24,   -30,   -49,   -41,   -37,   -36,   -44,   -39,   -46,   -28,   -19,   -11,    -2,    -2,     0,     0,     1,     0,     1,     0,     1,    -3,    -7,   -12,   -22,     1,    -2,     0,   -29,   -10,    -5,    -1,     3,   -16,   -15,   -12,   -22,   -11,   -17,     1,     3,    -4,     5),
		    61 => (   -2,    -3,     3,    -1,    -4,     3,    -4,     3,     0,    -2,    -4,     1,     1,     2,    -4,     0,    -4,    -4,    -2,     3,    -3,     0,    -1,    -4,     1,     5,    -2,    -2,     5,     0,     1,     0,     0,     2,     0,     1,     1,     2,    -1,    -2,    -8,    -8,     7,     2,    -7,    -5,     0,     4,     4,    -3,     0,     2,     4,     1,     3,     4,     0,     3,     3,     1,    -3,    -3,    -2,     4,    -3,    -4,    -1,    -1,   -19,   -19,   -18,   -39,   -39,   -17,   -11,    -2,    11,   -13,    -9,    -3,   -11,   -10,     3,    -2,     2,     1,    40,    27,     5,    -7,     1,    16,     6,     4,    -6,    -4,   -31,   -79,   -60,   -47,   -32,   -29,   -19,     0,    -2,    -5,    45,     8,    -3,   -12,    -2,     5,     5,    -4,    34,    28,    12,   -10,   -19,   -11,   -30,   -14,   -26,   -29,   -50,   -54,    25,    12,    19,    14,    11,    10,     2,    12,    12,   -15,   -26,   -31,   -26,   -22,     4,    -4,    26,    39,    24,     7,    -8,   -14,   -59,   -36,   -56,   -53,   -52,   -31,     1,    12,    -8,   -14,   -34,   -18,    -8,    10,    22,    -1,   -20,   -33,   -29,   -28,    -2,    -1,   -21,    17,    34,   -17,    24,    37,   -23,   -55,   -62,   -59,   -30,   -11,    -2,   -11,    -7,     3,   -13,    -8,    12,     0,     2,    -6,   -26,   -26,   -16,   -15,    -5,   -29,   -35,    -6,   -23,    26,    28,    34,   -41,   -41,   -90,   -51,   -28,   -12,    -2,     2,    14,    12,    -1,    18,    21,     4,   -18,   -11,   -30,   -21,   -18,   -13,     0,   -28,   -29,    10,   -22,    19,    24,     8,   -26,   -30,   -38,   -44,   -50,   -24,    -2,    14,    13,    12,     5,    11,    10,     3,   -13,   -23,   -42,   -17,   -35,    -5,     3,    -3,   -27,     6,   -13,   -18,    21,    31,    18,     7,    -8,   -50,   -15,   -38,    -3,    23,    38,    10,    14,     3,    -4,   -15,   -14,   -11,   -26,    -8,    -2,   -10,    -4,    12,   -29,   -10,   -14,   -26,    -1,    24,    -9,    -6,    16,    -5,   -17,   -32,    -2,     8,    14,    11,    -7,   -14,   -36,   -48,     2,    -4,   -23,    -1,     0,    30,     2,     2,    -6,    14,    -2,    23,    16,   -33,   -45,   -17,    11,   -12,   -46,     1,     5,    11,    10,     1,   -16,   -41,   -15,    -9,     1,   -10,    -6,     0,     1,    24,     0,     3,   -13,    23,    -6,    30,    28,   -10,   -17,     3,    -4,   -17,   -13,    11,    20,     5,    10,    13,   -24,   -33,   -10,    24,    -7,   -13,   -21,    17,    -2,    21,    -3,    -1,    -7,    16,     9,    12,    24,     7,    15,    17,    -9,   -22,   -19,     0,    21,    -2,     5,    22,   -41,   -67,   -36,    20,   -15,   -17,   -23,     1,     4,     4,    -3,    -1,    15,    10,    33,   -16,   -18,   -50,    15,    -2,     4,   -13,   -14,     8,     8,   -11,    13,    -9,     3,   -31,   -21,    34,    20,    -3,   -11,    27,    32,    -1,     2,     0,     3,    34,    16,   -39,    -2,    -6,    17,     2,    -8,     9,    -2,     7,   -14,   -13,    23,    16,   -45,   -48,   -15,     4,    -2,   -18,   -23,    15,    15,    -7,     0,     5,    15,    -7,    -2,     3,     0,   -28,     2,    -1,   -35,     6,   -12,    12,    -5,    -4,    23,     4,   -26,   -49,   -27,    12,     1,    13,    16,     7,    -1,    -7,    -5,     3,     2,   -29,     8,    -3,     5,    -9,   -13,   -16,   -24,    17,     3,    11,    -4,   -19,    -5,   -39,   -34,   -26,   -19,     6,   -12,     1,     9,    15,    -4,    -4,    -5,    -2,    -5,    -7,   -11,   -38,   -28,   -29,    -6,     0,    -5,     8,     4,     9,    -6,   -15,   -35,   -34,   -22,   -32,   -28,     4,     1,    15,     5,    17,     2,    20,    -4,    -3,    16,     9,    -1,   -31,   -10,   -19,    -4,    14,     3,    10,    -5,    12,    -1,     3,   -25,   -17,   -10,   -31,   -23,    -3,   -18,    17,    24,    28,     6,    18,     0,     0,    16,    -2,    15,    -8,    -5,   -16,     0,   -15,     3,     1,   -10,     8,    16,    -7,    -3,   -30,    -2,   -11,    18,   -10,    -5,    11,    35,    30,     4,    -3,    18,    24,    19,    15,     8,    21,   -13,    -3,     1,   -10,     8,   -17,    -1,     1,     4,     4,   -19,   -39,    -1,    14,    33,    11,    -3,    18,    30,    16,     1,    -2,    15,    23,    15,    14,    -5,     9,     4,   -25,   -21,    -7,   -17,   -17,    -2,    -1,    19,    32,    14,     3,    35,    16,     1,    -5,     6,    22,     4,    -4,    10,     1,     5,     4,    -1,    -4,    -7,    -5,    19,    27,    34,    37,    -4,    -8,    -4,     8,     9,    39,    16,    25,    19,    -3,   -30,   -31,    -8,    -9,    12,    27,    40,    -4,     2,     1,     2,   -10,   -37,   -35,   -32,    -4,    -3,    35,   -13,   -10,   -11,     3,     2,    24,    -5,    -3,    -6,     7,    -2,    14,     2,   -15,   -12,    17,    12,     0,     3,     2,     4,    -8,   -19,   -15,   -12,   -52,    -2,    24,   -65,   -53,     0,    -6,    18,    -8,   -28,   -53,   -29,   -16,   -27,   -19,   -14,   -11,    -4,     3,     0,    -4,    -4,    -1,    -2,     2,    -7,   -18,   -39,   -49,   -43,   -44,   -17,   -24,   -42,   -43,   -23,   -12,    12,   -26,    -2,    -7,    -4,    -8,    -1,    -1,     5,    -5,    -4,    -3,    -1,     3,     4,     0,     3,     3,    -1,    -3,    -2,    -7,   -21,   -18,    -1,    -3,   -16,    -6,   -10,     3,     5,    -4,     1,    -1,    -2,     1,     1,     2,     1,     4),
		    62 => (   -3,     2,     1,     2,     4,    -2,     1,     1,    -1,     0,    -5,    -2,    -3,     3,     8,     5,     4,    -3,     4,     5,     0,     3,    -2,     0,    -4,    -1,    -4,     0,     4,     2,    -2,    -4,     0,    -1,    -4,     3,     2,     8,     4,    -2,     0,     1,    -2,   -13,    13,     6,     1,   -21,    -5,    -5,     0,     0,     1,     4,     0,     4,     3,     2,    -3,     1,    -7,    -4,     5,    -2,     5,    -5,    10,    36,    28,    44,    18,    -6,   -12,   -14,   -25,   -62,   -46,   -11,   -10,    -4,     0,     7,    -1,     0,     0,    -3,    -5,   -17,   -16,    11,    25,    -3,    -6,    19,    -9,     5,    -8,     3,     0,     7,    21,     1,   -33,   -28,   -31,   -19,    17,     2,    -1,    -2,     4,    -1,     4,     4,   -12,    10,    12,    17,    43,    41,   -11,     3,    23,    24,    17,    37,    26,    23,     1,     4,     4,   -18,     6,    10,     6,   -27,   -30,   -10,   -18,    -5,     3,     4,     7,     2,    -5,   -18,   -14,    26,    -4,   -14,     9,     4,    14,    11,     1,    13,    14,    -2,     3,    -4,   -22,    14,    32,     4,   -15,   -17,   -20,   -10,     2,     1,    12,     8,    -8,   -29,     9,    11,    -6,     1,    -5,   -10,     0,    -6,    13,    -2,    -1,   -16,     7,   -21,     3,    13,    42,     9,   -15,   -22,   -11,    -6,    -3,     1,    -4,    21,    -1,    -9,   -29,    -2,    13,    -5,    11,    -1,     4,     9,    24,    18,    -2,   -12,   -13,   -26,     7,     0,    19,   -30,   -24,   -33,    -7,    -8,   -14,    11,    10,     3,    21,   -14,   -22,   -11,     7,     0,    20,    19,    -4,   -12,   -17,     4,     4,     2,    -5,    -1,     1,    -2,     4,     1,   -16,   -19,   -23,    -6,    -1,   -11,    38,   -10,    17,    22,   -27,     3,    -2,     1,    -2,   -17,     4,   -45,   -73,    -7,    11,     8,    -2,    -5,    -1,    -1,    -1,    14,   -34,   -18,    10,   -11,    -3,    -7,    22,     9,    -6,    -2,   -10,    25,     9,   -18,   -16,   -19,   -39,   -57,   -27,   -22,     3,     0,   -13,    -3,   -20,     7,   -34,    16,   -14,    -9,    14,    -6,     1,     1,    -9,    17,    19,    -7,     0,    -5,    -7,   -43,   -33,   -54,   -62,   -64,   -14,    -7,     1,   -19,   -24,   -19,    -7,   -11,   -16,    25,     1,     1,   -12,    -2,     3,    -3,   -13,    -8,    -2,    -5,   -18,   -53,   -42,   -49,   -48,   -37,   -46,   -17,    -2,   -18,    13,    -3,   -21,   -19,    -3,     1,   -15,    17,    -3,     8,    22,   -10,     1,     3,    16,     0,   -11,   -28,   -48,   -70,   -79,   -76,   -39,   -32,   -15,    22,   -12,   -14,    10,    -1,   -11,   -29,   -23,    -8,   -20,     4,    -9,    -2,    23,     3,     0,    -7,    -9,    -2,    -3,   -33,   -39,   -54,   -58,   -39,    -7,    -5,     2,     6,   -19,   -18,    -2,    -6,   -26,   -18,   -23,    -4,     1,    -7,    -8,     2,    15,    16,    -4,   -12,    -1,    -4,   -34,   -25,   -10,   -21,    -7,    17,    23,    14,   -11,     9,    -7,   -15,    -4,   -18,   -27,   -19,   -35,     4,    -2,   -11,    -5,    14,    16,    33,    -4,     0,    -2,   -14,   -29,   -19,     1,   -21,   -12,     8,     6,    10,     2,     3,     5,   -34,    -6,   -21,   -40,   -21,   -34,   -10,     1,    -2,   -10,    37,    17,    13,     2,     1,     3,    -4,   -24,    -7,   -27,   -13,    -4,     2,     4,    12,    19,    10,    -4,   -12,   -18,   -31,   -46,   -28,     4,    -1,   -26,   -26,   -19,    18,    -6,    14,     4,     3,   -10,     9,    23,    -6,    -5,    -7,    24,    15,     6,     7,    29,    -7,    -6,   -40,   -30,   -23,    -7,   -10,     3,     5,    -1,   -18,   -13,    49,   -18,    33,     3,    -4,     8,    22,    20,     3,    -2,    17,    32,    -7,    15,    14,    29,    16,   -20,   -14,   -22,   -32,    -9,    -3,     1,     0,   -23,   -29,    17,    18,    28,    36,     0,    -2,    23,    27,    27,    25,   -24,    11,    -3,    -3,     7,    14,    21,    11,    -1,    16,     3,    21,   -27,     4,     7,    10,    -1,    -4,    16,    19,    25,     5,    -2,    11,    28,    24,    18,    14,   -15,   -11,   -11,     7,     7,    -1,    14,    -5,    -1,     7,    16,   -13,     2,    24,     5,    15,    17,    16,    47,    53,    17,    -2,     1,    -2,    25,    24,     7,     0,    -5,     3,     9,   -11,    12,     4,     7,    -2,    15,    17,     4,   -38,    -9,    13,    17,    -6,    10,   -15,    -2,     7,   -21,   -11,    -4,    -2,    -4,     5,   -14,    11,    -1,     8,    25,    -2,    -5,    12,     0,   -12,    10,    26,     7,   -24,    18,     8,     0,    19,    13,    20,    17,    12,   -15,    -1,    -3,     0,   -17,    -9,   -18,   -29,   -49,   -71,   -45,   -19,     2,     6,     9,     9,    36,     3,   -17,     7,    23,    22,   -20,    13,    54,    32,    32,    12,    13,    -4,     1,    -3,    -7,    -5,    -8,   -15,   -12,   -24,   -45,   -46,    -9,    -3,    -8,    -1,    25,    29,    15,    42,    -4,   -41,     3,     9,     7,     1,    16,    15,    12,     4,    -3,     1,    -5,     1,    -2,    -4,   -13,   -11,   -13,    -6,    -4,   -20,    -1,   -27,   -27,   -18,   -44,   -30,   -21,    -9,    -4,    -3,   -15,     2,    -5,    -4,     1,     4,     5,     4,     2,     4,     4,     4,    -5,     3,     3,     3,    -4,    -3,    -2,    -4,     1,     3,    -4,    -4,     3,    -4,   -12,    -9,    -2,    -4,     1,    -3,     1,     4),
		    63 => (    3,     4,     4,     0,     1,     3,    -4,     0,    -2,    -4,    -1,    -3,    -3,    -2,    -1,    -6,     5,    -2,    -5,    -2,     1,    -2,     0,    -4,     2,    -4,     5,    -3,     5,     1,    -1,    -2,     3,    -5,     1,    -3,    -2,     3,    -4,   -10,    -8,   -12,   -14,   -12,    -7,   -22,   -11,    -1,     3,    -3,     4,     1,     0,    -1,     1,    -1,     3,     1,     3,    -3,     0,    -1,     0,   -10,   -36,   -33,    18,    16,   -13,   -26,   -36,    -1,   -12,    -9,    -5,    -7,   -26,   -20,   -16,   -19,    -9,     0,     0,     5,     5,     4,    -1,    -9,    -2,    10,    10,    27,    21,    -2,   -11,    20,    18,    15,    33,    11,   -18,    -8,   -15,   -12,     7,     0,   -43,   -64,   -32,   -23,     3,     3,    -3,    -4,   -16,    18,   -33,     4,    32,    12,     6,   -12,   -10,    -9,     4,    16,    25,     0,    -1,   -31,   -21,    -8,   -13,     9,     5,   -79,   -71,   -37,   -32,     4,    -3,     2,    -5,    -1,   -12,    -8,    16,     2,   -15,   -26,    -5,    20,    24,     4,     9,    -5,     9,     6,    -3,     9,    10,    37,    17,    25,    20,   -67,   -12,     3,     3,    -3,    13,     4,    15,    -7,     8,    23,   -29,    -2,     9,    27,    10,    10,   -15,   -15,   -10,     6,    11,     0,    29,    34,     1,    -5,    17,   -47,   -35,    -9,     3,     7,     2,    14,    45,    14,    31,    11,     3,    -2,     8,    23,    13,     2,    17,    15,   -25,    -8,     2,    22,     0,     6,   -27,    -5,     8,   -44,   -56,   -17,   -11,     0,     1,     6,    15,     6,    -8,   -15,     4,     3,     3,     9,    -2,   -15,    20,    11,     8,   -16,    13,    32,    15,    23,   -17,   -11,   -10,   -57,   -55,    -9,     3,   -19,    -5,   -10,    12,    11,    -2,    -9,     2,    -9,   -14,    -1,    -2,     8,    17,     9,    22,    17,    10,     9,   -10,   -13,   -10,   -14,   -66,   -70,   -65,   -23,    -1,   -25,   -17,   -16,    -5,   -19,   -22,    -3,    -9,     3,    -9,     2,    16,    14,   -14,     0,     8,    32,     8,   -28,    -5,   -46,   -25,    -6,   -44,   -33,   -50,   -21,    -4,   -23,   -26,     4,   -10,    -9,    -8,     9,    -1,   -15,    -1,     8,     2,   -12,   -14,   -13,    -1,    47,    20,     0,    -7,   -24,   -24,   -22,   -60,   -77,   -44,    -4,     0,   -15,   -32,     0,   -11,     3,    -5,   -16,   -10,    -3,    -1,     9,    22,    -1,   -11,    -6,    12,    27,    22,    25,    16,    -7,    -6,   -10,   -80,   -40,   -20,     0,    -3,    -9,   -24,     0,   -25,   -18,   -14,     0,    -1,   -22,   -10,    -2,    20,    -4,    -7,   -16,    30,    25,     5,    20,    12,     5,   -17,   -10,    -6,   -50,   -38,   -13,    -7,    10,    -1,   -11,   -24,    -3,     1,    -3,    -8,   -14,     3,    10,     5,    -5,   -15,    -9,     7,    28,    21,    36,    15,    24,    -4,    -4,    13,   -53,   -35,    -6,    -1,     8,    -1,     0,    -9,    32,    30,     1,    -1,    -9,   -18,    -3,   -15,    -3,   -19,   -12,     9,    14,    11,    23,    13,     6,    10,     7,    25,   -36,   -20,   -11,     0,     5,     1,    11,    -2,    10,    33,    17,    -8,    -1,    -3,     3,     6,   -13,   -17,   -18,    19,    29,    18,     7,    25,    20,    -4,   -14,    -1,   -49,   -53,   -19,    -2,    -1,    -2,    25,    -6,    -5,    29,    32,   -15,   -12,    -3,     2,    12,    -7,   -28,     3,    20,    19,    -5,   -13,    -4,    -4,    -8,   -11,   -54,   -50,   -24,    -6,   -13,     4,     7,    26,     2,    -5,    24,    11,     3,     8,    17,     8,    -1,   -31,    -9,    16,    17,     0,   -13,     0,     7,     5,   -12,   -20,   -48,   -50,   -12,   -13,     2,   -21,    -5,     1,    23,    24,    16,    27,    12,    11,    16,    -2,   -35,   -39,   -19,    -1,   -30,   -32,   -10,    -5,    -3,   -13,    19,     4,   -30,   -46,   -45,   -23,    -2,   -11,   -13,    -8,     8,    29,    18,    22,    -5,     7,    10,    14,   -36,   -30,   -19,   -19,   -35,   -37,   -20,   -12,   -14,   -29,    26,    -4,    -8,   -34,   -10,    -5,    -2,    -3,    11,     3,    -7,     9,    19,     3,    -5,     0,    13,    33,     6,   -26,    -4,     2,    -1,   -14,    -3,     6,    -7,     0,     9,    -2,   -24,   -37,   -17,     4,   -10,    -8,    16,     1,    -6,     9,    15,   -10,     7,    -6,    32,    37,    23,   -20,    -8,    20,     3,     5,    13,    -7,    -1,    -2,    23,   -10,   -48,   -31,   -26,    -4,    -1,     5,     6,     5,     0,     0,    -6,     4,     5,    20,    32,    39,     8,    25,    19,    26,    14,     9,    20,     2,    -5,     8,    -6,   -20,   -22,   -28,   -39,    -1,     0,     0,   -10,    25,     1,    -6,    -1,    23,    33,    34,    36,     4,     7,     9,    17,    19,    32,    11,   -11,   -18,     1,     5,    -6,    -1,   -44,   -33,   -17,    -4,    -3,     1,     3,   -14,   -13,    24,    21,    22,    24,    30,    17,    -5,     9,    -1,    14,    20,    24,    22,    14,    19,    21,    -1,   -22,   -60,   -38,   -13,    -8,     1,    -5,     5,     0,   -14,   -33,    23,    15,    18,   -25,   -26,     6,     5,   -10,   -28,   -23,   -12,    10,     5,    -5,    -9,    -9,   -22,   -21,   -14,    -5,     2,     2,     0,    -5,     0,     2,    -1,    -1,   -10,    -3,     2,    -8,   -17,   -21,   -22,   -11,   -20,   -22,   -15,    -1,    -5,   -14,   -18,   -14,   -10,    -6,    -1,     1,    -2,    -4,    -3),
		    64 => (   -2,    -2,    -5,    -1,     3,    -3,     3,     3,    -2,    -1,    -4,    -4,    -7,   -10,    -3,    -4,     1,    -5,    -4,    -2,    -1,    -2,    -5,    -1,     0,    -1,     1,     4,    -1,     5,    -3,     4,     1,    -3,   -18,   -14,   -10,    -7,   -20,   -16,    -5,   -18,    -7,   -13,    -9,     1,     3,    -1,    -4,    -3,    -2,    -7,     1,    -2,    -1,    -1,     3,    -1,    -1,     4,    -3,    -1,   -23,   -19,   -24,   -37,   -34,   -40,   -24,   -17,    -7,    -8,    -6,    -6,    -8,    -5,   -17,    -4,    -7,    -9,    -4,     1,    -2,     3,     0,    -3,     3,     2,   -11,   -14,    -5,   -11,   -35,   -51,   -28,    -2,   -12,   -30,   -22,     0,     0,    -6,    23,     8,   -12,    -4,   -16,     1,    12,    -2,     5,     0,    -4,     0,    -5,   -10,   -15,     0,     3,    -5,   -11,   -19,     0,    -7,   -14,   -19,   -14,   -18,   -12,   -16,    -1,    11,   -12,    -9,     7,    31,    12,    11,   -17,    -9,    -1,     4,    -1,    -7,    -6,   -20,    -5,   -19,    10,     0,    15,   -31,   -54,   -70,   -59,   -17,    23,    17,   -29,   -30,   -18,   -21,    -5,    22,     2,    14,   -16,    -5,     4,     3,    -4,   -23,   -18,    -6,    16,     7,    10,    21,   -22,   -54,   -62,   -94,   -67,   -11,     7,    20,    -8,   -43,   -14,     3,    20,    26,   -11,   -27,     7,   -12,    -5,   -23,     0,   -19,   -18,     1,    -3,     0,    21,    32,    11,   -32,   -79,  -108,   -35,    19,    13,    16,   -38,    -5,    12,    24,    52,    15,   -35,   -32,    -8,   -31,   -12,   -19,    -7,   -24,   -21,    -9,    11,     0,     8,    32,    13,   -20,   -94,   -70,   -19,     7,    25,    -3,   -32,   -22,     6,    20,     6,    15,   -40,    -5,   -25,   -25,     2,    -8,    -3,   -27,   -18,    -5,   -18,    15,    23,    22,    16,   -12,   -35,   -27,   -11,     0,    10,    -9,    -9,     0,    -1,     3,     1,    21,   -16,   -10,   -17,   -10,    -3,     4,     1,   -28,    -3,     0,    -5,    11,    16,    34,    23,     3,   -33,   -43,    -7,    18,     6,     1,     2,    -5,   -16,   -15,   -12,    -3,    13,     8,    -9,   -15,     3,    -8,    -5,   -18,     6,    10,     7,     3,    24,    33,    13,   -15,   -30,   -29,   -20,    -8,    -4,     1,   -15,    -8,     3,    -6,     3,   -12,    -5,    12,   -12,   -28,     4,    -8,     5,   -37,   -14,    -4,    13,    -7,     5,    21,    11,    -3,    -4,     5,    -6,     8,    -1,     2,    -3,     7,    18,    -4,     2,   -29,   -25,    -5,   -13,   -27,    -4,    -1,   -10,   -24,   -28,   -19,    14,    10,    -6,    23,    10,     0,     0,    12,     4,    13,    -1,     5,    16,    29,    -6,     5,     5,   -38,   -38,    -1,   -15,     4,    -4,     7,   -29,    -7,     2,   -11,   -13,     8,   -19,   -13,    -1,    -5,     2,    -6,     8,    23,     6,    18,    16,     4,     6,    16,   -14,   -42,   -31,     6,    33,     3,     4,    -2,    20,     3,    24,    -3,    20,    -2,    21,   -14,   -11,   -17,   -21,     1,   -11,    16,     5,     1,    -7,     4,   -29,    -5,     7,    17,   -24,    12,    41,     5,     2,     1,   -15,    14,    -5,   -22,   -18,    12,    -4,     6,    -4,   -11,    -7,    -7,   -19,     7,    -5,    -2,    -2,   -16,   -44,     0,     5,    -3,    29,    36,    12,    -5,     4,    -2,    -7,     2,     2,   -16,   -15,     8,     6,     2,    -9,   -12,   -17,   -12,   -23,     7,     1,    -9,     0,   -23,   -19,    15,    -4,     7,    14,    39,    31,   -10,    -2,    -1,    -7,    -4,    -4,   -22,   -17,     4,    -2,     0,   -19,   -31,   -32,   -10,   -15,    10,   -15,   -11,     7,    -8,   -12,    -4,    -7,     3,   -15,    -7,     2,    -9,     5,    -6,   -13,     6,   -10,   -18,    -6,     9,   -12,   -11,   -16,   -29,   -26,    -1,    -4,    15,    -3,   -13,    22,    -8,   -27,   -10,    -2,   -12,   -15,   -20,     1,   -10,     4,    -1,     0,   -14,   -18,   -18,   -17,    12,    -8,    -9,   -22,   -11,   -31,   -12,    -6,     3,     6,    -4,     3,     8,    -4,     6,    11,     2,    -5,   -32,    -1,     0,     3,     4,   -16,   -19,     0,    -1,    -7,    12,     5,   -10,   -19,   -46,   -28,    -5,    20,     5,    -5,    -6,    -1,     6,     2,     0,    -9,    18,    -1,   -35,   -17,    -2,     3,     2,     2,   -12,   -18,     2,     5,    -3,     9,   -17,   -28,   -32,   -21,    -5,     5,     5,   -11,   -24,    -5,    23,     2,     7,    11,    28,   -14,   -14,    10,    -1,    -3,     3,    -4,    -5,   -11,   -14,     2,    -2,   -10,    -3,   -11,   -37,    -6,     9,     7,    -3,   -12,   -25,    11,    17,   -13,    25,     2,   -12,   -29,    10,     3,    -1,    -1,    -2,    -2,     1,   -14,   -12,   -11,   -18,     4,    -4,   -12,   -15,   -11,    -5,    10,    14,     0,     0,     8,     5,     6,     9,    20,   -14,   -34,     3,    -9,     5,    -2,     4,    -2,     0,    -6,    -3,   -12,    -8,     9,    -6,   -18,   -17,    -1,    13,   -27,   -15,   -14,    10,    10,     5,    20,    12,   -11,   -12,   -15,    -8,    -7,     3,     4,    -5,    -3,   -10,    -5,   -10,    -4,    -1,     5,     2,   -14,    -9,    -8,   -56,   -62,   -58,   -30,    -4,   -13,   -34,   -44,   -40,   -50,    -2,   -14,     0,    -4,    -1,     3,     3,    -1,    -2,     3,     1,    -8,   -18,   -20,   -12,    -9,   -20,   -20,   -18,   -20,    -7,   -21,   -33,   -25,   -20,   -23,   -26,   -27,    -1,     2,    -1,    -1,     5),
		    65 => (   -4,     4,     2,    -1,    -4,     0,    -1,     3,    -5,    -5,     2,    -2,    -3,    -1,     1,     2,     2,    -2,    -5,    -4,     3,    -5,    -4,     3,    -4,    -3,    -4,    -3,    -1,    -1,    -4,    -2,     1,    -1,    -3,     4,     4,    -1,    -7,    -2,    -5,    -6,    -8,    -9,   -10,    -8,   -10,    -1,    -4,    -2,     3,     3,     1,    -4,    -1,    -5,     0,     2,    -5,     4,    -5,     0,     1,    -3,    -8,    -2,    -5,   -23,   -22,   -25,   -31,   -15,   -19,    19,     1,    10,    24,    -7,    -2,    -7,   -10,    -6,    -4,     0,     1,    -4,    -1,    -1,     4,    -4,   -10,    -8,   -13,   -19,     4,    -8,   -18,    -7,    -6,     7,   -17,    17,    13,    13,    31,    33,    21,   -23,   -18,     9,    32,     3,    -1,     4,   -11,    -7,    -7,   -11,   -28,   -13,   -25,    20,    19,    -1,     3,   -28,   -16,    -8,   -31,    -8,    17,   -14,   -14,     8,    -1,   -11,    -4,    24,    19,   -18,    -3,     4,   -17,   -12,   -10,   -16,   -52,   -55,   -13,    21,     5,    -2,    11,    25,    -5,   -53,   -20,   -15,   -21,   -11,    22,    13,    13,   -13,   -13,    15,    24,    -8,    -4,    -5,    21,   -11,   -18,   -39,   -51,   -54,   -28,    -6,    15,    -7,    27,    26,    -3,   -16,   -18,     0,    -4,     8,    25,    10,    21,    -2,     1,    44,    45,    15,     5,    -5,    20,   -24,   -13,   -13,   -45,   -44,   -25,    15,     2,    -2,    21,    18,   -15,    14,    23,    24,    26,    28,    32,     7,    20,    -2,   -12,    19,    45,     1,    -2,   -10,   -20,   -19,   -11,   -48,   -40,   -20,    -4,    -6,   -14,   -11,    -2,   -13,     2,    14,    21,    26,    45,    35,    26,    -5,     7,    17,    -2,    -5,    24,    14,     2,    -1,   -32,   -34,   -32,   -30,   -19,   -17,   -25,     0,    -7,    -9,   -16,   -11,   -25,   -25,   -13,    26,    11,    -4,   -20,   -16,    -2,    -8,   -12,    19,     4,    23,     4,    -6,    -3,    -6,     5,   -18,    -7,   -35,   -14,    11,   -15,     0,     2,   -15,   -33,   -75,   -78,   -61,   -48,   -67,   -58,   -21,   -27,   -60,   -27,     2,    26,    29,    -3,    -2,     1,    -6,    34,     1,   -35,   -22,   -13,     1,     1,   -11,     1,   -11,   -18,   -48,   -62,   -86,   -79,   -73,   -81,   -50,   -40,   -50,   -32,   -17,     4,    26,     2,    -3,     1,     9,    17,   -15,   -30,   -12,   -10,    -6,    10,     3,    -1,    25,     4,    -3,   -13,   -33,   -22,   -33,   -39,   -54,   -53,   -41,   -32,   -14,    -3,   -13,    -1,    -5,     1,    15,     8,   -11,    -5,     2,   -12,   -18,    -7,   -10,    -5,    12,    15,    12,   -12,   -13,   -16,   -19,    -5,   -42,   -69,   -42,   -34,   -11,    -2,   -14,     1,    -8,    -6,    22,     7,   -18,    -8,    10,     4,     7,     0,     6,     8,    -3,    -9,     5,   -12,    -7,   -13,    -2,    20,    -6,   -15,   -12,   -13,    -8,    -3,    -4,     7,    -7,   -24,   -15,     9,     1,    16,   -16,    -9,    16,    -3,     1,     6,   -12,    -4,    -8,     8,   -10,    -1,   -12,    10,    25,   -11,    -7,    10,     2,    -7,   -15,     2,    -5,   -15,   -14,    -7,    -3,   -17,   -27,    -1,     3,    10,    13,     4,    13,     1,   -16,    -1,     5,   -25,     4,    -4,   -11,   -26,   -32,    -1,   -15,   -25,   -17,     0,    -5,   -20,     0,     3,   -20,   -24,    -9,   -19,    -6,    18,    16,     8,    19,   -11,    -8,    -7,    -6,    -9,     3,    11,   -14,   -20,   -39,    -6,   -18,    -5,   -22,     1,    -5,   -17,     7,     7,    -2,   -32,   -46,   -31,   -40,   -20,    14,    -6,    -5,   -26,   -22,    16,     7,     5,     0,    21,   -18,   -14,    -1,     6,    -4,   -21,   -13,     4,     0,   -13,   -21,    33,    -1,     0,   -22,   -24,   -55,   -50,   -57,   -20,     4,   -15,   -31,     0,    15,     5,    -6,    19,   -18,   -16,    14,    15,   -11,    -3,    -6,     1,    -6,   -10,   -11,     6,    16,     6,     4,    -8,   -30,    -4,   -22,   -39,    -5,    -6,     6,   -13,     4,     5,    15,    13,    -7,    -3,     9,    -3,    -5,   -10,     4,     1,    -4,   -24,    -2,    24,    14,     3,     3,    -1,     8,    11,    -2,    -3,    12,     5,     3,   -11,   -11,     5,    21,     4,   -13,    14,    10,    -9,    -5,   -16,     1,     4,     3,   -27,    25,    11,   -15,    -7,   -12,     8,    31,    24,    20,     5,   -15,     9,   -10,    -6,     8,    -3,    -1,     5,    -1,    -2,    30,    -2,    -8,    -4,    -4,    -1,     3,    11,    32,    28,    14,    20,     3,     5,   -19,     7,    16,     7,     2,    -4,     3,   -16,    -8,    -5,     4,     5,     0,     8,    32,    -6,   -20,     3,    -4,     5,     4,   -17,     6,    -9,    -9,    -2,     1,    -7,     2,     4,    -9,    -6,    -3,     2,     1,   -15,   -10,    12,    -7,   -17,     7,    41,    10,    16,   -23,   -13,    -2,    -4,    -5,    -4,    36,   -28,   -28,   -11,   -17,   -26,     3,   -15,   -12,     4,    21,    -7,    -6,   -44,     8,     9,     5,    13,    34,    51,    25,    15,     0,     1,     0,     0,     3,     0,    -3,    -4,    -9,    -8,    -9,   -14,   -25,    -6,    18,    22,    11,   -42,   -49,   -41,   -43,   -20,    10,   -16,    14,    12,    -5,    -4,     0,    -2,    -3,     5,     0,    -2,     1,     0,    -5,     1,    -3,    -5,    -8,    -1,     2,     5,     8,   -11,    -1,    -1,    -1,    -7,    -3,     2,    -6,   -12,    -5,    -3,    -2,     5,     1),
		    66 => (    0,     2,     1,    -3,     4,     4,    -1,    -2,     3,    -5,    -1,     1,    17,    20,     3,    -4,    -1,     0,    -4,    -3,    -1,     4,     2,     4,     4,    -3,     1,     0,    -1,     4,    -3,    -4,     1,     1,     9,     9,     4,     2,    22,     3,     9,    24,   -11,   -10,    -5,     5,    13,    21,    23,    19,    17,    15,    -1,     5,    -1,     0,    -1,    -4,     1,    -6,     7,    15,    10,    -2,     5,    19,    17,    17,    11,    17,    14,    -7,    15,    15,    21,    33,    28,    16,    47,    32,    24,    19,     1,     1,     4,     3,   -28,    15,    -3,    28,    31,    29,    40,    41,    47,    47,    61,    39,    53,    37,    10,     4,     5,     4,   -15,   -20,   -14,    -1,    19,   -39,   -33,     1,     3,    -4,   -21,     2,    16,    25,    27,    39,    19,    41,    36,    19,    35,     6,    41,    34,     9,    15,     7,    21,    26,    14,    -7,   -10,   -12,   -26,   -10,    30,    -5,    -2,   -11,   -23,    35,    16,    21,    25,    16,    18,    32,     7,   -18,    16,    34,    17,     5,    25,     3,   -10,     6,   -22,    -4,     2,    28,    13,    26,    10,     2,     0,     0,     2,    27,    10,    29,    16,    -4,    12,    -7,   -16,    10,     8,     8,     3,     2,     1,   -32,     7,    -3,   -19,   -19,   -17,    -4,    11,    25,    35,     2,    -4,    -2,   -10,    27,    19,    10,    10,     2,    -9,   -15,    -7,   -23,   -30,    11,   -11,    -4,   -10,   -10,     3,   -10,    -6,    -7,    -6,    10,     3,    22,    23,    -3,   -11,   -14,   -53,    31,    10,     6,   -12,     1,    16,   -14,   -15,    -9,   -18,     1,   -24,   -43,   -18,   -11,    -4,    10,    11,   -10,   -19,   -19,   -42,    -3,   -33,     0,    -4,   -18,   -29,    24,    -6,   -17,   -12,     4,   -10,   -15,   -18,   -27,   -32,     0,     2,   -17,   -41,    -7,    -8,    -4,    20,    -4,    -5,   -29,   -52,   -32,   -28,    -3,    -4,   -20,   -16,     7,     3,   -18,   -19,    -4,   -11,    -7,   -26,   -33,   -15,     4,   -13,   -36,   -22,   -30,   -22,     4,     2,   -24,   -21,   -35,   -38,   -32,   -31,    -1,    -5,    -4,   -32,     7,     4,    -2,    -5,   -16,    -6,   -13,   -25,     3,    -3,    -5,   -22,   -18,   -16,   -19,   -10,   -10,     2,   -21,    -5,   -16,   -32,   -35,   -24,     5,    -4,   -15,   -30,    -5,     8,    22,     7,    -8,     8,    -2,     4,    -8,    12,   -17,   -11,   -27,   -17,   -24,   -18,    13,    10,   -15,    14,    21,    -2,   -47,   -24,    -2,     3,   -11,   -26,   -12,    10,    -3,   -12,   -12,    21,    26,    17,    17,     9,    12,     4,    -6,   -31,    -9,    13,    14,    16,   -10,    16,    11,   -15,   -49,    -1,     0,    -2,    -5,   -26,   -36,    12,   -15,   -25,     8,     9,    26,    26,    27,    14,     6,   -18,    -4,   -18,     8,     9,     5,    12,    12,   -14,    -7,    26,   -39,    -8,     0,    -2,   -15,   -17,   -40,   -14,   -13,    -5,   -12,    -4,     7,    13,     0,    31,    20,   -13,   -14,   -33,     2,    17,    -2,     5,   -24,     3,     0,    22,   -17,   -47,     3,    -1,   -23,   -18,    -9,     8,     7,    11,   -11,    14,    13,     5,    -9,   -17,   -11,   -10,   -12,   -15,    22,    24,   -10,    -8,     7,    -1,    -7,    17,   -25,   -38,    -5,     1,   -27,   -27,   -18,    23,     1,     9,    -5,   -18,   -10,    -5,    -9,   -16,     3,    10,    10,    17,    13,    16,    13,    -6,    -5,   -11,    -6,    15,   -24,   -54,     4,    -3,   -26,   -42,    -8,    -3,   -18,     4,    -2,     5,    17,   -28,    -2,    -4,     0,   -20,     2,    16,    42,    34,     3,   -13,     1,     7,     5,    26,     2,   -23,     3,     0,   -31,   -34,     4,    12,    11,    -4,     2,     2,    31,    32,    18,     8,     5,     9,     1,    23,    -1,    34,    -3,    -2,    -6,   -13,   -27,     8,   -16,    -1,     1,    -2,   -28,   -42,    -2,    -2,     1,    13,     5,     8,    27,    29,    24,   -16,     7,     7,     6,    16,    18,    15,    16,    -2,    -3,   -31,   -37,   -10,   -10,    -1,    -3,    -5,   -36,   -38,   -29,   -34,   -10,    23,    28,     0,    14,     1,    42,    19,     8,     5,    34,    21,    18,    11,     7,   -11,    -7,   -33,   -17,    -2,    -3,    -5,     1,     3,   -26,   -30,   -54,   -67,   -89,     0,     1,    17,     9,     5,     2,     0,     3,    23,    27,    38,    24,     3,     8,     7,   -27,   -24,   -59,   -16,    -6,    -4,    -1,     4,     4,   -33,   -41,   -46,   -43,    -6,   -11,     2,   -18,     5,    20,    -5,    10,    22,     2,   -18,     5,     1,     3,    14,   -33,   -41,   -39,   -27,   -32,     5,    -4,     2,    -3,    -5,   -13,   -15,   -23,   -43,   -59,   -77,   -53,   -68,   -33,   -33,   -21,     6,    11,    16,    34,   -52,    -8,   -28,   -24,   -22,   -17,   -11,    -5,     0,     3,     3,    -2,    -2,    -4,   -10,   -17,   -17,   -12,   -16,   -19,     7,    15,    -9,    -8,   -14,   -24,   -24,   -13,   -39,   -36,    -7,   -19,   -19,   -15,     4,    -2,     4,     2,     4,     0,    -1,    -4,    -7,     3,    -6,    -2,    -6,    -4,    -9,    -3,     1,    -2,    -8,    -1,    -5,     0,    -6,    -5,     5,    -4,    -5,     3,     3,     2,     4,     0,     2,    -3,     5,     2,     2,     0,    -1,     5,    -2,    -3,    -4,     2,     2,    -3,     0,    -2,    -4,     1,     1,    -5,    -6,    -3,     2,    -4,    -1,     2,     1),
		    67 => (   -4,    -4,     3,    -3,     1,     2,     2,     3,    -5,    -4,     4,     2,     4,     1,    -1,     0,     5,     3,     3,     4,    -2,    -4,     3,     4,     2,     4,    -4,    -5,     3,    -3,    -1,     0,     2,    -2,     4,    -2,     3,     2,    -2,    -5,    -5,    -7,    -8,   -19,   -19,   -12,    -1,     1,     1,    -3,    -2,    -3,     3,     3,     1,     3,    -3,    -3,     5,    -3,     0,    -2,    -5,    -2,    -8,     6,    -4,   -18,   -28,   -12,   -13,   -12,     4,    -1,    -4,    -5,    -6,    -6,    -2,     5,     1,    -1,     1,    -3,    -4,     3,    -3,     0,    -7,   -15,   -17,   -28,   -12,    -5,   -12,   -19,   -34,   -35,   -25,   -24,   -16,   -12,    -5,     1,    -4,     4,   -10,    -3,    -8,    -7,     4,     0,     4,     0,     0,    -3,   -13,    -3,   -21,   -21,   -30,   -37,   -53,     2,     5,     2,    -8,   -25,   -59,   -44,   -33,   -34,   -26,     3,   -17,   -21,   -23,   -14,    -6,    -4,    -3,    -4,    -1,   -13,   -19,    -8,   -39,     2,    39,     8,    -8,     0,    12,    -5,    14,     4,     6,    -1,    30,    -2,   -20,   -10,    -8,   -18,   -31,    -5,    -7,    -2,    -2,     1,    14,   -10,   -10,    -8,   -25,    11,    17,    27,    13,    -4,    -7,    -7,    -9,    12,     6,     1,    19,     7,   -37,   -17,     2,   -20,   -20,   -14,   -15,    -8,     4,    11,    16,     0,     9,     0,    11,    10,    14,    11,    -3,   -10,   -20,   -21,   -23,    -2,    19,    20,    15,    24,    36,     6,   -15,   -16,   -27,   -15,   -14,    -8,   -20,     6,    38,     2,    16,    11,     6,    25,    23,     2,    -4,    -9,    -6,   -17,     2,    23,     6,     5,    10,    12,    24,    13,    -3,   -35,   -23,    -5,   -10,    -7,     7,     8,     9,    19,    18,   -27,    -7,     1,     8,    -2,     7,   -15,    -9,     7,     1,    -6,     7,    21,    -6,    -5,    11,   -18,   -10,   -22,   -14,    -3,   -19,     7,     6,     3,    -6,     5,    26,    -7,    -6,     4,   -11,     9,     6,   -17,   -33,     6,    -3,     4,     4,    -5,     1,     5,    -6,   -24,    -6,   -18,   -18,    -3,   -14,     1,     7,     7,    -4,   -20,     0,     4,   -10,    15,     7,   -10,     4,     0,   -33,   -22,     0,    29,    -3,    -1,     0,    -2,   -20,   -14,   -19,   -39,   -21,   -23,   -18,     7,     3,     3,   -16,    -5,   -15,    -4,   -16,    14,    -3,   -22,   -12,   -37,   -38,   -26,   -15,    19,    -9,   -26,    -8,   -34,   -20,   -20,   -37,   -36,   -40,   -10,   -12,     3,    -2,    13,    15,    -6,    -5,    -4,   -13,    -1,     2,   -15,   -21,   -35,   -69,   -45,   -24,    -5,   -13,    -1,   -10,   -32,   -28,   -28,   -33,   -44,   -39,    -5,   -23,   -11,    -1,    16,     5,    17,    -2,    12,   -27,   -14,   -26,   -41,   -72,   -57,   -37,   -27,   -21,     1,   -20,     7,    16,     4,   -11,     8,   -24,   -29,   -11,    -6,   -19,    -7,     4,    -2,    -1,    13,    10,    -6,   -19,   -50,   -31,   -28,   -40,     4,    -7,    -5,   -24,    -1,    -2,    18,    21,     5,    13,    12,    -6,     3,     4,    10,    -6,    -9,     2,     2,     1,   -13,    -8,     0,   -32,   -16,    28,   -10,    -9,    25,     8,    -1,    -5,    21,     9,     4,    19,   -12,    -4,   -20,   -13,    -6,    -5,   -31,   -15,    -4,     4,     0,   -15,   -12,   -19,   -35,   -17,   -13,    -7,     1,   -22,     2,    -6,     2,    -7,     8,     6,    18,    11,     1,   -35,   -37,   -30,   -25,   -10,   -48,   -27,   -33,     6,     2,     7,   -18,   -16,    -5,   -13,     2,   -11,     6,    -2,     3,   -21,    15,     6,    26,    -2,    28,   -15,    10,    16,     3,   -24,   -31,   -19,   -37,     3,   -23,    -2,     2,     1,    -2,    -5,   -33,   -13,   -12,    11,    -9,    -9,   -24,   -11,   -11,    24,    35,   -15,   -14,   -12,    10,    17,    18,   -11,    -4,     7,   -15,   -20,   -17,    -1,    14,    -7,    -1,    -6,   -27,   -21,    -1,     7,    10,    -5,   -50,   -15,    -7,    10,     8,   -14,   -26,   -11,    -4,    15,    -2,   -12,   -41,   -22,   -12,   -21,     3,    -6,     3,    -6,   -10,    -8,   -28,   -39,   -35,     8,   -10,   -17,   -27,    -6,     1,    14,     5,    21,   -28,   -12,   -18,   -11,     4,   -14,   -49,   -27,   -26,    -2,    -1,    -7,     2,    -4,    -3,    -6,   -23,   -32,   -31,   -18,   -24,   -13,   -26,   -16,    18,     4,    15,     4,     8,   -19,   -10,   -14,   -41,   -62,   -45,   -26,   -15,   -25,     2,    -1,     5,    -7,   -17,   -35,   -36,   -32,   -48,   -41,   -56,   -38,   -33,   -19,    -9,    -9,     1,    -6,   -30,   -44,   -31,   -28,   -30,   -28,   -22,     7,   -15,   -23,    -4,    -5,    -4,     3,     0,   -14,   -35,   -42,   -41,   -61,   -57,   -42,   -28,    -7,     0,     7,    22,    -4,    -7,   -40,   -25,    -3,   -11,    -3,   -19,   -12,   -13,    -3,    -1,    -3,     0,   -23,     0,     3,   -15,   -23,   -33,   -33,   -52,   -31,     9,   -14,   -12,    -4,    27,     3,     7,    -2,    14,    19,    13,    -8,   -15,     0,    -2,    -4,    -2,     1,    -3,     0,    -1,   -12,   -12,    -4,    15,     9,     9,   -13,    -9,    13,    20,    10,     4,    -1,     7,    56,    46,    28,     8,    -5,    -8,    -2,     0,     0,     0,    -3,    -2,    -1,     2,    10,     2,    -2,    -9,     1,    20,    28,    17,    13,    12,     5,    22,    20,    34,    50,    32,    15,    -2,   -10,     4,     1,    -4,    -3,    -5),
		    68 => (    3,     5,     4,     1,    -2,    -4,     2,    -5,     1,    -3,    -5,    -1,    -2,     2,     1,     3,     3,     2,    -1,     1,     1,     1,    -2,    -1,     0,    -5,     5,     2,     4,    -2,    -2,    -3,     4,     3,     4,    -4,     2,     0,     4,    -2,     1,     0,    -1,    -4,   -21,   -18,     1,     0,    -2,    -5,    -4,     2,     1,    -1,     3,    -2,    -1,    -5,    -4,    -3,    -5,     1,     2,    -4,     5,    -6,   -11,    -3,     0,    -4,     2,    -2,   -11,    -1,     0,     0,    -4,   -11,    -5,   -10,    -2,    -4,     4,     4,    -4,    -2,     0,    -2,    -4,    -9,    -5,   -11,    -8,    -7,     0,     0,    -4,     1,   -17,   -12,    -4,    -2,     6,    -4,   -10,     2,     5,     4,    -4,     1,    -8,     3,     4,    -3,     2,    -8,    -5,    -5,   -15,   -15,     4,     1,    -3,    15,    15,   -10,    -1,   -26,   -21,    -5,     8,     2,     6,    -9,   -10,    -1,    -7,     2,     1,     0,    -4,    -5,     0,    -9,   -23,   -28,    -1,    -4,     1,     1,   -12,    -6,   -12,   -11,     3,    -6,   -17,    -7,    -9,   -11,    -3,    -8,   -13,    -7,    -4,    10,     0,    -8,    -4,     1,   -10,   -20,    -4,     4,    -4,    11,    -3,   -10,   -16,   -24,    -9,   -23,   -13,    -1,    -2,     2,    -6,    -8,    -6,   -14,    -6,    -4,    -4,    -7,    -5,     0,     2,    -2,    -8,     0,     5,    23,     4,     6,     3,    -5,    -6,   -14,     3,     2,     6,     9,     7,     4,     2,     5,   -15,    -5,     4,     1,     7,    -1,     2,    -5,    -2,   -11,    -4,    19,    29,    32,    12,    -4,   -18,   -13,    -4,     7,     3,     5,    -2,   -12,   -16,    -9,    -9,    -9,     2,     4,     5,    -6,    -5,     3,    -9,    -2,     1,   -13,   -17,    15,    25,    29,    11,   -10,   -26,   -16,    10,   -16,   -16,    -9,   -13,   -24,   -21,    -5,   -10,    11,    12,    13,     4,    -1,     1,    14,    -7,    -6,    -3,    -9,   -17,     9,     7,    23,    19,    12,   -13,     3,    11,    -3,     0,    -9,    -9,   -13,   -11,     0,    -8,     1,     5,    -2,   -10,   -10,    -1,   -14,    -7,    -8,     0,    -2,   -22,   -12,   -10,    -2,    19,    24,    16,    23,    17,     5,    -5,    -9,   -13,    -7,    -7,    -9,   -19,    -2,    -6,    -5,     4,    -5,   -11,    -7,    -1,   -18,     1,     2,   -13,   -28,   -22,    -5,     2,   -10,     9,     4,    16,     2,     0,   -20,   -21,     0,     0,    -4,    -4,   -14,   -13,    10,     4,    -5,    -8,   -13,   -14,   -22,     1,    -6,   -20,   -31,   -12,   -19,   -19,   -20,   -19,   -17,    -9,     3,     2,   -12,     5,     6,     2,   -13,   -12,   -22,   -18,    -3,    -3,    -5,   -13,   -22,   -13,     7,    -8,    -5,     4,   -31,   -13,   -12,   -17,   -25,   -23,   -34,   -17,   -24,   -14,    -1,    -5,   -18,   -19,    -2,     1,    -8,   -19,    -7,    -3,    -4,   -16,    -7,   -35,    -4,     1,     5,    -6,     6,     1,    -7,   -12,   -22,   -14,   -20,   -15,    -8,   -11,    -1,    -2,    -6,    -2,    -6,    -2,   -12,    -1,   -14,   -11,   -12,   -14,     7,   -12,   -15,     3,    -7,    -2,     8,    -1,    -7,   -16,    -9,    -4,   -18,     0,     4,     0,   -10,   -20,   -22,     8,     9,   -10,    -7,    -3,     0,     0,   -10,    -9,     4,   -16,   -12,     5,     0,     0,    13,    -4,   -12,   -10,    -8,   -13,   -13,    13,    15,    -2,   -15,   -15,   -24,   -13,     7,     1,   -11,    -8,     5,    10,   -14,    -6,    -8,    -4,    -7,    -1,    -4,    -3,     2,   -10,    -8,   -11,    -8,   -14,   -12,     5,     1,     6,     1,   -20,   -16,   -16,    12,     4,    -5,   -18,    -8,    16,    -4,    -8,     3,    -1,   -14,     2,     2,    -6,    -2,   -11,    -5,    -4,    -7,   -28,    -1,    11,    12,    -2,     2,   -14,   -17,   -17,    -3,    14,     5,    -5,     2,     9,    10,     0,     2,   -10,   -11,    -4,    -1,   -10,    -8,    -9,    -6,    -3,    -9,   -18,    -3,     6,    15,     7,   -18,   -22,   -15,   -21,    -4,     7,     2,     0,    -1,    15,     4,    -5,    -1,   -13,     1,    -7,    -8,    -3,   -14,    -4,    -5,   -18,   -13,   -11,    -8,    -6,     5,     7,    -4,   -11,   -10,   -20,     3,     7,     3,     2,     4,    16,     0,    -6,    -7,    -6,    -1,   -16,    -6,    -6,   -10,    -6,   -12,   -10,    -7,   -11,   -14,    -3,    -3,    -6,    -4,   -10,    -7,   -12,     6,    -3,    -2,     0,    11,     5,    -5,   -17,    -6,    -2,     1,     4,     4,    -1,    -8,    -8,   -15,   -15,   -11,    -5,   -11,    -2,   -17,    -7,     9,    -7,     0,     7,     1,    -5,     1,     8,    15,     6,    -9,    -1,     0,   -22,     0,    -3,     5,    -6,     1,    -4,   -10,    -9,     4,    -8,    -2,     0,   -15,   -14,   -15,     5,    11,    13,   -12,   -20,   -13,    -1,   -13,   -15,    -5,    -5,    -7,    -3,     4,     2,    -3,    -8,    -7,    -8,    -9,   -11,   -13,    -9,     1,    12,    -9,   -11,    -8,     0,     5,     1,    -3,   -10,    -8,   -15,   -12,     0,    -2,    -6,    -3,    -9,    -4,     0,    -2,    -1,    -2,     0,    -8,    -6,   -13,    -7,   -15,   -13,   -12,   -14,   -10,   -19,   -16,    -5,    -1,     0,   -20,   -24,    -2,   -16,     0,     2,     3,     0,     1,    -1,     5,     4,     1,    -2,     2,    -1,    -3,    -2,    -8,    -7,    -3,     1,    -7,    -5,    -3,    -8,    -6,   -14,    -3,    -2,    -2,    -4,    -4,    -1,     4,    -4,     1),
		    69 => (   -3,    -4,     3,     4,     4,     4,     0,     5,    -5,     3,     5,     4,    -1,     2,     1,     2,    -4,    -3,     5,    -3,     1,    -2,     2,    -1,     1,    -4,     0,     1,     1,     3,     5,    -4,     1,     0,    -3,    -9,   -11,    -9,    -8,   -13,   -15,   -23,   -12,   -27,   -23,   -24,   -12,     1,     3,    -4,   -12,     1,     4,    -4,    -4,    -3,    -4,    -2,    -4,   -18,   -21,    -4,    -4,   -21,   -27,   -12,   -13,   -20,     2,     0,   -57,   -32,   -29,   -18,   -32,   -23,   -43,   -48,   -35,   -29,   -18,    -9,     4,     1,     1,    -1,    -2,   -24,   -31,   -27,   -17,   -29,   -64,   -80,  -107,   -96,   -64,   -83,   -77,   -83,  -109,   -94,   -30,   -41,   -67,   -58,   -48,   -28,   -24,   -15,     5,     3,     4,    -3,   -13,   -21,   -35,   -44,   -63,   -44,   -49,   -54,   -33,    -9,     4,    -5,   -17,   -17,   -15,   -31,   -57,  -113,   -72,   -59,   -59,   -31,   -26,   -43,   -31,     2,    -2,     1,   -13,   -20,   -16,   -26,   -27,   -18,   -39,     7,     7,     2,    14,    31,    10,    12,    26,    26,    -4,   -16,   -33,   -14,   -66,   -28,   -41,   -42,   -29,    -7,    -2,     4,   -13,   -43,   -32,   -39,   -21,   -13,    -1,    20,    21,   -10,    -8,    30,    13,    31,    49,    30,     7,    11,    -7,    -4,    -8,     7,     1,   -14,   -32,   -38,     1,   -15,   -28,   -36,   -23,   -42,    -6,    -4,    -7,     8,     7,    -5,    18,    36,    34,    29,    59,    35,     0,    11,    18,    -2,    10,     9,     0,     3,   -35,   -29,   -25,   -33,   -25,   -28,   -31,    -3,    12,    -6,     0,    10,     3,     2,    24,    21,    32,    49,    39,    27,    24,    29,     2,    12,     8,    19,    20,     1,   -33,   -18,    -5,   -23,   -33,   -35,    21,     8,    20,    10,    11,    22,     4,    -6,    10,    28,    26,    16,    12,    10,     8,     7,    23,     0,    -2,    -9,   -11,   -36,   -43,   -29,    -2,   -16,   -47,   -22,    21,    22,     1,     4,    -3,    -3,     1,    -2,    16,    11,     6,   -20,     1,   -12,     0,    -1,     6,   -22,   -13,   -11,   -28,    18,   -46,   -18,    -2,   -73,    -1,   -16,     6,    25,    10,    -9,   -22,    -6,    -6,   -17,     0,   -28,   -23,   -25,    -1,     7,   -19,    -9,    16,   -10,   -31,   -20,   -27,    -3,   -38,   -15,     1,    -8,    -5,   -15,    17,    10,     8,   -10,   -24,   -25,    -9,     0,   -21,   -27,   -13,   -21,   -11,     6,   -15,   -23,     5,   -17,   -15,    -3,   -32,   -53,   -32,   -22,    -5,   -15,   -23,   -16,     8,    -8,     6,     4,     1,   -15,    -4,   -15,     1,    -8,   -13,   -24,     6,     0,    -7,   -12,   -16,     1,   -19,   -18,   -14,   -39,   -24,    -7,    -9,   -14,   -14,    -3,    11,    -6,    -3,     7,     1,    -2,     2,    -9,    13,   -23,   -15,     9,     2,     0,    10,     8,    -2,   -15,   -22,   -44,   -20,   -46,   -28,     0,     0,    -2,   -33,   -14,     6,     4,    12,     3,    17,    11,   -17,   -23,   -20,    -6,    12,     9,    18,    10,    16,    25,    30,    11,     5,   -33,   -18,   -44,   -10,   -29,     3,    -8,   -23,   -15,     0,    18,    18,    -5,     8,     2,    -6,   -27,   -27,    -8,    22,    15,     3,    20,    -7,    15,    24,     5,    -1,   -23,    -8,   -56,   -30,   -33,    -1,    -1,   -33,     3,   -20,     6,   -17,    -8,    -1,     7,    -9,   -17,    -5,   -11,    15,     5,     4,     8,   -13,     1,     7,   -11,   -45,   -53,   -16,   -68,   -40,   -23,    12,     1,   -39,    29,   -18,   -17,    -4,     0,   -29,   -14,   -17,   -23,   -35,    -5,   -15,    -9,    13,     7,   -30,     6,     2,   -23,   -15,   -17,   -23,   -53,   -34,   -15,     3,    -8,   -33,    14,    -4,   -17,   -24,    -9,   -31,   -12,     0,    -9,    -6,   -17,    -1,   -18,    10,   -10,    -6,     4,    -3,   -20,     0,    18,   -11,   -35,   -26,   -10,     2,   -10,   -63,     5,   -23,     7,    -2,   -41,   -11,   -20,   -11,   -13,   -26,   -18,   -13,   -19,     4,     4,   -12,     4,   -17,   -26,     1,    35,    31,    15,   -19,     1,     4,    -3,   -53,     7,    -9,    10,     9,   -10,   -14,   -27,     7,    -5,   -19,   -13,    -3,   -10,    21,    18,    -4,   -18,   -29,    -4,     8,    26,    23,    -4,   -51,     2,     2,     0,   -41,    15,   -15,    -2,   -11,   -17,    -1,   -13,     0,   -22,     8,   -11,    19,     4,    24,    22,     2,   -18,    -9,     4,    31,    31,    25,   -37,   -37,    -2,     0,     3,    -6,     8,   -14,     3,     5,    30,    13,     1,   -11,    -4,     2,    11,    25,    21,    16,    11,     9,    -1,    -8,    -4,    12,    25,    38,   -17,   -26,     3,    -5,    -1,   -19,   -27,   -10,    12,    35,    44,    27,    19,     7,    15,     6,    11,   -23,   -14,   -17,    11,    44,    21,    23,     4,   -18,     5,     8,   -17,    -2,    -2,    -2,     1,    19,   -23,    -4,    17,    30,    40,    27,    25,     1,    10,    -6,   -17,    13,    -7,    -4,    29,    23,    11,    20,    -9,    -4,   -15,     0,     1,    -7,     2,    -1,    -4,     1,    18,     1,    10,    20,    36,    -8,    10,    -1,   -14,    11,   -10,    27,    25,    11,     1,    12,    -5,    36,     8,   -12,    23,     9,    -1,     4,     0,     3,     2,    -2,     3,    -1,   -18,     7,     5,     7,    -1,     9,    14,    17,    10,    14,     5,    14,   -21,     0,     7,   -12,   -29,   -21,   -19,     2,    -2,     5,    -4),
		    70 => (    1,    -3,    -2,     2,     5,    -2,    -3,     1,    -1,     4,     0,    -3,     0,     0,    -4,    -3,     3,    -5,     1,     1,    -4,     4,     0,    -2,     5,    -1,    -2,    -1,     3,     5,     5,     0,     0,     0,     0,    -1,     3,    -5,    -3,     0,     4,    10,    -6,     2,    -4,     2,     3,     0,     1,    -1,     4,     5,     0,     1,     1,     1,    -1,     0,     2,    -3,    -3,    -4,    -6,     2,    -8,    -8,    -1,    -9,   -12,   -20,    -8,     4,   -10,   -14,    -6,    -4,     0,    -5,    -1,    -5,    -3,     3,    -5,    -2,    -5,     5,    -5,    -4,    -2,     7,    -9,   -10,   -11,   -39,   -21,   -13,     2,    14,     7,   -21,    -4,    -3,     1,     2,    -9,   -21,   -21,   -10,     4,     2,    -2,    -4,     3,     4,     5,     2,    -8,   -34,   -11,    -2,   -12,    -5,    -7,    21,    28,    32,    15,     9,   -26,   -32,    -8,     5,   -25,   -28,   -14,    -9,    -9,   -17,    -9,     0,    -3,    -2,   -10,    -4,    -7,   -22,    -8,     2,     3,    -1,     4,    10,    34,     9,     9,    16,    -6,   -30,   -22,    15,   -15,   -30,     2,     6,    -2,   -24,   -20,   -12,     5,    -6,    -3,    -7,     6,     9,    12,    11,    13,     4,     0,    29,     4,    -4,     4,     1,    20,    13,   -15,     0,   -11,    -7,    -4,    -7,    -5,   -35,   -18,    -7,     0,    -3,    -8,   -19,     4,    13,    18,    15,     5,    13,     3,    15,    -3,     4,    23,    13,    26,     8,     7,    10,    14,     9,   -18,    -7,    -7,    -7,   -20,   -15,     4,    -4,    18,   -15,    14,     1,    10,   -12,    -2,    19,    15,    -5,   -12,    19,    15,    -5,   -14,   -15,    18,     1,     7,    18,    -4,     1,   -16,   -11,   -30,   -12,     4,    -1,    25,    -4,    -5,   -11,   -20,   -18,    14,    17,    21,    -3,    -7,    18,    -3,     2,   -10,    -3,    -9,    22,    -4,   -11,    -8,   -11,   -20,   -20,   -24,     4,    -1,     4,    24,     6,   -14,    -3,   -16,   -19,    12,    11,    -3,    -1,     1,   -21,    -6,    13,     2,   -11,   -19,   -17,   -22,   -12,   -12,    12,    -5,    -9,   -19,     2,     2,    26,     1,   -13,   -17,    -4,    -8,   -12,    -3,    -5,    11,   -12,   -38,   -57,   -43,    -7,   -13,   -20,   -20,   -21,    -8,   -11,    -8,    -8,    10,   -12,    -9,   -11,     2,     0,    -4,    -8,   -18,   -23,   -10,   -21,   -11,    -4,   -16,    -2,   -46,   -56,   -65,   -30,    15,   -10,   -15,    -6,     4,     3,    -4,   -10,   -24,   -17,   -17,   -12,    -1,     4,     7,    16,    -7,     0,     3,   -13,   -10,     6,     7,     1,   -34,   -56,   -25,   -12,     1,    10,    -6,   -11,     8,    16,    -6,    -7,   -20,   -16,   -24,    -6,     0,     2,    -5,    14,     9,    -2,   -11,   -10,   -18,    13,    29,    -1,   -33,   -24,   -19,   -23,   -28,    -4,     6,    -2,     4,    14,     4,    -8,   -14,    -2,   -22,    -5,     0,     1,    -7,     8,    15,     4,   -31,   -11,     4,    22,    37,     1,   -16,   -29,    -9,   -22,   -48,    -3,    -3,    -6,    18,    10,    18,   -13,   -17,    16,   -18,   -19,    -3,     1,    -3,     9,    10,   -16,   -23,   -13,    -3,     8,    18,    17,   -22,   -13,   -18,   -12,   -59,    -3,    -9,    -8,    14,    -8,    12,   -11,   -26,   -10,   -41,   -10,     0,    -5,   -12,     6,     5,   -12,   -20,    -6,    -2,    10,    18,     5,    -6,   -31,   -42,   -76,   -32,    -2,   -18,    -6,     8,   -11,     1,     2,    -9,   -15,   -30,     1,     2,    -2,   -10,    -2,    -4,   -18,   -22,   -16,   -14,     9,    20,     6,   -10,   -27,   -57,   -60,   -40,   -22,    22,     0,    15,    -8,    -2,    -1,   -14,   -15,   -21,    -7,    -4,     5,    -9,    -5,    -5,    -8,   -24,   -16,    -8,    26,    10,    -7,     4,   -13,   -26,   -19,   -10,    -7,     1,    -2,    10,    -2,   -14,     4,     3,   -38,    -9,     0,     4,     4,    -2,   -11,     9,    18,   -28,   -16,   -14,     1,    11,    22,   -18,    -6,    22,     1,    -9,    -6,     4,   -13,     2,     7,   -16,    11,     4,   -29,    12,     4,    -2,     4,    -1,    -4,    -6,    -1,   -36,    -8,   -18,   -11,     3,    14,    19,    19,    13,    17,   -17,   -12,    -6,     3,    14,     3,     2,     7,     7,    -4,    10,    14,     0,     0,    -1,    -7,   -12,    -5,   -16,    -8,    -9,    -1,   -11,    15,    -3,    11,    15,    -3,     7,    -8,     1,    11,    16,     8,     5,     9,    -4,     2,    10,     8,    -1,     2,    -4,   -14,     1,    -5,   -23,   -33,   -11,    13,    -4,   -10,    -5,    18,    12,    24,    33,    33,     9,   -18,   -16,    -7,    -4,   -13,     5,   -19,    -8,     1,    -1,    -4,    -7,     2,    13,    -7,   -16,   -14,   -23,   -10,    -9,   -12,    -9,    -8,   -12,     0,    -2,     5,    -3,   -16,    -7,     1,     1,    -8,    -6,    -2,     2,     0,     3,     4,     4,    -2,    -5,    -1,   -10,    -2,    -5,    -3,    -4,    -7,    -6,    -9,    -2,   -36,   -27,   -29,   -15,   -20,   -24,   -16,   -14,    -3,    -5,     4,     1,    -1,     1,    -4,     3,    -1,     0,   -14,   -20,    -2,    -5,    -1,    -9,    -7,    -5,   -18,   -23,   -19,   -18,   -29,   -31,    -6,   -26,   -19,    -4,    -3,    -5,    -5,     0,     4,     1,     5,    -5,    -2,     4,     3,    -3,     2,    -4,    -4,    -5,    -6,     2,   -10,    -5,    -3,    -4,    -4,    -4,     0,    -3,    -9,    -7,    -5,    -3,     1,    -1,    -2),
		    71 => (   -3,    -5,    -4,    -3,    -2,    -1,     1,     0,     1,    -5,    -2,     2,     2,    -3,     4,     2,     2,     2,     5,     1,    -5,     1,    -3,    -5,    -3,     4,    -5,     4,    -3,    -3,     2,     3,     2,     2,     3,     3,    -5,     2,    -3,     2,    -3,    -2,    13,     5,    10,     0,    -6,    -4,    -4,     3,    -3,    -4,    -1,     3,    -4,     2,    -3,     4,    -2,    -2,    -4,     3,     2,     3,   -16,   -17,   -10,    -9,   -23,   -12,   -17,     0,    23,    -2,    -7,    -6,   -15,   -37,   -25,   -17,    -7,    -8,     0,    -3,     3,    -3,    27,     2,     1,    -8,    -8,    -3,   -16,   -24,   -27,   -34,    -2,     3,   -33,    -9,    16,    18,    19,    17,    19,    21,    -8,    -2,    -6,    -2,    -2,     5,     2,    -3,    21,    22,     6,     9,     2,    -2,     9,     0,     8,    -3,    -2,    10,   -18,   -25,    -3,     7,    12,    20,   -11,    17,    -9,     3,    -5,   -16,   -22,    -9,     4,     3,    12,     4,     6,    10,    -1,    -4,   -16,   -11,   -11,     2,    18,     1,    14,    16,     6,   -23,    -2,    12,    10,     9,     7,     5,    -5,   -17,    -4,   -10,    -2,    -1,   -15,   -14,    -5,     7,     3,    -3,   -43,   -63,   -27,     2,    -6,   -12,    -9,    -5,     2,   -25,    16,    -4,     4,    16,    10,     4,    -2,     1,   -11,    -6,     3,    -4,   -19,   -17,   -21,     8,     9,   -20,   -40,   -19,     0,   -15,    -5,   -18,    -4,   -21,   -14,   -10,    10,     5,    11,    24,     8,    -5,   -10,     2,   -21,    -4,    -2,    -7,   -26,   -18,   -27,    -8,    28,     5,   -32,   -14,     3,    -6,    20,    18,     2,    -7,   -12,   -16,   -23,   -30,     2,    13,    17,   -10,   -16,    -2,   -22,    -1,    -1,     0,   -14,   -22,   -16,    -2,     4,    17,    11,     3,   -21,   -11,    -9,    11,     3,    -2,   -18,   -16,   -28,   -40,   -16,    -6,     7,    18,    -7,    25,    20,    -9,    -3,    -8,   -16,   -10,   -12,   -13,   -21,   -12,    14,    -9,   -24,    -8,     4,    20,     5,   -19,    -6,     2,   -20,   -10,   -27,   -33,    14,    16,   -12,    20,    17,    17,    -1,    -1,    -6,    -5,   -11,   -13,   -20,   -19,   -27,   -32,   -27,    -2,     5,     0,    -8,   -20,   -17,     1,   -24,   -19,   -11,   -15,    13,    17,   -10,    18,    11,    30,     4,     4,    -7,   -10,     1,    -4,    -1,    -1,   -20,   -10,    -4,     3,    17,    16,    -4,    -8,     3,    23,   -28,   -26,   -10,    -9,   -12,    -5,    -1,    25,    31,    37,    -3,     2,    -2,     0,    -2,    11,     8,     4,    18,    19,    -9,    -7,    -6,   -27,    -2,    -5,     4,     5,   -37,   -35,   -23,   -20,   -23,   -34,   -22,    33,    26,    -2,     5,    -3,     1,     7,    -7,    11,    12,    -6,    38,    33,    12,   -21,   -31,   -25,     4,    -4,    18,    -2,   -17,   -30,   -12,   -18,   -15,    -7,    -3,    -2,     3,     0,    -1,    -3,     1,    -8,   -12,    -9,   -20,    10,    15,    34,     1,   -11,    -9,    -3,    -4,    -3,    11,    -3,    -7,   -22,   -22,   -26,   -19,   -19,   -24,    -2,    -1,    -9,     2,     2,     2,   -12,    -1,     8,   -18,    -1,    14,     8,     6,   -20,    -3,    -5,     4,   -25,     0,   -10,   -20,   -39,   -26,   -39,   -24,   -20,    -2,   -25,   -14,    -5,     5,    -1,    -2,   -13,    -1,     8,   -10,   -25,    -8,   -19,   -25,   -45,     6,    18,     5,    -3,     1,   -19,   -38,   -31,   -14,   -25,   -19,   -10,    -7,   -14,   -17,   -27,     9,    -2,    -7,    -3,   -21,   -18,   -28,   -34,   -35,   -57,   -44,   -49,   -21,    -5,    21,     4,     3,   -11,   -33,   -18,   -16,   -14,   -14,   -14,   -21,   -10,   -17,    -7,     1,    -3,     3,   -14,   -16,   -42,   -16,   -29,   -12,   -31,   -35,   -49,   -32,   -23,    23,    18,     2,    -4,   -18,    -8,   -20,   -14,    -1,     3,    -8,    -8,   -11,    -1,    -3,     2,    -7,     8,    14,    -7,     7,   -10,   -14,    12,    11,     1,     5,   -26,    25,    18,    17,    11,    33,     4,    17,   -17,   -21,    -3,     8,   -12,    -9,    -2,     8,     0,   -11,    17,    24,    13,    21,    19,    -2,   -10,     4,    -8,   -21,   -17,    10,    12,    24,     1,    26,     8,    23,     7,   -33,   -18,   -10,    -4,   -17,     0,     9,     7,   -34,   -17,    31,    42,    25,    13,     4,   -14,   -23,   -13,     1,   -11,    -6,    40,    16,   -11,     6,     3,    10,     4,   -17,   -19,   -13,    -3,     1,    -1,     4,     5,    -7,   -15,     5,     2,    16,   -20,   -29,   -12,   -33,   -25,     5,    -2,     0,     9,     4,     1,     4,    -6,     3,   -13,     0,    -7,   -10,   -21,    27,    -2,     3,     2,     0,    -8,     2,    -2,    -7,    -7,   -19,    19,    17,     4,    -9,   -34,   -30,     7,    -6,    12,   -20,   -52,   -24,   -18,   -27,   -19,   -25,    32,    35,     5,    -3,     1,    -4,    -6,    -1,    -4,   -10,    -5,    -6,   -12,   -15,   -28,   -22,   -44,   -21,   -33,   -25,   -49,   -34,   -24,   -36,   -11,    -7,    -8,     0,    -5,    -8,     0,     0,     0,    -1,    -3,    -4,    -7,    -2,    -9,    -2,   -11,    -1,     0,   -34,   -25,    11,     7,    21,   -33,   -11,    -9,     0,    -8,    -1,     2,     5,     0,     4,     5,    -3,    -1,    -1,     0,     5,     5,    -3,     0,    -5,     5,   -10,    -9,    -5,    -6,   -12,   -11,    -9,    -1,     4,     3,    -4,     4,    -1,     1,     1,     0,    -3,     3),
		    72 => (   -4,    -2,    -1,    -5,    -2,     5,    -2,     2,     2,    -1,     3,     3,   -11,   -11,     7,     4,     4,     5,    -5,     3,    -1,     4,     0,     3,    -3,     2,    -2,    -1,    -2,     0,     1,     1,     1,     2,    -6,     0,   -22,   -14,   -21,   -28,   -19,   -27,   -13,   -18,    -7,   -13,   -19,   -40,   -28,    -9,    -7,    -9,     5,     1,     1,     3,    -3,     0,    -6,    -5,   -17,    -2,    -3,   -26,    -9,    23,    20,    -3,    -6,   -41,   -33,   -53,   -37,    -9,     1,    -8,   -45,   -13,   -16,    -6,    11,     4,    -3,     4,     0,     2,    -7,   -20,    -9,     5,     2,     0,     9,     9,    15,    -1,   -22,   -50,   -37,   -42,   -42,   -34,   -37,   -33,   -37,   -28,   -18,    -7,     2,     1,     5,     2,     3,    -4,   -14,    -2,     3,   -10,    12,    11,     4,    -7,    17,     3,   -15,   -44,   -38,   -31,   -36,   -22,   -35,   -35,   -22,   -26,   -17,   -15,     1,    -3,   -16,    -7,    -4,     3,   -10,     0,    11,   -15,    22,    21,    23,     2,    13,   -12,    10,    -1,   -17,    -3,   -44,   -44,   -31,   -19,   -11,   -22,   -29,    -9,   -17,    -5,    -3,    -9,    -4,     1,    -3,     3,     9,    25,    16,     4,    14,    17,     0,    -5,    -4,    12,    -4,   -19,   -22,   -23,   -23,   -11,    -9,   -22,   -22,   -17,   -27,    -9,    -8,    -8,     0,    -2,    -1,   -10,    -4,    -4,   -18,    -9,     2,     6,   -21,    -2,    -6,    -5,   -14,   -16,   -21,    -6,   -23,   -27,   -25,   -33,   -36,   -39,   -28,   -17,   -16,   -10,   -16,    30,    -6,     1,   -28,    -8,     7,    -7,     2,   -10,    10,    -9,   -12,    14,    14,     3,    -9,    -8,   -18,   -21,   -41,   -43,   -35,   -34,   -39,   -16,   -22,   -10,    -4,   -14,    -9,     9,   -32,    -5,     1,   -11,    -1,    -2,     7,     3,     6,     3,    41,    12,    -6,   -18,   -24,   -20,   -27,   -25,   -52,   -13,    34,   -29,   -10,   -13,     0,   -11,    -8,    -4,   -38,    13,    -2,    -1,    -1,   -15,   -17,    -8,     5,    -7,     9,    26,    20,   -15,   -23,   -14,   -15,   -26,   -26,     5,    20,   -15,   -22,   -19,    -1,    -3,   -28,   -11,   -15,   -11,   -11,    -8,   -12,     0,     7,    28,   -16,   -25,    -5,     8,     2,    -7,    -4,   -21,   -25,   -36,   -20,     3,    -5,   -21,   -39,    -4,    -3,    -5,   -33,    -5,    -3,     9,   -21,   -38,    -5,   -13,   -20,   -12,    -3,    -1,   -11,    -4,    11,    -5,    -3,   -26,   -21,    -7,     5,   -33,    -9,   -12,   -18,     3,    -3,    -5,   -26,    -1,    -6,    -8,   -30,   -40,    -9,   -16,   -29,   -17,   -10,     2,   -13,    10,     2,     5,   -13,   -15,     8,    24,    31,     5,    -9,    -6,    20,    20,     3,    -2,    -6,    -8,   -22,    -2,   -35,   -25,   -10,   -23,    -8,   -11,     0,     7,     5,     8,    12,    -1,   -14,     0,    10,    25,    15,    -4,    -8,     1,    40,    20,    -1,    -7,    22,   -17,    -5,    -3,    -5,   -20,   -12,    -4,     5,     1,    18,    28,    10,    13,     0,    -6,    -6,     2,    13,     3,   -13,   -21,     0,     7,    11,    24,     3,     1,    23,    -5,    13,   -18,     3,    -5,   -32,    -8,     6,    18,     3,    14,    12,    11,    22,    12,     2,    11,    -2,    10,     9,    11,     8,    14,    -5,    23,    -5,    -2,    35,     5,    19,   -10,    18,     2,    -8,     4,    12,    15,    -2,     3,    17,    16,    18,    13,    18,    26,    16,    20,    -8,     5,    -1,   -10,   -26,    22,    -3,     2,    15,    12,    10,     8,    27,    -3,   -14,     4,    14,    16,   -11,     6,    -8,    12,     7,     3,    16,     9,     4,    16,    13,    19,    31,    16,   -19,    15,     1,   -18,     2,    28,    -4,    17,    12,     7,    -2,    20,     5,    -4,   -16,   -12,    -6,    15,    -1,    -1,    -9,   -13,   -14,     0,    18,    31,    18,    10,    17,    36,    -2,    -8,     6,    20,     2,    -6,     4,    -9,    10,    -4,     1,    -3,    -4,     2,     5,    -1,   -25,   -36,   -31,   -30,   -26,    -7,   -14,    -7,    -8,   -25,    14,    -2,     4,    -1,    -4,    11,     8,     6,    30,     1,    -1,    -3,    18,   -16,     6,   -11,   -14,   -15,   -47,   -70,    -9,   -14,   -23,   -28,   -30,   -41,   -41,   -21,   -19,    -1,     5,     3,    -2,    -2,    -2,    10,     6,   -13,   -14,   -16,   -21,    -9,   -10,   -19,   -16,   -43,   -67,   -63,   -19,   -11,   -25,   -38,   -46,   -34,   -34,   -28,   -45,     0,     3,    -5,     4,    -5,    -6,    -9,   -12,   -20,    -1,    -1,   -29,   -32,   -58,   -49,   -65,   -53,   -62,   -59,   -41,   -44,   -41,   -44,   -38,   -53,   -41,   -23,   -42,     4,    -1,     4,   -13,    -4,   -47,   -13,   -30,    -8,     4,   -22,     3,   -14,   -90,   -64,   -56,   -47,   -53,   -59,   -50,   -48,   -46,   -48,   -37,   -38,     6,    16,    15,     0,    -2,     1,    -2,     2,   -12,    -9,    -2,    -7,   -35,   -47,   -52,   -32,   -51,   -47,   -33,   -40,   -41,   -31,   -24,   -41,   -42,   -35,   -10,   -10,     0,     8,    10,     2,    -1,    -4,    -4,     2,     0,   -15,   -25,   -25,   -36,   -45,   -33,   -11,   -14,   -16,   -24,    -9,   -19,   -16,    -9,   -29,   -15,   -10,   -18,    -4,    -4,     1,     1,    -3,    -3,     1,     2,    -4,    -1,    -3,    -5,    -1,     4,    -7,   -12,    -2,    -7,   -17,   -10,    -2,    -9,    -8,   -14,    -8,   -11,   -11,   -10,    -4,     5,     5,    -1,     0),
		    73 => (    4,     1,    -4,     2,    -4,     3,    -2,    -4,    -4,     1,     2,     5,    -6,    -3,    -8,     0,    -2,     4,    -4,    -5,     3,     2,     1,     1,     3,    -5,    -1,     0,    -3,     3,     3,    -1,     1,     0,    -3,     1,     0,     1,    -5,    -5,    -4,    -7,   -13,   -10,    -7,    -6,    -2,     2,     0,     1,     3,     0,    -3,    -2,     4,    -1,    -3,    -1,    -3,    -1,    -2,     2,     1,    -5,    -8,   -14,   -40,   -39,   -39,    -8,    -8,    -1,    -6,    -6,     3,     0,   -12,    -3,     0,    -9,    -4,    -1,    -1,     0,    -3,     0,    -1,    -1,     0,    -8,    -5,    -1,     6,     1,    -6,   -22,   -14,   -21,   -28,   -31,   -29,   -12,    -9,    -5,    -8,   -10,   -15,   -20,     0,     0,    -5,     1,    -3,    -1,     4,     2,     0,    -3,    -8,   -29,   -21,   -52,     6,    18,    -4,    -4,    16,     4,     0,    -4,    -2,    -1,    -5,    16,    32,   -21,   -22,   -19,    -2,     0,    -2,     0,     3,    -3,     1,   -17,   -12,   -17,   -38,   -41,   -15,    18,    14,   -18,    -8,   -10,     0,   -13,   -10,   -16,     2,   -19,    -7,   -14,   -13,   -46,   -15,    -4,     0,     2,    10,     7,     0,   -14,     5,    -9,    -5,    11,    26,     7,    -4,     9,    -6,     6,     9,   -19,    -8,   -23,     2,     0,   -15,    -2,   -11,   -22,   -33,   -10,     5,     4,     3,    -2,     4,   -46,   -36,   -16,     4,     3,    -1,   -21,     6,    32,     2,   -14,   -16,    -6,     1,    -7,    -7,   -14,    -9,   -23,   -34,   -21,   -25,    -3,    -1,    -3,    -3,    -8,     0,   -32,   -23,     2,     5,     5,   -10,    -7,    16,    14,    -4,    -9,     3,    -9,    -7,    -3,    -4,    -5,    -1,   -13,   -60,   -18,   -40,     5,    -5,    -7,     3,    -9,   -19,   -18,    -8,    11,    -4,     5,    12,    24,    15,    -6,    -5,   -13,     8,    14,   -10,     3,     5,    -4,     7,     5,   -48,   -18,   -23,   -20,     1,   -11,    -3,    -5,   -10,   -19,    -7,   -19,     9,     2,     8,    25,    14,   -23,   -27,   -10,   -13,    -9,   -16,     6,    21,   -16,     5,    -2,   -45,   -38,   -35,   -16,    -4,   -15,     0,    10,    23,    15,     6,     0,    22,     4,   -23,   -26,   -88,   -34,   -14,   -18,   -13,    -4,   -13,     4,    14,    26,    -3,    12,   -37,   -26,   -16,     3,    -2,   -10,    40,     7,    28,    18,     1,   -32,   -26,   -43,   -44,   -60,   -45,    -5,     2,    -9,    -8,   -18,   -11,    -4,     7,    18,    16,    13,   -25,     6,   -13,     0,    -2,   -15,   -19,   -24,   -27,   -23,   -19,   -68,   -60,   -46,   -25,   -15,     4,    24,    24,   -15,     2,    -4,    -7,     2,    -4,    -8,    -8,    -4,   -27,   -18,   -22,    -7,     0,     5,    12,   -11,   -19,   -52,   -51,   -59,    -7,    17,     9,    -9,    -1,    13,    -2,     6,    -5,    12,     1,   -19,   -23,   -13,   -13,     2,   -16,   -36,   -22,    -7,    -5,     2,     0,    -5,   -26,   -56,   -73,    25,    24,     4,     6,    10,    21,    20,    18,     5,    -4,    -3,     3,    -5,   -29,   -18,   -34,   -14,   -16,   -21,    22,    -6,    -3,     4,    11,    -9,   -11,   -20,    -8,    -9,    13,    18,    19,    21,    17,    14,    17,    -4,    -1,   -12,    -3,   -14,   -33,   -22,   -21,     3,   -10,   -13,    -7,    -7,     4,     4,    10,     7,   -25,   -25,   -12,   -18,    -6,     8,    29,    11,    29,    26,     6,   -27,   -19,     1,    -7,    -2,   -33,   -23,   -17,   -12,   -37,   -14,    -4,    -3,    -9,    -6,     3,    10,   -23,   -43,   -48,   -15,   -23,    -2,    11,    20,    26,     4,     1,   -11,   -12,   -21,     9,    -3,     4,   -12,   -13,   -32,   -38,    -6,    -4,    -4,    -4,   -13,     2,    -2,   -36,   -34,   -40,   -36,   -48,   -35,   -43,   -17,   -31,   -11,   -22,   -11,    16,    10,    20,     3,   -17,     7,   -17,   -34,   -38,    -2,   -18,    -6,     3,   -12,     7,    25,   -10,    -3,   -38,   -61,   -65,   -97,  -128,   -95,   -75,   -27,    -3,   -12,    -3,    17,    24,    14,     5,    -9,   -17,   -45,   -35,   -23,    -6,     4,    -6,    -4,    19,    41,    25,     0,    -4,   -25,    -5,   -19,   -20,   -30,   -21,   -15,     1,     9,    -1,    -1,    12,     0,    12,    -5,   -12,   -30,   -23,    -9,   -11,     5,    -3,     2,     5,    23,    42,    39,    29,    18,    16,    10,    22,     9,    -8,     5,     5,     6,    11,    -4,    -6,    -2,   -12,    -8,   -22,   -14,   -24,   -14,    -2,     0,     3,     4,     4,   -10,    28,    28,    25,    21,     4,    -7,    11,    -1,    16,    28,    -1,    14,   -29,     5,    -3,   -19,    13,     4,    -7,    -7,   -25,   -16,    -3,     5,    -3,    -2,     6,    18,    36,    -6,    19,    16,     2,     3,    14,    16,    11,    13,    -2,    -5,   -11,     7,   -52,   -14,    11,    13,    19,    19,   -32,    -9,   -13,     1,     3,    -2,     5,   -20,     1,    54,    35,    29,    12,    17,     2,    -8,     3,    -7,   -20,    -9,    -7,   -19,   -53,   -11,   -15,   -33,   -13,   -40,   -24,   -13,   -17,     4,     2,     4,     0,   -16,   -31,    -1,     3,    -7,    -6,   -26,     0,     3,   -10,     4,     0,   -27,    -3,    12,     9,   -13,    -7,   -11,     4,    -3,    -4,    -2,     3,    -1,     5,    -3,    -5,    -1,    -3,   -12,    -4,    -3,    -3,   -30,   -26,   -21,   -14,   -18,   -19,   -19,     1,    -3,    -9,   -21,   -19,    -4,   -16,     1,    -4,    -2,     0,    -1),
		    74 => (   -2,    -1,    -5,     0,     1,     4,    -1,     2,     5,     3,     3,     5,    -4,   -16,    -3,    -1,    -4,    -1,    -5,     5,    -3,    -4,    -1,     2,    -1,     5,    -3,    -1,     0,    -1,     5,    -4,     4,     4,   -19,   -18,    -7,   -17,   -30,   -17,   -36,   -22,     9,   -55,   -49,   -35,   -10,    -2,   -23,    -4,     0,    -8,    -5,     2,     2,    -3,    -1,    -3,    -8,   -21,   -31,   -21,   -10,   -28,   -18,   -18,   -48,   -62,   -47,   -11,     7,   -15,   -28,   -23,   -32,   -42,   -42,   -27,   -28,   -34,    -9,   -21,     3,    -5,    -4,    -1,   -13,   -39,   -63,   -21,   -24,    -3,   -43,   -50,   -30,   -42,   -72,   -24,     7,    -5,   -19,   -28,   -38,   -12,   -10,   -20,   -12,   -35,   -41,   -17,    -2,     2,     0,     0,    -7,   -55,    -6,     2,     3,     9,    -3,   -29,   -21,   -20,    -6,    14,    18,     8,     4,    13,    20,     1,   -11,     4,    41,     2,    -4,    -8,   -38,   -11,    -3,     2,   -14,   -25,     5,    12,     8,    34,    18,    14,    13,    -6,    12,    21,    32,     8,    -2,    23,     8,    28,    -6,    18,    18,    31,    31,    17,   -36,     0,    -3,     2,   -12,    -7,    21,    14,     5,    35,    29,    31,    19,    11,     6,    32,    40,    52,    31,     7,   -14,     0,    13,     2,    -3,    31,    40,    12,     8,   -21,     0,   -20,   -18,    10,    22,    11,    22,    36,    16,    74,    48,    66,    36,    40,    37,    34,    20,    23,     8,    26,    11,   -11,    -8,     4,    16,   -16,    42,   -29,   -21,   -24,    26,    12,    12,     2,    28,    15,    -2,    62,    36,    40,     6,    -8,    -3,    10,   -12,   -12,   -12,    -4,     6,     4,   -28,   -10,     0,    11,    19,   -32,     2,   -10,    20,   -17,     3,   -15,   -21,   -10,   -10,    -1,    11,   -27,   -10,     4,    -8,     4,   -20,    10,    -5,    -7,    -6,    -7,   -34,     0,    -7,   -20,   -19,   -17,     3,   -13,    11,   -11,   -11,   -23,   -41,   -18,   -19,     6,   -11,   -32,     0,   -26,   -22,   -11,   -10,    -2,   -26,     0,   -32,   -17,    -8,   -20,   -44,   -13,    -3,   -25,     5,   -22,    11,   -17,   -21,   -17,    15,   -31,     4,   -13,   -28,    -9,    -4,    -9,   -15,    -5,     3,    17,   -22,   -20,   -53,   -22,   -15,   -33,   -53,   -13,   -22,   -41,    -3,     5,     4,   -17,   -29,    -8,    -4,   -20,    -4,     3,   -15,     9,    31,    15,   -29,     1,     6,    12,    -7,   -13,     0,    16,    -7,   -21,     4,    25,   -20,   -34,    -1,   -10,   -28,   -26,   -29,    -3,     2,    29,    17,   -13,     9,    29,    36,    -4,    10,     5,     0,    15,    17,    -5,     2,   -16,   -19,    -9,     3,    14,   -10,    -4,    -5,    16,   -50,   -34,    -1,    -1,    -1,    46,    26,    15,    26,    19,    12,    -8,   -11,    -4,     7,     6,    -9,    -4,   -21,   -26,    -6,    -4,    -1,    20,   -28,    -4,    -5,     4,    22,     5,    25,    -2,    17,    22,    27,    13,     4,     5,    23,    16,     5,    -3,    12,    24,    -6,   -11,     2,     2,    23,    14,   -10,    -3,   -18,   -28,     3,     1,   -31,     7,   -13,   -13,   -12,   -10,     1,    -1,    14,    14,     2,    -1,     6,    -4,     8,    10,     5,    11,    24,    17,    17,    -4,    11,     5,   -17,   -12,     1,    -2,   -20,   -26,     1,     2,   -14,    24,     4,    -5,   -27,   -11,     3,   -18,    -5,   -18,    20,    -5,    -8,     6,     1,    18,     7,    33,    10,   -40,    -7,   -13,   -21,    -4,    -7,     1,     3,    19,    10,     3,   -22,    -9,   -26,   -19,    10,   -12,     3,   -12,   -15,   -31,    -9,    25,    42,    26,    16,    28,    19,   -10,   -18,   -25,     1,   -19,   -28,    56,   -14,   -10,   -16,   -28,   -11,   -24,   -30,   -30,    -3,     2,     9,    14,     6,   -32,    -1,    13,    14,    10,    18,     3,     6,    -3,    -7,   -20,     3,    -6,   -14,    14,   -18,   -27,   -30,   -33,   -17,    13,     2,     3,     0,    -5,     1,    11,    18,    -4,    20,    19,    30,    19,     8,    -6,   -30,   -34,   -15,    -4,    -8,    -3,   -21,    18,    13,   -12,   -20,   -16,     5,     8,     0,     9,   -21,   -10,    -7,    13,    15,    12,    -4,    25,    55,    43,    44,    13,   -10,   -47,   -32,     1,    -8,    -8,    -9,   -27,   -58,   -31,     0,    10,    24,   -10,    30,     4,    -6,    -1,   -22,   -13,    22,    21,    -1,    42,    48,    53,    34,    28,     2,    -1,    -9,    -6,     5,     3,    -1,   -38,   -50,   -92,    16,    25,    39,    25,    44,    33,    14,     1,    -7,   -13,     8,    -3,    20,    46,    45,    19,   -19,    20,     0,    29,    -9,    -1,     1,     3,     2,   -14,   -48,    -8,    38,    42,    11,    30,     5,    35,   -11,    -2,    -2,   -32,   -15,   -17,    24,    41,    -1,   -14,    -7,    -3,   -25,    24,   -24,    -2,     1,    -1,   -15,    -1,    41,    56,    18,   -15,   -11,     5,    21,    18,   -20,    11,   -26,     8,     4,    -6,    -7,    -5,    -7,   -10,    -9,     5,   -10,   -27,   -20,     4,     2,    -5,     0,   -36,    62,    53,    31,   -11,   -22,   -35,   -62,   -12,   -18,   -20,   -12,   -45,   -48,   -32,    -8,    -3,   -36,   -73,   -65,   -17,     4,    -4,     5,     3,     0,    -5,     2,    -2,    -7,    -1,   -21,   -24,   -16,   -19,   -25,   -31,   -25,    -8,   -19,    -8,   -39,   -58,   -46,   -27,   -30,   -14,   -21,     2,     5,     1,     0,     0),
		    75 => (   -3,     4,    -4,    -1,     0,    -2,    -3,     3,    -2,    -4,     1,    -1,     4,     2,     1,    -4,     5,     1,     3,    -1,     3,     2,    -1,    -1,     4,     2,    -3,    -3,    -3,     0,    -4,    -1,    -4,     4,    -1,    -1,     4,     3,    -4,    -5,    -8,   -15,   -11,    -7,    -6,   -15,   -11,    -1,    -2,    -6,     2,     2,    -5,     5,    -3,     2,     1,    -2,    -4,    -4,     1,     1,   -11,    -7,   -24,   -25,   -29,   -30,   -15,   -19,   -47,    -7,     6,     5,    -4,    15,    26,     1,     0,     7,   -12,    -2,     4,     0,     1,     1,    -5,     7,    13,   -20,   -24,   -25,   -15,    -8,    -8,   -13,     3,     7,    15,    17,    14,    -2,   -17,   -13,     5,    15,     4,    13,     6,     4,     6,     5,     3,    -3,     0,    11,     0,    -2,    13,    20,     6,    20,     1,   -24,   -15,    -2,     9,    20,    23,     3,    -1,   -15,    -4,     1,    11,    14,    11,    15,    -9,   -14,    -5,    -2,     3,     3,   -13,     1,    19,    10,    13,     2,    -5,   -19,   -22,    -5,     1,    -6,    -1,    -1,    -3,    25,    18,    -1,    16,    16,    15,    12,   -11,   -12,     2,    -5,   -21,   -14,     9,    13,    27,     8,     2,    -3,     0,   -12,   -15,    -7,    -2,    -1,    -5,   -11,     6,    26,    27,    19,    14,     8,    14,    14,    10,     5,    -4,     2,     2,   -17,     4,    32,     4,     6,   -12,    -6,    -8,    -4,    -8,   -11,    -2,   -12,    -1,    -5,    -7,     2,    12,    -5,    15,    13,    29,    17,    12,    14,    -4,   -15,   -17,   -28,     6,     1,     1,     3,   -10,     3,     1,    13,     9,     9,    -2,   -17,   -16,   -24,     5,     6,    -8,     2,    23,    30,    14,    21,    13,     7,    -1,    -7,   -35,   -25,     3,     5,     2,     2,   -11,    -7,    11,    16,    24,    18,    -8,   -10,   -20,   -19,    -8,     1,     9,    24,    29,    28,    23,     5,    19,     6,     3,    -2,    -6,   -37,    -1,    -1,    -3,    10,   -10,     4,    -1,    23,    31,     3,    14,     1,   -23,    -8,     2,    14,    27,    40,    38,    29,    27,    14,     2,   -14,     4,    -5,    -3,   -24,     8,    -1,     5,    10,    13,    -4,    -9,    22,    18,     2,    15,   -14,   -20,   -31,    24,    21,    37,    15,    17,    18,    25,    22,     4,   -16,     2,     2,     0,   -28,     8,    13,    14,    14,    25,    17,   -15,     0,     6,     2,     4,    -7,   -21,    -2,    12,    25,    14,     1,    -5,    15,    10,    10,    24,   -17,    -5,     0,    -3,   -31,     1,     9,    11,    21,    15,    21,    28,    12,    10,    -8,     1,   -20,   -12,   -10,     0,    21,    18,    20,    -1,   -13,   -13,    -1,    19,   -16,     4,     0,    -7,   -41,    -4,     5,    15,    18,    17,    13,    30,     3,     6,     2,     0,   -16,    -8,     8,    28,    22,    19,    15,    12,   -11,   -19,   -18,   -13,     1,     5,    -6,   -10,    -4,     8,    14,    -1,     7,    16,    24,    28,    -3,    -2,     2,    15,     3,    -1,    11,    17,    23,    13,    12,     7,     1,     4,   -20,   -12,   -26,    -1,    -8,   -18,    -2,    10,    36,     9,     6,    15,    16,    15,   -17,     3,     5,     3,    11,   -12,     3,     1,     4,    20,    36,    17,     1,    -9,   -20,   -15,   -32,    -3,    -2,   -15,     8,    13,    34,    23,    20,    25,    22,    -8,   -10,   -16,     1,    17,   -12,     3,    -4,    -4,    -2,    15,    10,    18,     4,    -5,   -21,   -35,   -37,    -1,     1,   -22,     4,     6,    30,    22,    17,    27,    22,    -2,   -21,   -33,     9,    11,     1,    -2,    -9,   -11,   -16,    -5,     1,    -3,     9,    10,   -15,   -42,   -23,     5,    -5,    16,     2,     7,    15,    16,    31,    21,    -2,   -12,   -12,   -18,    10,     1,     4,   -11,     4,    -5,     3,     3,    -2,    -2,    14,     6,   -16,   -45,   -19,     5,    -3,    11,     9,     8,     6,    17,    21,    26,     0,   -10,   -16,     3,     2,   -10,    -7,    -5,     3,    14,    14,    -7,     7,     9,    17,   -18,    -4,   -31,    -2,     0,     1,     3,     3,     5,    14,    18,    24,    23,    18,     1,    10,     6,     5,     0,    -6,    -1,    -2,     6,    15,    18,     2,     6,     4,   -20,    -1,   -19,    -4,    -3,    -2,   -22,    -2,     8,     5,    17,    11,    25,    14,     7,    24,    12,     3,     2,     3,    -9,   -11,    -9,     4,     6,   -12,    -8,   -11,   -27,     2,    17,    -3,     0,    -1,     6,     0,   -12,    -2,    11,    19,    12,     7,    -1,    12,    10,    11,     7,    -8,   -29,   -21,   -11,   -11,    -5,   -20,   -12,   -20,    -7,     8,    14,     2,    -5,    -4,    -6,     1,   -16,    -8,    14,     6,     6,    13,    14,    10,     5,    -7,     5,    -1,   -18,   -14,    -6,   -15,   -18,   -14,   -11,    -9,     5,   -33,   -11,     1,     3,    -1,     3,    16,   -30,   -24,    -3,     8,   -11,   -18,    18,     9,    10,     5,     0,     8,    11,    20,    15,    -4,    12,     6,    22,     6,     1,    -1,    -3,     0,    -2,    -4,     0,   -15,   -23,   -31,   -36,    -6,    -1,    -8,    -7,    18,    -4,     5,    16,    10,    10,     3,    -8,    -4,   -16,   -12,     4,   -19,     0,     0,     4,    -2,    -2,    -5,    -4,    -3,    -8,    -6,    -3,    -1,    -3,    -1,     4,     1,    -8,    -4,    -7,    -4,    -1,     3,    -3,   -12,    -7,   -25,   -19,    -7,    -3,     4,     3,    -2),
		    76 => (    2,    -1,     3,    -2,     0,    -2,    -5,     1,     3,     4,    -2,     2,     1,     2,    -2,    -4,     2,     1,     2,    -1,     4,    -2,     2,    -1,    -5,     2,    -3,    -1,    -2,    -4,    -2,    -1,    -2,     4,     6,     9,    15,     8,     5,    10,     9,     5,    -5,    -7,   -12,     3,    -2,    -2,    27,    11,     5,     8,     3,     2,     0,     1,     2,    -2,     6,     5,    23,     8,     0,    16,    20,     2,    -7,     1,    -1,     5,   -12,    -6,    -7,     8,    -1,     6,     9,    34,    41,    33,    30,    14,    -4,    -2,     2,     0,   -11,   -10,    -2,     0,     1,    -4,    -3,    -2,    -7,    -5,   -31,   -29,   -30,   -16,   -19,   -25,     7,    31,    31,    20,     8,    29,    30,     3,   -24,    -3,     4,     3,    -8,     1,    11,     5,   -10,   -14,   -16,    -3,    -9,   -14,   -27,   -36,   -40,   -31,   -13,   -17,   -13,     3,     4,    24,     2,    28,     9,    -8,    15,    18,    -5,    -2,   -12,   -15,    10,     5,    -6,    -9,    -6,    -3,   -17,   -23,   -25,   -23,   -18,    -8,   -12,    -5,     0,     2,    -7,     8,    16,    25,    29,    26,    33,    19,    -4,    -3,     1,    -3,     4,     6,    -7,    -4,   -15,    -4,   -16,   -15,   -11,   -17,   -31,   -34,   -28,    -6,    -6,     7,     1,    -7,     4,    21,    29,    16,    13,    28,     3,    -3,     2,    -2,    13,     6,   -16,    -3,    -2,    10,   -23,   -24,   -21,   -37,   -25,   -38,   -12,     2,     6,   -10,   -11,     4,   -12,   -12,     8,    16,    11,    30,    -1,    -1,    -2,    -7,    17,     1,   -26,   -12,    -7,    -4,   -30,   -32,   -38,   -36,   -30,   -22,     6,     3,     9,     2,     0,    -7,   -10,    -5,   -27,   -14,    24,   -16,     3,    -4,     0,   -13,    23,    -3,   -24,    -3,     7,    -5,   -27,   -33,   -35,   -35,   -20,     9,    11,     5,    -3,     5,    -6,   -11,    -9,   -20,   -25,   -17,   -13,    -8,    -2,    -4,    -1,    -8,    16,    -6,   -16,    -4,    -4,   -25,   -52,   -40,   -28,    -6,    -2,    11,    -9,   -13,   -26,   -33,    -6,    -9,   -18,   -21,   -17,   -14,   -12,   -16,     1,    -3,     5,   -12,     7,     4,   -27,   -24,   -22,   -51,   -30,   -28,   -13,     1,    11,     0,   -13,   -40,   -51,   -32,   -32,   -19,   -14,   -18,   -26,    -3,    -6,    -9,    -5,    -2,    -5,   -19,     5,    -7,   -20,   -26,   -31,   -30,   -33,     2,   -11,    10,    -3,    -8,   -13,   -27,   -45,   -32,   -26,   -15,    -8,   -10,    -2,    -7,   -16,    -7,     4,     3,    -3,   -12,    -4,    -5,   -17,   -19,    -1,    -9,   -10,    -6,     8,    12,    -8,     3,     2,    -1,    -7,    -9,    -5,   -32,   -18,    -3,    -3,    -1,   -17,    -5,     1,     0,     2,   -10,   -12,   -13,   -10,     3,    16,   -13,     4,    -8,    12,     3,     4,   -14,     8,    -1,    -5,     2,     3,   -20,   -36,   -30,    -3,     1,    -7,    -9,     1,     0,   -10,    -5,   -14,   -18,    11,     8,    -8,     5,   -10,     9,    18,    -2,    -6,    -9,    -3,     9,     3,   -13,   -23,   -24,   -32,   -14,    -9,    -6,    -5,   -14,     3,     2,    -9,   -12,     4,   -16,    -7,    -4,     5,     2,     0,     3,    10,     7,     1,     5,    -5,   -12,     6,     3,   -19,   -30,   -17,    -8,   -12,     3,   -10,    -7,    -4,    -3,   -11,   -20,    -6,   -21,   -16,     2,     6,    -3,    23,   -11,    -8,   -22,   -15,   -11,   -14,   -20,    19,    12,     3,   -17,    -5,   -10,   -13,    -9,   -12,   -24,     3,    -4,    -4,    -3,    15,    -8,   -18,    -9,    -1,     3,    -1,    -9,   -19,   -15,     0,     8,    -1,     0,    22,    32,    22,     0,    -8,   -14,    -7,    -1,   -23,    -3,    -1,    -3,     3,   -12,    11,   -11,   -13,     2,   -18,     8,    -5,   -19,    -7,   -26,     0,    15,     5,    10,    27,    20,    17,     3,   -20,   -14,    -3,     1,    -3,    -9,    -3,    -3,    -7,   -13,    14,     1,    19,    10,    -7,    -4,     1,    -9,    -9,     0,    26,     5,    -9,   -11,    -1,     4,     0,   -10,   -16,   -15,     1,    -2,    -3,     0,     3,    -3,   -14,   -11,     6,    -1,     1,     1,    15,   -15,     9,    21,    18,    12,     9,     1,    -4,   -13,   -13,   -18,   -25,   -22,   -16,    -6,    -2,    -3,     1,    -3,     0,     0,    -6,     2,    -5,   -10,   -35,   -10,    16,    -7,     2,    17,    27,    11,   -19,   -20,   -10,   -23,   -17,   -20,   -20,    -5,    -5,   -15,   -10,   -14,     2,     4,    -4,    -4,     1,   -11,   -15,    -7,   -19,    11,     9,     4,    11,    17,    15,     4,    -4,   -11,    -5,   -29,   -23,   -18,    -1,    -5,    -1,     2,   -10,   -12,    -4,     2,     2,     3,    -2,    -2,    -7,    -9,    -5,    -6,   -14,   -12,    -6,   -11,    -5,   -12,    -5,    -4,     6,     0,    -1,   -14,    -5,    -7,    -5,     3,     1,    -6,     1,    -2,    -4,     5,    -4,    -4,     0,   -17,   -21,   -22,   -12,    -7,    -3,     1,     1,    -4,    -5,     2,    -6,    -2,    -4,    -5,   -15,    -6,    -4,    -9,     0,    -2,     1,    -3,     4,    -5,     0,    -2,    -3,    -9,    -8,    -6,    -5,     0,   -10,    -8,    -4,    -1,    -1,    -1,    -3,     2,     0,     2,   -11,    -4,    -8,     0,     1,     4,    -3,     3,    -4,     2,     5,     3,     3,     4,    -4,     5,     4,     3,     3,     2,    -2,    -1,    -6,    -1,    -3,    -6,     2,    -1,    -5,    -8,     2,    -1,     0,    -4,     1,    -5),
		    77 => (    1,    -2,    -3,     2,     3,     1,    -5,     4,    -1,     1,    -3,     5,    -2,     5,     3,     1,     1,    -1,     0,    -3,    -3,    -5,     4,     3,     1,    -1,     4,     0,     3,     2,    -2,    -1,    -1,    -2,     0,     4,     3,    -1,    -7,    -1,    -2,    -3,    -5,   -17,   -22,   -14,     4,     4,     5,     0,     0,     0,     3,     0,     0,     5,     3,     4,     1,    -3,     0,     4,    -1,    -5,    -1,     0,   -13,    -8,    -2,    -3,    -4,    -4,     0,     1,    -5,     0,     0,    -2,     0,    -4,    -3,    -1,    -2,     3,    -2,     1,    -5,    -4,    -5,    -3,    -2,     3,   -12,   -12,   -11,   -15,    -7,   -11,     3,   -15,   -18,   -35,   -10,   -18,   -11,    -9,   -19,    -4,    -7,    -4,    -4,     4,     2,     0,     2,    -3,   -14,    -7,   -12,   -33,   -27,   -23,   -32,   -49,   -56,   -42,   -29,   -55,   -41,   -46,   -43,   -26,   -27,   -11,   -37,   -22,   -13,   -10,    -4,    -4,    -5,     5,    -5,   -20,    -4,    26,    22,    16,    35,    34,     1,    14,     5,    11,    -8,    -1,    -5,   -19,    -1,   -11,   -20,   -41,   -42,   -31,   -40,   -34,   -10,    -4,     3,     0,    -3,   -12,    -7,    14,    19,    27,    28,    -1,     5,    16,    24,    25,    31,     8,    27,    20,    14,    16,    19,     5,    13,    -2,    -5,   -12,     1,   -10,     0,     4,    -7,    -3,   -11,    -9,   -13,    20,    -6,     5,    -3,    18,    30,    29,    11,    18,    11,    28,     3,    10,    15,    -2,     2,    -4,     4,    -5,    -7,    -5,   -13,     8,    -1,    -7,    -8,   -22,   -20,   -17,   -28,   -25,   -28,    -2,     3,    -8,     3,     6,    -3,    11,    -7,     1,   -18,   -10,   -22,   -21,   -20,    -8,   -14,   -16,     0,    -2,    -6,     5,     1,   -17,   -29,   -22,   -46,   -15,   -28,   -18,   -15,   -22,   -12,   -20,     2,   -22,     1,    -5,   -17,   -12,   -13,   -18,   -15,    -5,   -16,    10,    -2,    -8,   -18,   -17,    -1,   -20,     0,   -13,   -21,   -13,   -26,   -15,   -41,   -49,   -50,   -13,   -10,     4,    -7,   -11,    -3,   -35,    -9,   -28,   -19,    -9,   -19,     9,    -2,    -4,   -17,    -2,   -15,   -16,   -17,   -30,   -39,   -33,   -52,   -35,   -57,   -34,   -26,    -9,    -1,    -7,   -13,   -13,   -11,   -10,    14,    17,   -14,   -31,   -17,    14,    -1,     1,    -9,     5,    -1,   -14,   -22,   -41,   -34,   -47,   -32,   -41,   -32,   -20,   -17,    -6,    -2,   -24,   -29,   -11,   -15,     3,     5,    -6,    -1,    -2,   -10,    14,     4,    -2,     7,     0,    -6,   -15,   -10,     2,   -18,    -3,   -14,    -7,    -8,     0,    -3,     3,    10,   -12,     2,    -6,    16,    17,    -6,   -19,   -15,    -1,   -18,   -16,    -4,    -1,     0,    -7,    12,     0,     8,    18,     0,     2,     5,    11,    15,    10,    11,    10,    10,     1,    10,    34,     0,     3,     9,   -35,   -21,   -13,   -13,     4,     1,     0,    -8,     3,    17,    13,    12,    20,    19,    -5,     8,    -2,    -8,     3,     0,     9,    22,    13,    -3,    -7,   -16,     4,   -12,   -40,   -41,   -26,    -4,   -10,     5,    -3,   -10,   -11,     4,     1,    -4,   -25,    -1,    -2,    -3,   -16,    -1,     5,     4,    18,     8,     0,    -2,    -6,     4,    -8,   -23,   -31,   -37,   -23,   -16,   -13,    -3,    -3,   -12,   -11,   -17,    -9,    14,   -18,    -7,    -3,    -8,    11,     1,   -10,     7,    -6,   -16,   -15,    -1,    -2,    12,    -4,     5,    -6,     7,    10,    19,   -26,     1,     1,    -4,   -12,     0,   -12,   -14,    -7,     0,   -23,   -14,    14,     7,    -9,    -5,    -5,   -40,   -27,    -5,     2,   -14,   -17,   -23,   -19,    -6,    14,    27,   -24,    -3,     2,     4,    -6,    11,   -17,    -3,   -30,   -32,    -7,   -14,     1,   -15,   -12,    -5,   -20,   -53,   -22,    -2,    -7,   -43,   -53,   -26,   -30,   -14,    17,   -13,    -8,     4,     6,     5,    -4,   -14,    -5,   -10,   -21,   -16,    -9,    -1,    12,   -14,   -13,   -10,   -23,   -31,   -15,   -43,   -40,   -16,   -22,   -25,   -13,   -29,   -34,    -7,    -4,    -2,     1,    -3,    -1,   -11,    11,     0,     4,    -9,     2,     3,    -2,    17,     7,   -11,    -6,   -16,    -7,   -24,   -17,   -34,   -23,   -11,    -7,   -16,   -17,    -6,     2,     2,    -2,    -7,    -7,    19,    -1,    -7,     6,    11,    -2,    -1,     2,    -1,    10,   -25,    -2,    11,    -1,   -11,   -31,   -39,   -25,    -6,    -1,   -25,    -8,   -12,     2,     3,    -3,    -7,   -33,    -3,   -22,     4,    -3,     0,   -13,    -7,    -4,     1,    16,   -10,   -10,   -27,   -30,   -19,   -18,   -36,   -17,   -18,    -1,    -2,    -2,   -13,    -2,     0,    -1,    -8,   -22,    -9,   -17,    -2,    16,     9,     4,   -22,     3,     9,    13,    -4,    18,   -29,   -31,    -6,    -6,   -30,   -32,   -24,     5,    -5,   -17,    -8,     4,     3,    -5,     5,     9,    10,     5,   -23,     6,    12,   -26,    -4,    12,    15,   -11,    -7,   -21,   -36,   -19,   -11,   -13,   -21,   -15,    -8,    -1,     1,    -6,    -1,     1,    -1,     3,     1,   -17,    -6,   -14,    -2,    21,    22,    14,     1,     2,    17,    16,    20,     0,    -1,     2,     3,     5,     3,     0,     1,    -1,     2,    -4,     4,    -3,     1,     0,    -3,     4,     6,     1,     2,    -3,     7,    -2,    -9,    -2,     6,     6,     5,     0,    -1,    -1,     6,     5,    -2,     0,     3,     7,     4,     3,     0,    -2),
		    78 => (   -5,    -3,     1,     4,     3,     4,    -2,    -1,     1,     0,    -2,     5,     2,    -3,     4,     2,    -2,     3,     1,     2,    -3,     0,     4,    -4,    -5,     2,     3,     4,     3,     4,    -4,    -3,    -4,    -4,     0,     0,     5,     2,    -1,    -4,     3,     2,    -3,   -14,   -25,   -18,    -2,     1,    -1,     0,     1,     4,    -3,    -5,    -3,     0,     3,    -4,    -1,     3,     5,     0,    -2,     2,    -7,   -13,   -28,   -21,    -7,    -4,    -6,     0,     1,    -7,   -10,    -5,    -6,   -12,   -19,    -8,    -9,    -7,    -1,     2,     0,     0,    -8,    -1,    -2,   -16,   -11,   -25,    14,     8,    -5,    -9,    -1,    -9,   -16,    -9,    -5,   -13,    -2,    -6,    -8,    -7,     1,     5,     0,    -7,   -13,     4,    -1,     2,     1,    -1,   -15,   -25,    -2,     1,    -7,   -24,   -23,   -29,    -9,    -9,    -2,   -21,    -8,    17,    18,   -10,    -7,   -11,   -16,   -13,    -2,    -9,     5,    -7,     4,    -5,    -3,    -3,   -15,   -19,     5,     4,   -14,   -26,   -20,   -15,   -18,    -5,    -7,    -1,     1,     3,    12,     6,     2,     0,    -8,    -4,    -3,    -5,    -4,   -14,     1,     4,   -12,   -24,    -5,   -20,     0,     4,    -2,    -2,   -15,   -13,     3,     4,    -1,     9,    -4,    -3,     2,     1,     3,     0,     3,    -2,    -1,    -1,    -3,     2,     1,   -21,    -9,    -1,   -13,    -9,     7,    -1,     4,     5,    10,    -1,     2,   -14,    -2,    17,     4,    -4,    14,   -13,    -3,    -2,    -5,   -10,    -7,    -8,    -5,    -5,    -8,   -11,   -10,     1,   -12,    -8,    10,     1,    -3,    -1,     5,    -2,    -7,    -8,    -1,    17,     9,   -19,     4,    -5,   -18,    -7,    -5,     2,    -3,     7,    -2,     2,     0,    -7,   -20,     0,    -5,   -25,     5,    -6,     6,    -2,    -2,   -17,   -12,    -6,    -3,    14,     6,   -19,     6,     1,    -4,    -1,    -1,    -8,   -15,    -3,   -11,   -25,     1,    -6,   -18,     5,    -5,   -22,   -21,     2,    -3,   -15,     3,     1,    -5,   -16,   -21,     7,   -13,     6,     2,     0,    -4,   -11,   -12,   -19,   -15,    -5,    14,   -18,     1,     3,    -9,    -1,   -11,   -22,   -20,     6,    -6,   -19,    -7,   -12,   -18,   -24,    -8,    12,    -1,     0,    11,     5,    -6,   -23,   -14,     9,    -1,     0,    20,   -20,    -4,     3,   -12,   -11,   -16,   -11,   -14,    -1,    -1,   -13,   -13,   -12,    -9,   -21,   -21,    13,    10,     5,    10,     5,    -1,     4,     7,   -13,    -7,   -10,    -8,   -29,    -3,     0,   -17,   -11,   -19,   -18,   -14,    -4,    -8,     1,   -26,   -18,   -26,   -29,   -13,    -1,    -6,     2,    16,     5,     2,     7,    -7,   -10,   -13,   -16,   -16,     1,     1,    -1,     2,   -11,    -2,   -11,   -23,    -9,    -6,     0,    -1,    -8,    -4,   -36,    -9,   -12,   -24,   -14,    -9,     2,    -1,    -5,   -16,   -16,   -14,    -5,   -46,    -6,     0,     4,     0,    -8,     0,    -1,   -12,   -13,   -10,     4,    -1,   -14,    -3,   -26,    -1,     1,    -9,    -2,    -7,    -9,    -8,    -6,    -9,   -13,    -6,    -3,   -41,   -15,    -1,    -2,    -3,    -6,     3,    -7,    -8,    -1,    -5,   -13,    -7,    -8,   -15,    -6,     8,     0,    -8,     2,    -8,   -10,   -10,    -5,   -12,    -9,    -5,     1,   -22,   -15,     3,     0,    -3,    -6,    -1,    -7,   -10,    -5,    -9,   -23,   -22,   -16,   -25,     3,    13,     8,    -7,   -16,    -4,    -2,    -2,    -6,   -11,    -5,    -1,    -4,     0,   -16,     1,     2,     0,   -11,    -1,    -8,    -6,     0,   -12,   -17,    -5,   -19,    -1,     9,     4,    -2,     5,   -16,     1,    -4,    -8,   -15,    -3,    -7,     4,    -2,     1,    -9,     1,    -4,   -14,   -15,     3,    -6,    -4,   -14,   -22,     0,    -6,    -9,     8,     7,     0,    13,    15,    -6,    -3,    -7,   -12,    -6,    -7,    -2,    -2,     0,   -23,   -19,     0,     2,    -5,    -3,     2,   -15,   -10,    -8,   -11,     7,    -2,    -8,    -4,    -7,   -17,     1,    -4,    10,     2,    -6,   -22,   -14,   -13,    -6,     1,    -5,   -18,     5,   -18,    -8,    -6,    -1,   -10,   -18,   -14,   -24,    -1,    15,    -1,   -19,     3,    -8,   -17,   -22,     0,    19,     3,     4,   -11,    -4,    -9,    -8,    -7,     1,   -21,     0,    -9,    -9,    -3,    -8,    -2,   -16,    -7,   -10,    -6,    10,     8,     4,     3,    -8,   -16,   -17,    12,    12,     1,    -3,    -7,   -19,   -16,    -8,    -8,    -4,   -14,     3,     1,     2,    -7,    -2,    -7,   -14,   -12,    -9,   -14,     0,    10,     9,    27,     8,     3,     0,    24,     0,    -6,   -24,   -11,    -8,   -11,    -5,    -6,    -1,   -25,     2,     1,    -3,    -3,    -7,    -1,    -6,   -16,   -11,   -14,    -8,   -11,   -12,     3,    -1,     4,     5,    12,   -24,   -23,   -20,   -18,    -7,    -2,    -5,   -17,    -4,    -4,     1,    -1,     4,   -13,   -11,    -4,     1,    -8,   -15,   -15,   -14,   -14,   -35,    -4,     6,     3,    14,   -24,   -33,   -23,   -15,    -3,    -6,     0,     2,    -1,    -9,    -8,     2,    -1,     2,     4,    -4,     3,   -11,   -11,    -8,     0,   -13,   -19,   -23,   -20,   -27,   -36,   -18,    -8,    -1,    -3,    -7,   -28,   -16,   -14,    -4,     1,     4,    -1,     2,     3,    -4,    -2,    -2,    -4,    -1,    -8,     1,    -6,    -3,    -6,     1,     3,   -11,    -1,    -3,   -13,   -17,     0,     2,    -5,    -3,    -3,    -5,     1,    -2,     3,     4),
		    79 => (    1,     0,     4,     0,    -2,     5,    -4,     1,     1,    -4,    -2,     1,     5,     2,     3,     3,     3,    -5,    -1,     0,     1,     0,     2,    -1,     0,     4,     2,    -2,     3,     3,    -1,     0,     3,     3,     5,     4,     5,     4,     1,    -7,    -9,    -7,     3,     2,     2,    -2,    -2,     1,    -5,     0,     3,     3,    -3,     0,     4,    -4,    -1,    -3,     2,    -3,     4,     0,    -4,    -1,    -1,    -7,    -5,    -6,    -2,    -4,   -10,    -4,    -4,    -4,    -3,    -3,     0,     2,     3,     3,     0,     0,    -1,     2,     1,    -1,    -3,     1,     4,    -3,    -3,    -5,    -9,    -5,   -12,   -22,    -5,   -13,   -18,   -15,   -17,    -2,     9,    15,   -10,    -6,   -11,    -5,    -2,     0,     4,     1,     0,     4,     3,     1,     1,    -4,   -19,    -5,    -6,   -15,   -17,    17,    12,    13,     1,   -14,   -16,   -25,   -32,   -29,   -34,   -16,   -12,     3,     1,   -18,   -11,    -4,    -4,     2,     1,    -4,     0,     1,    -3,    -8,   -32,   -40,   -26,    26,    -1,     3,    -7,    11,    35,   -11,    -5,    -6,    12,   -18,   -19,    -9,   -12,   -17,   -19,    -3,     0,   -14,    -6,     0,    -5,   -22,    -2,   -33,   -12,   -17,   -10,   -14,    10,    10,    19,    10,     5,     9,   -10,   -24,   -29,    -6,   -13,    -9,    -4,    -9,   -11,    -8,     5,    -4,    -8,     3,    -4,   -32,   -31,   -60,    22,   -37,     8,    23,    12,    10,     9,   -12,   -10,   -30,   -57,   -27,   -15,   -14,   -13,   -12,    -7,    -7,   -11,   -10,    -8,   -26,    -9,    -6,   -10,   -19,   -40,   -45,    28,    -8,    20,    24,    21,   -14,   -36,    -7,   -25,    -8,   -19,    11,    -7,   -16,    -9,   -17,   -18,   -13,   -31,     0,     0,   -17,    -9,    -5,   -25,   -23,   -57,    -9,    24,     0,    13,     2,   -29,   -27,   -20,     2,    -6,    10,   -21,     9,    -3,   -20,     5,   -12,    -9,   -22,   -14,    -6,     2,    -6,     2,     3,   -13,   -10,   -24,    15,    26,    17,   -12,     6,   -20,    10,    37,    23,     0,    18,    26,    15,   -18,   -40,   -17,   -25,   -11,   -17,    -2,   -16,    -5,   -10,     1,    -4,   -11,   -14,    -7,    -1,    17,     5,     2,     2,    20,    26,    34,    12,    22,    28,     7,     1,   -16,   -19,   -26,   -22,    -5,   -19,     1,   -14,     5,    -2,    -8,     1,    -5,   -14,   -24,   -12,    -6,    -8,    -6,     6,     0,    18,     0,     2,     8,    10,     1,     5,   -10,   -13,    -1,   -37,   -36,   -14,   -19,    -6,     2,    -6,    -6,   -21,   -13,   -12,   -24,    -5,   -10,     6,   -22,    -7,    -4,    13,    -1,    25,    19,     0,   -40,   -15,   -19,   -26,    -7,   -14,   -18,   -12,   -19,     1,    -2,    -5,   -13,   -16,   -12,   -12,   -25,   -10,   -32,    -4,   -21,   -13,    -3,    13,   -13,    -7,     7,     5,   -16,   -28,   -18,    -5,    15,    -6,    -1,   -17,    -7,    -4,     3,     4,    -5,   -13,    -3,    -9,    -7,   -50,   -43,     1,    11,    18,    17,    -5,    -4,   -20,    10,     9,   -34,   -27,   -34,     5,    12,    -9,     4,   -10,    -8,   -11,    -2,    -3,    -9,    -6,    -1,   -10,   -11,   -25,   -59,   -51,   -29,     0,    -7,   -32,   -21,   -19,    -2,   -18,   -16,   -45,   -28,    -7,     8,    -1,     6,   -13,     2,    -5,    -1,    -2,   -13,     1,     1,    11,     9,   -13,   -20,   -38,   -48,   -75,   -39,   -24,    -9,   -15,   -10,   -14,   -19,   -40,   -23,    -8,   -20,   -20,    11,    -5,    -7,    -6,    17,     4,   -12,    -7,    -8,   -17,   -12,   -15,   -20,   -23,   -33,   -63,   -26,   -14,   -10,   -23,   -10,    -5,   -22,   -34,   -47,   -20,   -22,   -31,   -15,    -2,    -5,    -9,     4,    -8,    -3,     0,    -5,   -27,   -32,    19,   -18,   -24,   -29,   -40,   -12,   -12,    -7,   -12,   -16,   -26,   -12,     0,   -36,     6,    -2,    -6,   -10,    -8,   -10,     5,     0,    -9,    -6,    -5,    -6,     6,   -22,     7,     8,   -10,     1,   -14,    -7,    -9,   -15,   -23,   -15,   -20,    -2,   -10,   -31,     0,    11,    -2,    20,     6,    -3,     1,     0,     4,   -13,    -7,    10,    15,   -30,     1,    16,    32,     9,    -3,    -7,    -7,   -27,   -21,   -25,    -4,    -2,     1,    -9,   -15,    -4,    19,    13,    14,   -16,     1,     3,    -4,   -28,   -16,     0,    -9,   -32,   -21,    16,    21,     1,    17,     2,    -1,    -4,   -14,    -2,    -5,    10,     4,    -3,   -13,   -10,     9,    26,   -21,    -4,    -4,     4,     5,    -2,   -12,    -3,   -17,   -18,   -25,     1,    16,    14,    23,    10,    10,    13,     9,    -2,    -5,    11,    -3,     7,   -22,     8,     6,    20,    -7,    -3,     3,    -3,     1,    -2,   -26,     0,     1,    -6,     0,     9,    -2,    10,    -4,   -19,   -12,    -1,    -7,     6,    -1,   -20,   -26,    13,    -1,     1,     5,    -2,    -4,    -5,    -3,     0,    -2,     8,   -10,     1,    -1,    13,    23,    -1,     6,   -15,   -17,   -18,   -20,    -7,     1,     4,    20,   -22,   -29,    15,     4,    13,    13,    -1,    -3,     2,    -1,     1,     5,    -2,    11,     5,    -2,    -8,     3,   -39,    -3,    21,     8,    -3,    -3,    30,   -10,   -31,   -24,   -14,   -18,    -4,     2,    -6,     7,     8,    -2,    -4,    -3,    -1,     4,     4,    -4,    -8,    -6,     3,     5,    -8,   -11,    -5,    14,     2,    -9,     1,    14,    26,   -16,     2,     0,     2,    -6,    -3,     1,    -4,     4,     3,    -3),
		    80 => (    0,     5,    -5,     5,    -2,     2,     1,    -4,    -3,    -4,    -1,     2,    -4,     4,     2,     5,    -4,    -5,     5,     4,     0,     5,    -2,     0,    -1,    -4,    -5,     2,    -3,     4,     3,    -2,     5,     4,    -2,     5,    -2,    -4,    -4,     3,     3,     6,    -8,    -3,     3,     2,    -6,    -1,     1,     1,     0,     0,    -1,    -3,    -3,     0,    -4,     1,    -5,    30,    28,     0,     4,     6,    -5,    -8,    -3,   -22,   -18,   -31,   -34,   -31,   -19,   -22,   -18,   -22,   -17,   -18,   -21,   -13,   -17,    -8,    -1,    -3,    -3,    -1,     4,    37,    22,    11,    -6,    -9,   -15,   -13,   -14,    -8,   -11,    14,     4,   -10,     3,    -6,    -8,    -2,     5,   -34,   -24,   -21,    -1,    -6,   -17,    -4,    -1,     2,    -3,    -1,    -8,   -11,   -15,   -17,   -15,    -9,   -10,   -13,   -23,   -11,    -6,     5,   -13,     3,    18,     6,    18,    11,    34,   -10,    -1,   -12,   -20,    -3,     0,     3,    -7,     6,     3,     2,     7,   -29,   -35,   -29,   -32,   -45,   -25,     0,    -5,    -5,   -10,    10,    11,     9,    23,    14,    36,    -6,    -2,   -14,   -18,    -9,    -4,     3,    -7,    -5,     5,    24,     3,     4,   -25,   -45,   -38,   -41,    -7,    19,     0,     6,   -27,   -11,     1,     3,    -4,    27,    19,   -19,   -33,   -40,   -22,     0,    -3,    -2,    -4,    -8,    14,    28,     5,    -9,   -16,   -10,   -15,     5,     1,     2,   -17,    -4,    -9,    -7,    -1,    15,     8,   -16,    13,    10,    -6,    -9,   -29,     9,    11,    -9,    11,   -10,     3,    17,    12,   -12,   -14,   -21,   -32,   -29,   -12,   -11,    18,   -14,     8,    -5,     9,     6,     4,    17,    16,    11,   -21,   -28,   -30,    -6,    -2,    -3,    14,    -3,   -13,    16,   -10,   -17,    -8,   -40,   -13,   -26,    -9,    -5,    17,    10,   -18,    -4,     7,     0,     9,    -5,     8,    21,    17,     6,   -21,     2,     2,    -1,     8,    -1,   -20,    -8,   -33,   -13,   -16,     5,   -15,    -5,    16,    -2,     4,    12,     1,   -18,   -30,   -12,    25,    17,    22,    19,    18,     7,   -37,    -4,    -4,    14,   -11,   -10,   -24,   -24,   -18,    15,     4,    -5,   -10,     3,     3,   -13,    -6,   -17,   -38,   -46,   -44,     0,     8,     9,     1,    -2,    -6,    -1,   -20,    -3,     5,    13,    -5,    -6,   -10,   -17,   -17,    -3,    -4,    -6,    13,    15,    15,    17,     9,    -9,   -66,   -60,   -14,    12,   -20,    -5,     9,    32,    -3,    -8,   -17,     0,     4,    11,     9,   -17,   -13,   -11,     1,     5,     6,    11,     3,    14,     9,    11,     2,   -18,   -79,   -30,    15,    -2,   -17,   -21,     2,    63,    18,    14,   -16,    -4,     1,    -2,    -1,   -42,   -11,    -6,     8,    21,     0,     7,   -18,    -1,    -5,    -9,   -66,   -56,   -60,   -25,   -14,   -12,   -11,     6,     4,    27,     9,    -7,   -29,    -1,     1,     3,    -9,   -45,     7,   -15,     2,    23,     7,     8,   -26,   -10,    15,    -2,   -47,   -31,   -10,    -1,   -16,   -10,   -33,     4,     6,    17,    29,   -19,   -33,    -9,     5,     3,    -1,   -32,     8,    -1,    -1,    21,    14,   -12,   -12,     2,   -19,   -31,   -12,    -4,     2,    -9,     6,   -18,    -8,   -18,    -7,     2,    17,   -26,   -14,     2,     0,    -5,   -14,   -16,     6,    20,     9,    22,   -10,     7,    -1,   -14,   -43,   -30,   -18,    -5,   -14,    -1,    -3,     8,     8,   -22,   -15,     5,    15,   -29,   -15,     2,    -5,     2,   -10,    -2,     9,     3,     7,    19,    27,    12,   -23,   -43,   -34,   -14,     1,     3,    -5,    -1,     8,   -16,    -3,    -7,     8,     4,     3,   -13,    -8,    -6,     5,     6,   -27,    -9,    31,    -1,     2,    14,     7,    13,   -21,   -40,   -17,   -21,    -1,     6,   -16,     4,   -13,    -8,   -24,    -7,     8,    -1,    11,   -18,    -3,     4,     1,     7,   -38,     9,    27,     6,    13,    -4,    10,     9,    -4,     7,    -8,   -10,    -5,   -27,    -6,    -7,    -7,   -26,   -29,   -10,     3,    -4,     4,   -16,     5,     5,     2,     5,   -37,    10,     5,     4,    15,    22,     5,    10,     1,    -1,   -13,    -9,     2,    11,     0,    -4,   -20,   -25,   -35,   -37,   -22,    -6,    19,   -10,     4,     7,     2,    -4,   -42,     0,    -1,    19,    23,    10,     9,     7,     9,   -12,   -15,     3,    15,     1,   -35,   -28,   -12,   -15,   -42,   -25,    -5,    -3,    16,     2,     1,     5,     4,     0,    -7,   -30,   -33,     5,     3,     1,     4,    14,    17,    15,     2,    11,    12,   -21,   -33,   -21,   -31,   -28,   -40,   -18,     7,     1,   -23,     0,    -3,    -4,     0,    -2,    -9,    -7,    29,    37,    -2,    -9,     3,    20,    33,    22,    30,   -32,   -28,   -29,   -57,   -49,   -28,   -30,   -14,     4,    -4,    -1,    12,     3,    -2,    -4,     3,    -5,     0,     0,   -20,   -38,   -35,   -35,   -30,   -19,   -25,   -31,   -41,   -30,   -12,   -33,   -35,   -32,   -39,   -28,    -2,    -7,    -6,    -6,    -1,     0,    -4,     2,     5,     3,    -3,    -5,    -4,   -28,   -38,    -9,    -1,   -10,   -16,   -19,   -10,   -14,   -11,   -20,   -22,   -36,   -38,    -8,   -23,   -10,   -10,    -5,     0,     2,    -4,     3,    -4,    -5,     5,     4,     1,     3,     4,    -4,    -1,    -1,     1,     3,     3,    -2,     1,    -1,    -2,     2,    -1,    -6,    -4,    -6,    -7,    -5,     1,     0,     4,    -4),
		    81 => (   -4,     2,     4,     5,    -3,    -3,     1,    -4,    -4,     3,    -2,     5,     1,    -2,     5,    -1,     2,    -1,     3,    -1,     3,    -1,     4,    -1,    -5,     4,    -3,     4,    -2,     1,     3,     0,     0,    -4,     1,    -1,     1,     5,     0,    -3,    -1,    -8,     5,     6,    -3,    -7,     1,    -4,    -2,    -1,    -3,     2,     3,    -1,     2,    -3,    -3,     3,    -3,     5,    -1,     4,    -1,    -5,    -6,    -5,    -6,    -4,     0,     1,    25,    31,    66,    49,    24,   -16,     4,   -22,   -16,   -13,    -2,     4,     4,    -2,    -1,     0,    11,     9,    -5,   -17,   -35,   -12,    22,     7,   -14,   -25,   -21,    -5,    10,    37,    41,     8,     1,   -18,     1,    23,    -5,    -1,   -17,    -1,     2,    -2,     3,     5,    13,    11,    24,    10,    -7,    -9,    35,    26,    16,    -3,    -3,   -15,    -3,     9,    12,     6,    -8,    -8,    17,    23,    11,    17,    -3,   -13,   -12,   -16,    -1,    -5,    -3,    -4,    27,    52,    23,    20,    14,     5,     4,   -26,   -27,     5,    17,     4,    -9,     5,     2,     9,    17,    18,    16,     5,     3,    -6,   -14,   -14,     3,     2,   -33,     2,     4,    11,    23,     7,   -15,   -19,    10,    -6,     0,    -4,    -3,    -5,   -20,    14,     7,    24,    14,    -4,     6,    -2,    -2,    -3,    -8,    -3,    -5,     3,   -38,   -33,   -33,    -2,    13,    15,   -25,     5,    17,   -15,    -3,   -21,    -5,    14,    -4,     5,    13,    27,     4,    -3,     9,    -8,    -8,     1,   -16,    -8,    -1,    -3,   -42,   -26,   -31,    -6,     6,     1,    -7,    12,     7,     5,    11,   -20,   -22,     4,    15,     2,    16,   -22,   -13,   -10,     5,   -13,    -1,    -1,   -16,    -3,     2,    -2,   -41,   -17,   -20,   -22,     1,    11,    18,     2,     4,    31,    24,   -15,   -27,    -8,   -14,   -15,   -15,   -11,    -9,   -11,   -15,     0,    -6,     3,     3,    -5,     1,    -2,   -32,    -5,   -36,   -18,   -32,     3,    14,    21,     9,    34,     9,    -9,   -14,    -9,   -21,   -17,    -6,   -30,   -19,   -22,    -2,    -3,    -6,    -4,     6,     1,    -1,     7,    -7,    -3,   -30,   -16,   -28,     1,   -14,     9,     2,    18,     7,    -7,    -4,   -21,     2,   -22,   -20,   -27,   -17,   -13,     3,     0,    -4,    -4,    -3,     5,    -2,    -2,    -4,   -11,   -21,   -21,     9,    18,     4,     2,    -9,     3,    -2,   -17,   -21,    -6,    -7,   -23,    -9,   -27,   -40,   -18,    -9,    -9,    -5,    -6,     3,     9,     0,    -1,    -6,    -5,   -28,    11,    18,    19,    26,   -11,   -15,    -1,    -6,   -22,    -9,    13,    -7,   -16,   -18,   -58,   -27,   -23,   -19,   -16,   -14,    -2,    -2,    -1,    -2,     0,     3,    -1,   -24,    21,    18,    -4,    -8,   -33,   -43,   -25,   -15,   -13,     7,     9,    -1,   -14,   -24,   -38,   -34,   -39,   -26,   -17,   -10,   -15,     1,     3,    -4,     3,    -2,     7,    -5,   -20,   -12,   -12,   -22,   -29,   -37,   -38,   -44,    -3,    19,     4,    -5,   -16,   -22,   -50,   -29,   -30,   -24,   -25,   -58,    -8,    -3,    -7,     3,    -2,     7,   -12,   -11,   -11,   -17,   -17,   -38,   -21,   -23,   -40,   -35,    -3,    25,    19,    -6,   -22,   -18,   -39,   -34,   -41,   -15,   -28,   -19,    -7,    -5,    -8,    -2,    -2,    -2,   -21,    -5,    -9,   -16,   -29,   -30,   -28,   -32,   -69,   -38,   -31,    11,   -11,   -10,   -12,     2,   -15,   -20,   -15,     0,   -17,   -30,   -32,    -3,   -12,    -6,     3,     3,    -6,    -6,   -25,   -49,   -28,   -48,   -32,   -35,   -88,   -77,   -43,     0,   -15,    -7,     6,    -8,    -7,    17,    11,    25,   -12,   -58,   -13,   -13,   -10,    -2,     0,    -6,   -11,   -17,   -45,   -26,    -6,    -2,   -18,   -24,   -42,   -27,   -21,   -15,    11,    21,     3,   -18,    -1,     9,     0,    -2,    11,    -3,    -2,   -20,    -6,     3,    -5,   -13,    17,    -1,   -34,   -14,     6,     7,    15,    29,     4,    -7,     2,    11,    10,    27,    17,    40,    30,    25,    -1,    10,    12,     6,     4,   -15,     3,    11,     5,   -17,    18,    21,     8,    23,    20,    25,    25,    14,    14,    -2,     9,    10,    22,     6,    23,    37,    11,    14,    -3,   -18,   -10,     8,    16,   -19,     4,    11,     2,   -47,   -29,    14,    35,    11,     3,     6,    10,    10,     8,     5,     9,    -3,     8,    -9,     9,     5,    21,    22,    11,   -37,   -24,     5,    -3,    -2,     1,     5,     2,    -5,   -14,     7,    -7,    12,    -6,    -3,    -9,   -13,     2,     2,    15,   -17,   -28,   -37,   -30,   -10,     6,    17,    21,    -8,   -20,   -20,   -25,    12,     3,     0,     0,    -4,     1,    -9,   -14,   -20,    -4,     6,    12,    -6,    -4,   -35,   -23,   -45,   -38,   -34,   -21,   -13,    -4,     5,     9,   -12,   -16,   -22,    -4,     0,     4,     0,    -2,     5,    -6,    -2,    -3,   -10,    -4,    -3,   -22,   -10,   -14,   -20,   -23,   -15,   -30,   -22,   -26,   -31,   -26,   -31,   -25,   -20,    -9,     0,     2,     1,    -4,    -4,     5,    -3,     1,    -7,    -8,   -10,    -8,    -6,   -21,     1,    -4,   -11,   -17,   -11,   -21,    -5,   -22,   -13,   -18,   -13,   -11,    -7,     2,    -4,    -3,     3,    -2,     2,    -3,    -2,    -4,     0,     5,     1,    -1,    -1,    -3,    -8,    -8,    -1,    -6,    -5,    -6,    -6,    -5,    -4,    -1,     0,     0,    -2,     0,     2,     3,    -2,     5),
		    82 => (    1,     1,    -4,    -3,     0,    -2,     2,    -5,     5,     0,     0,     1,    -5,    -1,     6,     5,    -1,     1,    -3,     3,    -2,    -5,     4,    -2,    -5,     2,    -1,    -1,     0,     4,     5,    -1,    -4,     5,     3,   -12,   -19,    -8,   -17,   -16,   -19,   -34,   -14,     2,    17,     2,   -19,   -37,   -24,   -13,   -18,    -6,    -1,    -3,    -1,     1,     3,     5,     0,   -26,   -28,     4,    -1,    -5,     0,    31,    27,    12,     7,     9,     4,    12,    -1,    -3,   -14,   -24,   -15,   -11,    -9,    -1,     4,     6,     0,     1,    -1,    -3,    -2,   -29,   -37,    -5,    -1,    10,   -11,    13,     6,     5,    -9,    10,    21,    11,    11,     3,   -13,   -16,   -11,     4,   -20,   -47,     5,     7,     2,     1,     0,     3,    -8,     8,     7,   -12,     3,    -5,   -25,    12,    25,     4,     4,    15,    19,     6,    11,     6,    26,     3,    -1,    -9,   -23,   -11,   -15,    -5,   -11,    -1,     0,    -4,     7,    -2,    -3,     7,     7,   -24,    -2,     6,   -16,   -11,     6,     0,     0,    -5,    17,    -7,     4,   -12,    -8,    -7,   -15,    -8,   -32,    -1,   -13,   -11,    -2,     2,     3,   -12,   -12,     2,     1,    19,   -16,   -14,     5,    -9,   -22,    20,    -1,     6,    23,     3,     7,   -19,   -11,    -2,   -12,   -17,   -40,    16,    -8,    -5,    -4,     2,    -4,   -11,   -12,    -5,    11,     0,   -16,   -14,    14,     4,    -1,   -16,     1,    11,    -1,     3,   -27,    -6,    11,    18,    -4,   -40,   -15,     5,   -20,    -9,    -8,     7,    -8,   -17,   -10,   -25,   -15,     1,    10,     8,    20,    11,   -23,   -14,   -28,    -2,     0,     5,     9,    19,     1,     3,     2,   -19,   -33,   -40,   -15,    -6,    -1,    -8,    -4,   -14,    -9,   -33,   -28,   -36,   -43,   -11,     1,   -23,   -34,    -2,    -4,   -20,    -5,     7,    14,   -14,    -6,    22,    -1,   -18,   -18,   -21,   -14,   -12,    -4,     2,    -4,   -23,   -23,   -32,   -36,   -69,   -98,   -88,   -71,   -58,   -18,   -21,    -4,   -23,     2,    -9,    10,     2,    -2,    -8,    -2,    -9,   -30,   -24,   -11,    -5,    -1,   -13,   -13,   -27,   -26,   -33,   -49,   -59,   -79,   -67,   -56,   -31,   -23,   -33,    -7,   -22,   -15,   -35,   -34,     1,    -1,     3,    11,    -9,   -30,    -3,   -12,    -9,     5,   -16,   -33,   -25,   -42,   -30,   -28,   -37,   -10,    -9,    -5,     6,    -4,    -6,     4,   -15,   -26,   -31,   -23,   -12,    -7,    10,    22,   -24,   -25,    29,     3,    -7,    -5,   -14,     2,    -9,   -20,   -14,     5,    38,    16,    -4,   -10,     7,    36,    25,    10,     6,    -1,     1,   -13,   -17,    -3,    13,    29,    -2,    -5,    12,    -2,    -1,     0,   -15,   -21,    25,    16,    -3,    25,    38,    31,    22,    31,    24,    20,    32,    29,    -4,    15,   -27,   -14,    -5,    11,    -2,     6,     5,    -6,    17,    15,    14,     0,    -9,     5,    58,    25,    31,    19,    17,    15,    16,    27,     9,    15,     8,   -13,    10,    -5,     5,   -11,    -1,   -14,    -9,    -6,    16,    -3,    24,    45,    27,    -1,     1,     5,    24,    -9,    30,    46,    22,    10,    14,    18,     3,   -17,    10,    11,     9,     7,     8,    -3,     1,   -14,   -17,   -10,    -7,   -20,    33,    44,    18,     3,    -7,     3,   -13,    13,     9,    31,    -8,    14,   -11,   -16,     7,     0,    -6,    22,    15,    15,     2,    -1,   -15,    -3,   -34,   -24,   -28,   -36,     5,    10,    29,     3,    -4,   -18,     6,    -2,    23,    24,     0,     0,   -10,   -16,    -8,    -1,     6,    -5,    -1,    16,     4,    14,    21,    11,    -9,   -16,   -14,     6,    23,    13,    28,     2,   -17,   -17,    -7,    14,    13,    17,    14,     8,     4,   -13,     3,     1,    -6,   -15,    -3,     5,    -1,    17,    20,     3,    17,    18,     7,    27,    25,    20,    14,    -3,   -20,     2,    -2,    10,    31,    10,     2,    -5,   -18,   -11,   -20,   -27,   -23,   -23,    -4,    -1,   -19,   -13,    -3,    -6,     0,    -8,     6,    30,    -4,     9,    -1,    -5,    13,     0,     8,    13,     9,     8,     8,    13,   -16,   -19,    -5,    -6,   -24,   -17,   -16,   -18,    -6,   -16,    -1,    12,    20,     8,    17,     9,   -17,   -11,    -2,    -4,    -3,    -2,     6,    15,   -15,   -14,    -6,    -5,   -15,    -5,     4,    -9,   -22,   -29,   -10,   -18,   -21,   -27,    -5,     2,     5,    -7,    -9,   -12,   -29,   -32,    -4,    -4,    -5,     7,    25,    23,     4,   -25,    -6,   -16,   -30,    -9,   -18,    -2,   -37,   -20,   -34,   -13,   -17,   -22,   -39,   -18,    -1,    15,   -24,   -22,   -17,   -21,     3,     2,     4,   -13,    -9,   -10,    -4,    -9,   -20,   -23,   -40,   -46,   -34,   -27,   -44,   -34,   -29,   -28,   -12,   -18,   -39,   -47,   -27,   -43,   -26,     7,    13,    13,     1,     0,     1,    -7,     1,   -10,    -8,    -6,   -14,   -27,   -35,   -12,    -8,   -12,   -32,   -25,   -16,   -24,   -30,   -19,   -40,   -30,   -18,   -23,    -8,    -9,     8,    17,     0,     2,     3,    -2,     2,    -9,   -13,   -12,    -9,   -11,    -4,    -4,    -3,     0,    -1,   -13,    -7,   -32,   -24,   -20,   -14,    -8,    -7,    -4,   -10,     4,     0,    -2,     0,     4,     5,     0,    -1,    -3,     0,     1,    -4,     1,     4,    -9,    -4,    -4,    -9,    -2,    -3,    -3,     0,    -6,    -7,   -12,   -15,    -9,    -4,    -1,    -1,    -3,    -4),
		    83 => (    5,     1,     2,     3,    -2,    -2,    -4,    -4,    -3,     0,    -2,    -4,    -1,    -1,    -7,    -7,    -2,    -2,     3,     0,     4,     0,     3,     5,     2,    -4,     3,     4,     0,     2,     1,    -3,     3,    -4,     1,    -4,    -5,    -1,    -8,    -6,    -7,   -22,   -17,   -16,    -8,   -25,   -12,   -13,    -7,    -5,    -5,    -1,     5,     3,    -4,    -5,    -1,     2,    -1,    -1,   -11,   -10,   -12,   -13,   -25,   -32,    12,    -2,   -11,   -19,   -26,   -25,   -18,    -3,     3,   -22,   -30,   -39,   -36,   -30,    -5,     5,    -4,     1,    -3,     4,    -6,    -6,    -5,    11,    21,    57,    54,    21,    24,    23,    17,     7,    -4,    27,    36,    23,    20,    47,    83,     8,   -52,   -54,   -27,   -15,     1,     1,     4,    -2,   -33,     2,    11,    17,     6,    34,    44,     0,    24,    11,    13,    -4,    10,     1,    15,    25,    20,    21,     9,   -28,   -28,  -105,   -81,   -30,   -21,     2,     1,     4,    -5,    -3,    -3,    17,    39,    49,     5,    12,    19,    -9,   -16,     3,   -10,    -3,    23,   -12,    -5,    14,     4,    -6,    -8,     7,     8,   -40,   -18,     2,     3,     6,    11,    -2,    -5,    34,    53,    44,    21,    22,    10,     2,   -14,     7,    -2,    15,    12,     5,     5,    -3,     2,    -7,    -1,     5,    17,   -46,   -22,    -8,    -2,     3,     1,    10,    -5,     7,    49,    64,    33,     2,     4,    30,     4,   -17,     5,    -1,    12,    -9,   -16,     9,    -8,    -9,   -14,    -6,    14,   -42,   -26,   -12,   -15,    -5,   -19,    -2,     9,    35,     6,    17,     4,    -8,    -6,   -23,   -28,   -17,    -7,    26,    13,    16,   -20,    14,     4,   -18,    12,     2,   -13,   -27,   -25,    -2,     0,   -11,   -49,   -11,    51,    49,    21,    22,    25,   -12,    10,   -16,   -13,    -8,   -13,   -12,     3,    28,    13,    -5,     9,   -11,    29,    23,   -57,   -24,   -18,     3,    -5,    -2,   -53,     3,    11,    25,    30,    39,     0,   -11,   -25,   -30,   -16,   -26,    -8,   -14,    -2,    17,    20,     8,   -22,   -17,    10,    37,   -26,   -27,   -21,     0,    -4,   -19,   -24,    28,    43,    41,    25,    10,    19,   -10,    -4,   -23,   -24,    -7,    -2,   -22,     4,     5,    11,   -20,   -26,   -13,     2,   -11,   -68,   -48,   -23,    -5,    -5,    -6,   -25,    11,    28,    41,    29,    15,     4,   -17,     8,   -10,   -14,   -15,   -17,     4,     5,    -2,     4,     9,   -14,   -31,   -13,     2,   -43,   -30,   -10,    -3,     4,    -7,   -22,     2,    44,    31,    19,    15,    34,    -3,    13,   -11,   -15,    -5,    -9,    18,   -47,   -13,    21,    18,   -16,   -17,   -22,    13,    -8,   -47,   -11,    -4,    -1,    12,    -5,    10,    19,    32,    32,    -4,    14,     1,   -10,    -6,     0,   -13,     9,   -22,   -22,    -6,    13,    14,     9,     6,    -9,    13,    -8,   -65,   -29,     4,    -6,    13,   -11,     6,    15,    41,    25,   -23,   -12,   -26,    -2,   -18,    -8,   -18,   -15,    -8,   -22,   -24,    -8,    26,     3,     8,    15,    29,    33,   -67,    12,   -13,     4,     1,     6,    43,    40,    34,     5,    13,   -30,     1,     3,   -24,   -40,    -7,     4,   -10,   -24,   -18,    21,    32,     5,   -13,    15,     3,    22,   -75,   -32,   -17,     0,     7,    -9,    21,    26,     7,    -9,     5,   -11,    -7,   -18,   -18,     1,     0,   -24,   -15,     7,     7,    15,    30,    -5,     3,   -15,   -11,   -15,   -60,   -18,    -9,   -10,     7,    -3,    13,    34,    24,     0,    -2,    -9,   -24,     0,    -8,   -19,    19,     0,    18,    -2,    12,    30,   -15,    10,   -12,    -8,   -37,   -11,   -59,    -3,   -16,    -3,    -9,    10,     7,    13,    22,   -12,   -16,   -21,   -36,   -18,   -21,    -4,     6,    22,    20,     2,    19,    16,    -8,     9,    -5,    -9,   -14,     9,   -30,   -24,   -18,    -2,     8,   -25,     6,    12,    15,     0,    -7,   -22,    -1,   -18,   -15,    -7,     1,    20,    14,    38,    26,    -5,    -7,    17,    14,    16,    17,    -2,   -42,   -19,    -2,    -5,    -6,    10,    -2,     5,   -21,    16,    28,    -1,    -8,   -14,     0,     9,    18,    29,    31,    21,     9,    13,    28,    -2,    14,    23,    -7,   -33,   -41,   -22,    -4,    -5,     0,    22,    16,   -22,    13,    28,    32,    -6,     6,    16,     8,   -10,     6,    18,     9,   -14,    11,    -7,    21,     3,    19,    43,     9,   -26,   -29,   -17,    -4,     4,     4,     9,     2,   -12,    -7,    12,    28,    10,     8,     5,    14,    -2,    -9,    -8,    14,    10,    -3,   -11,   -18,     2,    43,    41,    20,    36,    15,   -23,     4,     2,     1,    24,    41,    36,     0,    27,    25,    18,    31,    11,   -10,    -9,     4,    11,    -9,    -2,     3,   -18,     9,    56,    35,    20,    23,   -36,   -21,    -7,    -1,     4,     0,     6,   -12,     1,    34,    27,    -5,    11,    12,   -15,    -7,    11,    35,     3,    -5,    -5,     6,    16,    18,   -15,   -43,   -50,   -48,   -38,   -11,    -8,    -5,     0,     4,     0,    -6,   -48,    22,    11,     3,    15,   -11,    -9,   -22,   -22,   -12,   -17,     1,    43,    47,    43,     8,   -10,   -18,   -52,   -25,    -3,    -3,     2,     4,    -1,    -3,     3,     2,    -8,   -15,   -14,    -7,   -11,   -31,   -27,   -22,   -18,   -30,   -26,   -17,    -2,    -7,    -2,   -22,   -28,    -8,    -9,    -6,     4,     3,     3,     2),
		    84 => (    0,    -1,     5,     3,     2,     1,     2,     2,     4,     0,     1,     0,   -16,    -9,    -6,    -8,     0,     1,     2,    -4,     3,     0,     2,    -1,    -2,     3,    -1,    -3,     2,    -3,     2,    -2,    -3,   -10,   -16,   -22,   -13,   -21,   -19,   -18,   -23,   -26,    -6,   -23,   -21,    -4,   -12,   -12,   -22,   -14,    -9,   -19,     0,     2,     3,    -4,     4,     3,   -11,   -18,   -25,   -30,   -27,   -28,   -45,   -39,   -55,   -60,     6,    12,    -1,   -30,   -27,   -35,   -52,   -29,   -58,   -27,   -28,   -19,   -10,   -13,     5,     2,     4,    -1,    -3,   -54,   -35,   -38,   -21,   -32,   -25,   -49,   -43,   -45,   -27,   -59,    -7,    -4,   -30,   -18,   -16,    -3,    21,     0,   -27,   -31,   -18,   -11,    -5,     0,     2,     5,   -23,   -52,    -5,     0,    11,     1,   -25,     2,    -7,   -36,    -4,    -7,   -17,   -22,   -11,    -3,    -6,     3,     0,   -16,     6,     8,    12,    -9,   -34,    -6,    -5,    -5,   -27,    -4,     1,    -7,    -2,    -6,    13,    -8,    19,     1,    22,   -17,   -10,   -25,   -17,    14,    -4,     3,   -23,    -9,     4,    -2,   -12,    12,   -14,    -2,    -2,     3,   -14,   -21,    10,    26,    17,   -23,    -8,   -27,    -3,     8,    -2,   -17,   -40,   -41,   -32,   -23,   -33,   -19,   -41,    -2,    -3,    -3,    -9,    -4,    -1,   -17,     4,   -47,   -18,     1,    12,    20,   -20,   -25,   -37,   -17,    -8,    -3,   -27,   -22,   -29,   -36,   -31,   -10,   -18,   -23,   -21,   -15,   -17,   -12,     6,    24,    21,   -30,   -16,   -41,    28,     8,    21,     8,   -35,   -38,   -41,   -17,   -35,   -23,   -17,    -4,   -49,   -28,   -28,    -7,   -11,    -6,   -20,   -23,   -15,    -4,    19,    22,     0,   -10,    -1,   -32,    23,     6,   -18,    -1,   -25,   -16,   -21,   -22,   -33,    -9,     1,   -12,   -28,   -11,   -17,    -7,     1,    13,    10,    23,    12,    16,    25,   -18,   -30,   -10,     5,   -20,    16,     4,   -13,    15,   -10,   -25,   -12,    -2,    -1,     1,    18,    -7,   -14,    20,    16,    32,    -8,     2,    14,    10,     8,    -2,    -4,     5,   -16,    -7,    -3,   -24,    -4,     0,     1,    29,     0,     2,     9,    31,    24,    15,    30,    -8,     3,    20,    32,     7,   -13,    -6,     0,     5,    14,    13,    -5,    -6,   -34,   -30,    -1,    -2,    14,    16,    -5,    22,    17,    13,    19,    24,    23,    22,    28,    11,    -9,    -3,     3,    -5,   -16,    -3,    -5,    12,    23,    12,    34,    20,    17,   -35,     3,    -5,    -3,    29,    13,    25,    10,    19,     1,    13,    15,    37,    33,    19,     1,   -10,    16,    11,   -20,     4,     5,    23,    17,    22,    18,    46,    42,   -20,     3,     6,   -44,    12,    42,    29,    14,    12,    25,    17,    14,    11,    22,     0,    -7,   -13,    18,    31,   -17,    25,   -12,    29,    15,   -13,    -1,    27,    27,    -5,    -2,     8,    44,    21,    -1,    24,     8,   -11,     6,    12,    15,    12,     7,     5,    -5,    17,    27,     5,    -1,    22,    -3,    -2,    27,    16,   -11,    18,    51,    -7,     0,     2,   -10,    28,     9,    21,    28,    21,    15,     6,    -2,    -8,     9,     1,    -6,    31,    10,    14,    29,    39,    11,     6,     0,     1,    -3,    16,    32,   -12,    -4,    -8,    13,   -11,    35,    26,    11,    16,     2,     4,     2,    -1,     2,    10,     9,    10,    15,     4,     3,    18,   -14,     0,     7,     7,     7,     5,    20,    -2,   -28,     0,    26,    12,    27,    -1,    -6,    -7,     9,    18,     2,    14,     4,    20,    23,     3,     4,     6,    11,   -10,    -8,     1,    -5,   -15,    -8,   -29,    -9,   -11,     2,   -19,   -14,    37,    -2,    28,     4,   -23,    12,     4,   -14,     3,     2,    -9,    18,     2,   -11,   -13,   -17,   -31,   -22,   -18,   -33,   -36,    -9,   -22,   -11,   -10,    -1,    -5,   -25,    25,    14,    -1,     2,     1,     6,   -20,   -47,   -26,   -34,   -16,    -7,   -21,   -10,   -25,   -31,   -26,   -46,   -35,   -26,   -33,   -11,   -51,    -9,     0,    -2,    -8,   -40,    12,    16,     6,   -22,   -37,   -12,   -22,   -32,   -19,   -27,   -20,   -32,   -14,    -1,   -12,   -20,   -33,   -12,   -27,   -14,   -22,     6,   -31,   -34,    -2,    -5,     0,     0,   -29,   -46,    -8,     0,   -36,   -39,   -35,    -7,   -10,   -25,   -27,   -16,    -9,   -18,   -22,   -18,    -7,   -24,     6,     4,    15,   -16,   -11,    -6,    -9,    -4,    -1,    -2,   -39,   -19,   -47,     0,    12,     3,   -28,    13,   -14,   -10,   -12,   -15,   -10,   -13,     1,   -15,    -5,   -14,     6,   -10,   -25,   -34,     3,    -2,     4,    -2,     1,     0,    -5,   -36,    -3,    10,    16,    14,     9,   -18,    -6,   -32,    11,    17,   -16,    -1,   -18,   -40,   -26,    -5,    12,    -6,   -19,   -57,    -9,   -14,     2,     1,    -3,   -11,    -7,     7,   -27,     7,     0,   -12,   -26,    -9,   -10,   -34,   -28,   -13,   -42,    -6,   -15,   -20,   -32,    -9,    -2,    14,    -5,   -36,   -17,   -12,    -1,     2,     4,    -1,   -30,   -14,    -8,   -30,   -35,   -15,   -16,   -50,   -36,   -25,   -52,   -47,   -34,   -46,   -18,   -11,   -50,   -68,   -65,   -58,   -16,   -15,    -5,    -4,    -3,     4,     1,     4,    -3,    -3,    -7,    -6,    -7,   -11,   -12,   -39,   -43,   -23,   -32,   -41,   -13,   -22,   -45,   -28,   -31,   -38,   -29,   -26,    -7,     3,    -3,     2,    -4),
		    85 => (    1,    -1,     4,    -5,     0,     0,     1,    -5,    -1,    -4,    -4,    -4,    -3,    -7,    -1,     3,     3,    -3,     2,     0,    -3,    -4,     1,     2,     5,    -1,    -4,    -4,    -3,     5,    -1,    -3,    -5,    -3,    -4,     4,     1,     4,    -8,   -19,   -17,   -21,   -15,   -14,   -21,   -19,   -25,   -31,   -17,   -16,    -7,    -4,    -5,     1,    -2,    -1,     1,     5,    -9,    -9,    -7,    -6,   -14,    -9,   -48,   -37,   -56,   -50,   -39,   -40,   -41,    -7,    -5,     8,    10,   -10,    11,     5,    -5,    11,   -18,    -9,     3,     3,     1,     3,   -15,    17,    24,   -15,   -53,   -42,    -8,     5,    16,   -28,   -34,    -6,   -18,    28,    20,    10,    39,    30,    33,    64,    51,    36,   -15,    16,    12,     0,    -2,    -1,   -18,    18,   -55,   -48,   -27,   -16,   -53,   -15,    17,   -14,   -13,   -25,     7,    25,    24,    39,    73,    34,    37,    44,    77,    36,   -25,     5,   -17,   -13,     2,     4,   -25,    25,   -59,   -20,   -17,   -15,     0,    18,    22,     3,   -16,   -26,    10,    10,    26,    35,    43,    46,    57,    11,    36,    11,   -14,   -18,   -26,   -29,     2,     2,    -6,   -56,    -9,    29,    28,    12,    25,    12,    11,     0,     1,   -25,    -3,     2,     6,    -2,    32,    51,    32,     1,    27,    23,    38,    37,     6,     7,    -2,    -8,    -4,   -62,   -34,   -14,    14,     6,     3,     0,     1,    22,   -19,   -10,   -12,   -38,    -9,   -13,    23,    39,    13,    18,    60,    49,    45,    11,    20,    36,   -16,   -19,   -26,   -66,   -20,   -24,    10,    16,    -5,    -1,   -22,     9,    15,    -1,   -14,   -28,   -38,    -6,   -12,    37,    27,    27,    51,    44,    28,     5,    15,    22,     3,     0,   -27,   -35,   -17,   -15,    -9,    10,     6,   -15,     5,     3,    -4,    -2,   -23,   -39,   -38,   -29,    -7,    32,     3,     9,    26,    35,    36,    18,     3,    -1,    -3,    -6,   -18,   -56,    11,    -1,   -23,   -25,     1,    14,   -23,    18,    16,   -14,   -23,   -17,   -44,   -36,    11,     5,     6,    27,    25,    39,    47,     9,   -13,   -14,    -3,    -5,     1,   -40,     9,   -19,     1,   -19,     6,    -8,   -11,    -2,     5,   -12,   -30,   -16,    17,     9,    -1,     4,   -21,    -7,    19,    34,    43,    28,   -15,   -11,     1,     0,    -7,   -30,    35,    -6,    -7,    15,    12,    19,    38,     3,    29,    -8,    -8,   -24,    -6,   -11,    -6,   -23,   -25,   -20,     1,     9,    11,    34,    50,   -16,     4,    -3,    -4,   -35,     3,     5,    -7,    24,     0,    -1,    13,    17,    22,    -7,   -18,    -5,    -8,   -19,   -29,     7,    -9,    19,   -22,   -31,   -32,   -21,    36,   -16,     1,     1,   -11,   -38,    21,    10,    31,    -4,     0,    19,    19,    17,   -10,     3,     7,    -3,    -1,   -12,     6,    -2,    19,    -6,    15,     0,    -7,   -38,   -39,   -16,     8,    -2,   -23,    -7,    27,    37,     3,    16,    -7,     8,    15,    -4,    -6,     2,    -7,   -37,   -12,     5,    -7,    -5,   -10,    -6,     3,    12,     9,   -17,   -31,    -9,     0,    -5,   -27,    -9,    10,    33,    42,    15,     5,     7,   -11,   -13,   -20,     1,    -9,   -20,   -32,     2,    20,     5,   -14,    16,    23,    -2,   -24,   -50,   -44,   -13,     1,    -7,   -34,    -6,    23,    43,    16,    53,    29,     1,    -3,    -9,   -38,    -7,     6,   -20,   -11,   -16,     5,     4,    17,     4,    19,     1,   -16,   -51,   -76,   -47,    -9,    -6,   -35,    -2,     6,    13,    46,    37,    34,    15,   -24,    -8,   -33,   -36,    12,     7,    -7,   -26,    -9,    -8,    20,    -5,    -4,     3,   -22,   -50,   -43,   -38,     4,   -13,    19,    28,     3,    26,    40,    18,     0,     5,     6,     7,   -16,   -26,     6,    17,     8,     7,   -11,     0,   -20,    11,    -2,    15,    17,    -9,   -51,   -29,    -2,    -9,    33,    24,    30,    55,    23,     1,    11,    24,     4,    12,    -9,    10,     2,    27,     7,     6,     6,     7,   -10,    -1,    -2,    17,   -22,    10,   -62,     3,    -2,    -6,   -27,    -4,    18,    35,    54,    12,   -10,     3,    -8,   -14,     5,     2,    -5,   -13,    -1,    -1,    10,    -3,     5,    10,     9,     3,   -14,     9,     8,     0,     2,    -2,   -50,   -26,    -5,     5,    -6,    22,     1,     7,    -4,    13,    -9,   -10,    19,    10,    12,    21,    -5,    23,    11,    -5,   -17,     4,     5,    16,    38,    -2,    -2,    -2,    15,    -7,     6,     2,    13,     9,    -9,    -7,    27,    13,    16,    24,    17,    16,    12,     7,   -42,   -15,     4,   -10,   -23,    -4,    24,    20,    45,    -5,    -1,    -5,   -27,   -18,   -34,    -4,     0,     0,    17,    21,     7,     9,    18,    26,    23,    16,    24,    10,    11,     1,    -9,    -7,   -10,   -28,     7,   -46,   -21,    -3,    -2,    -4,    -6,    23,   -50,   -47,    -1,   -10,     2,   -10,    -3,    -4,    -1,     8,   -16,    25,    28,    24,     8,    26,    24,    25,    46,    41,    31,   -12,    -2,    -5,    -1,     5,     2,   -17,   -28,   -35,   -45,   -62,   -30,   -12,    -8,    13,    26,    62,    33,    44,    12,     3,   -13,    12,     1,     2,    -1,   -34,   -13,    -1,     0,     2,    -4,    -3,    -5,    -2,     4,     8,    -6,    -7,   -10,    -9,     3,    -1,     5,    -5,   -50,   -24,    -7,    -5,   -15,   -13,   -32,   -41,   -28,   -23,    -5,     3,    -3,     5),
		    86 => (    0,     1,    -5,     3,     4,     0,     2,    -3,     0,     1,     3,     3,    17,    12,    -3,     0,     2,    -2,    -3,     1,     2,    -3,     1,    -4,     3,    -2,    -5,     0,    -4,    -2,    -3,    -5,     2,     1,    15,    19,    17,    20,    21,     8,    23,    17,   -26,     2,    -3,    15,    12,    19,    25,     8,     5,    -3,    -4,     3,     2,    -2,    -1,    -5,     8,    -2,    11,     4,    19,    13,    21,    27,    15,    12,    23,    12,     9,     1,    15,    15,    23,    26,    42,    36,    26,    12,     5,    13,    -5,    -4,    -5,    -2,   -17,    -3,     4,    18,    34,    38,    35,    35,    41,    32,    19,    29,    20,    -7,     3,    27,    25,    -1,     9,    33,    38,    35,    26,    -9,    -2,    -2,     1,     3,   -35,   -17,    15,    34,    42,    28,    10,    25,    38,    20,    29,    -3,     9,   -12,    15,    20,     5,    13,    30,   -13,     1,    17,    15,    17,    -6,    11,    -3,    -1,   -22,   -20,    18,    22,    16,    21,    25,    30,    35,    11,    18,    -2,     5,    -1,    19,    10,   -18,   -13,     3,    -9,    15,    17,    19,    30,    11,     7,    -3,     1,     0,    -8,    19,     6,    25,     9,     5,    29,    38,    10,   -10,   -12,   -11,    -7,     3,    -6,     9,     6,     6,    25,     8,    12,    13,    12,    -3,    -9,     1,     3,    -2,   -15,     9,    10,     4,    28,    19,    34,    16,     3,    -1,   -14,    -3,   -13,     0,     8,    32,     7,    22,     9,    -6,   -16,     9,    -2,   -13,   -23,    -2,    -3,   -15,   -23,    23,     8,    -7,     9,    16,    16,    16,     0,     8,   -14,     8,   -10,   -18,    31,   -15,     9,    17,    32,   -25,   -31,   -33,   -46,   -29,   -39,     2,    -4,   -23,   -25,     8,    -4,    -9,     3,    12,    -1,     1,    10,     6,    -6,     0,   -13,   -20,   -33,   -21,    13,    15,    -9,   -29,   -25,    -8,   -39,   -15,   -34,     2,     1,   -19,   -30,     6,   -14,   -12,   -12,    -9,     3,     4,   -12,     9,     2,     4,   -25,   -30,   -35,   -20,    11,     0,   -16,   -34,   -32,   -33,   -11,   -16,   -49,     0,    -2,   -18,   -38,    -4,    -3,    -1,   -19,   -31,   -12,    -6,     9,    12,    -8,   -20,   -16,   -12,   -10,    11,    12,    -1,   -14,   -23,   -14,   -19,   -12,   -37,   -14,    -2,     1,    -4,   -24,    -6,     4,    -9,   -21,   -48,    -3,    -2,     4,    -1,    -6,   -10,    -1,    14,    38,    31,     8,   -12,     6,   -17,    29,    10,   -13,   -37,   -13,    -2,     0,    -6,   -25,    -5,   -12,   -15,   -47,   -59,   -22,    -7,    -5,   -11,     6,   -12,     6,    20,   -10,    -5,    10,   -11,    10,    -2,    38,   -18,   -21,   -31,    -2,    -4,     0,    -5,   -27,   -24,   -11,   -30,   -29,   -36,   -20,    -2,     0,    -1,    -5,     1,    10,     3,   -13,   -23,   -12,   -13,     0,    12,    27,    -4,    -4,    -5,     0,     4,    -5,    -8,   -25,   -36,   -21,   -21,    -8,   -53,   -45,   -19,     1,    -5,    -8,   -13,    12,     9,   -20,   -17,     5,    -7,     1,     4,    -2,     0,    11,   -26,   -39,     4,    -5,   -13,   -45,    -7,    12,   -19,    -5,   -39,   -18,    -8,    -4,   -13,   -24,   -12,     2,     7,    -1,     7,    -3,    -5,     5,     3,     4,     9,     8,   -26,   -35,     0,     0,   -11,   -39,     8,   -12,    -1,     7,    -4,     4,     9,    16,   -13,   -30,   -18,    -9,     5,    -4,    11,     3,    -4,   -10,    -2,    20,    24,    17,   -18,   -44,     1,    -4,    -7,   -49,    -7,   -15,    -5,     3,     5,    22,    31,    27,    15,    -8,    -4,     7,     7,    20,    21,     8,    16,    16,    -7,    12,    17,    26,   -19,   -21,     4,   -13,   -41,   -37,     0,   -12,    15,    19,    23,     4,    45,    41,    30,     7,    13,    -1,     0,    -6,    -3,     9,     8,     1,    -3,    -5,     2,     0,   -14,    -8,     3,   -11,   -11,   -30,   -11,   -14,   -16,    39,    32,    34,    52,    42,    42,    23,    32,    34,    -2,   -18,    -5,   -22,     4,    -3,    -9,   -12,   -29,    -6,   -31,    -1,     5,    -1,   -28,   -13,   -15,   -27,   -16,    25,    73,    44,    35,    16,    24,    24,    29,     8,    -6,    -9,   -10,    15,     9,    -5,    -6,    -7,   -46,   -38,   -26,    -5,    -3,    -4,    -6,   -18,   -31,   -44,   -32,     3,    20,    34,    26,    21,    15,     3,     4,    -4,   -16,   -12,   -11,    -1,    13,    12,    -5,   -15,   -60,   -36,   -22,    -1,     5,     0,    -2,   -25,   -16,   -22,   -25,   -24,   -26,    -1,    -2,    -5,     1,    -4,    -4,    10,    10,   -26,    -9,    24,    15,    -7,   -26,   -41,   -48,   -17,   -18,    -5,    -1,     3,     2,     0,   -12,   -10,    -5,   -27,   -49,   -50,   -50,   -63,   -32,   -44,   -30,     1,    25,    33,    22,   -18,   -11,   -41,   -23,   -23,   -14,    -5,     2,     4,     3,     2,    -2,     3,    -5,   -15,   -21,   -35,   -25,   -18,   -22,     1,    16,     7,   -13,   -18,   -20,   -19,   -19,    -8,   -36,   -19,   -22,   -30,    -9,     1,     5,    -2,    -5,    -2,    -1,     0,    -9,   -12,    -2,     2,     0,     3,    -9,   -12,    -3,     5,    -7,    -9,     0,     4,    -1,     0,   -11,    -5,    -6,    -8,    -4,    -1,    -3,     1,    -2,    -3,     0,     4,    -3,    -2,     2,     2,    -4,    -1,    -4,     5,    -3,     1,     0,     0,    -1,     4,    -6,    -1,    -3,    -6,    -2,     4,     3,    -3,    -2,     3),
		    87 => (    2,    -2,     3,     1,     3,    -3,    -4,     1,     4,    -4,     3,     1,     4,     1,    -1,     1,     3,     3,    -2,     3,     2,     2,     1,     3,     5,    -3,     1,    -5,     3,     0,    -2,     4,     1,     1,    -4,    -4,     2,     0,    -1,   -11,   -17,   -13,    -1,   -22,   -40,   -35,    -2,    -2,    -1,     3,    -1,    -5,     1,     4,    -4,    -2,     0,    -3,     2,     2,    -7,    -1,     3,    -4,    -4,    -7,   -24,   -44,    -6,    -5,    -1,   -31,   -11,   -14,   -11,    -6,    -1,    -4,    -2,    -2,    -1,     3,     3,     4,     2,     0,     4,    -8,    -5,   -10,   -21,   -38,   -27,   -24,   -13,   -19,   -28,   -23,   -17,   -23,   -23,   -17,   -12,   -28,   -10,   -10,   -14,    -3,    -2,    -5,     1,     3,     3,     4,     0,     2,   -27,   -18,   -12,   -48,   -47,   -42,   -85,   -31,   -16,    -3,    -6,   -14,   -38,   -29,   -28,   -30,   -31,    25,     2,   -26,   -32,   -17,    -7,    -3,     4,    -5,     2,   -40,   -17,    37,     5,    24,    12,    18,   -17,   -45,   -50,    -1,   -19,   -31,   -16,   -30,   -39,   -20,   -16,   -12,   -18,   -46,   -19,   -28,    -3,     1,     4,    -2,    21,    28,    23,    36,    25,    26,    15,    19,    41,    -3,     3,   -25,   -23,   -26,   -12,    -6,   -20,     1,    -2,     1,    13,   -38,    -7,   -26,   -13,   -10,     0,     7,    28,     1,    44,    41,    48,    57,     9,    51,    47,    21,    19,    13,     7,    -9,   -15,    -2,     7,     2,     6,    -1,    42,    10,    -7,   -27,    -7,   -14,   -17,    -6,     1,     4,     5,    19,     9,    38,     8,    25,    24,    20,    34,     7,    14,    12,     1,    -4,    -7,     4,    -3,    -3,    32,     0,   -23,   -40,   -25,   -19,    -4,     1,    36,    17,    14,     2,     1,    13,    12,     1,     2,     8,    38,    21,    32,    15,     4,     1,    -6,     1,     9,     1,    20,     9,   -41,     6,    31,    60,    -3,   -17,    14,    -5,   -15,   -11,    -9,   -14,     9,     1,    -8,   -20,   -20,     3,    -6,    -3,     3,    18,    13,    -9,    11,   -16,   -12,   -13,   -15,    22,    30,    56,     4,   -10,    12,   -12,   -15,   -28,   -15,   -12,   -14,    -7,   -32,    -7,   -28,   -40,   -12,    -2,    -7,    -4,   -17,    -9,     4,   -24,     1,     9,   -30,   -39,   -29,     7,     1,    11,   -18,   -22,   -17,   -31,   -30,   -34,   -40,   -52,   -61,   -24,   -32,   -23,   -17,     9,    10,    -1,     5,     6,     4,    -7,   -17,   -19,   -70,    -9,   -34,     6,     1,     0,     9,   -26,   -48,   -19,   -17,   -26,   -29,   -22,   -28,   -21,   -11,   -20,    -9,    24,    -6,     9,    11,    -1,   -29,    17,   -13,    -3,   -36,   -22,   -28,   -15,    -6,     4,    -5,    -9,   -15,   -10,     0,     0,   -17,   -14,     9,     4,    12,     7,    13,    10,   -17,    26,    13,    24,    -2,    16,    -3,    11,     3,   -23,   -20,    -2,     3,    -2,    -5,     0,    -4,     0,    -1,    -8,   -24,    -4,   -15,    -8,    -1,     7,     3,     7,   -18,    15,    19,     1,   -25,    32,    -1,    14,    -4,   -21,    -7,   -18,     5,    -7,    -1,   -16,    -5,    -5,   -10,    -5,   -11,     0,    15,    -8,    11,    20,     0,    -4,    -3,    -3,     8,     3,    10,     3,    -8,   -17,     5,   -47,   -36,    -5,    -1,     5,   -29,   -27,   -31,   -20,    16,    19,     3,    20,    23,     7,    12,     0,     0,    -7,    11,    -6,   -23,   -10,     9,     1,     4,    -5,     3,   -19,     8,   -22,     5,     2,    -4,   -16,   -21,    -3,   -15,    21,     3,     4,     4,    -2,     0,    -3,   -13,   -15,   -19,    -8,   -22,   -11,    -4,   -26,    -8,    -8,   -12,   -23,    18,   -21,    -1,     4,    -5,    -3,   -19,   -31,    -9,     4,     3,    -4,   -19,     4,    -3,     6,     3,   -10,   -23,   -15,   -41,   -22,   -28,   -43,   -18,    -5,    25,    -5,   -27,   -12,    -4,    19,    -6,   -15,   -51,   -44,   -22,     0,     5,    -5,   -18,     7,    -5,     1,    -6,   -17,   -10,   -45,   -51,   -32,   -30,   -33,   -43,     3,     4,   -34,   -29,    -4,    -3,    -4,   -11,   -34,   -20,   -23,   -26,   -44,   -33,   -27,   -11,   -12,     1,     4,   -12,   -13,   -17,   -32,   -39,   -29,   -36,   -25,   -35,     0,    -4,   -15,    -6,     2,    -7,    -4,    -8,   -45,     2,   -10,   -14,    -7,   -36,   -30,    -7,    -5,    -5,   -12,   -21,     2,    -7,     2,   -17,   -13,   -24,   -73,   -58,   -39,   -21,    -5,   -28,    -5,    -4,    -2,   -16,   -55,    -6,    -2,     7,    11,   -36,   -15,    -1,    -3,     3,    -1,    -1,     3,   -10,    -4,   -34,   -12,   -22,   -30,   -54,   -24,   -22,   -12,   -28,     3,     0,     1,    11,    -5,    15,    16,    -6,    -8,    -7,   -15,   -26,     0,    -6,     3,    -2,    -8,   -18,    20,   -23,   -10,     9,    12,   -30,   -23,   -20,    -8,    -6,     1,     2,     3,   -14,    14,   -13,   -18,   -15,    34,    15,   -10,   -22,   -15,   -10,    -6,    -3,   -21,     0,    -2,    -8,     2,   -15,    -7,    -9,    -9,   -29,    -6,   -10,     5,     3,     4,    -5,   -18,   -64,   -48,   -56,   -15,    -2,   -13,   -19,   -33,   -24,    -8,     2,    27,     0,   -13,    -1,   -27,     3,    -5,   -10,   -18,    -3,     2,     1,     3,    -3,     4,     4,     1,     2,     4,    -1,   -11,     8,    25,    31,    21,    -6,   -13,   -18,    21,    24,    33,    28,    -7,    -3,    -3,   -14,     1,    -2,    -3,     0,    -4),
		    88 => (   -2,    -2,     1,    -2,    -3,     1,    -5,     5,    -3,    -2,     4,     3,     4,     3,     2,     3,    -3,     2,     3,     2,    -4,     4,    -2,    -1,     3,     4,     0,    -2,    -2,    -1,    -5,    -1,    -3,     0,    -4,     1,    -3,    -4,    -4,    -9,   -14,   -12,   -21,   -50,   -54,   -45,    -9,    -8,   -10,    -6,    -9,    -2,     2,     3,    -5,    -4,     1,     4,    -1,    -1,     1,     0,    -9,    -3,   -20,   -19,   -26,   -31,   -21,   -11,    -1,   -26,   -33,    10,    15,    -1,   -21,   -31,   -33,    -4,    -6,    -8,    -3,    -1,     1,     2,    -4,   -11,    -9,   -40,   -34,   -42,   -27,   -15,    10,    14,    17,     4,    -5,   -25,   -36,   -49,   -23,    -8,     8,    20,     2,    11,    12,   -12,    -5,     3,    -4,     2,     6,    -2,   -21,   -44,   -31,   -31,    17,     9,    35,    35,     6,   -33,    -1,   -16,   -15,     5,    -1,   -21,   -16,     5,   -20,     7,    13,    12,     8,    -9,     0,    -3,   -15,   -13,   -40,   -34,   -37,     2,   -12,    12,    26,    21,     6,    17,     3,    19,    21,    28,    11,     0,    -1,   -10,   -30,   -25,    15,     6,   -13,   -18,     4,     4,   -32,   -30,     8,   -27,   -36,   -22,    -3,    -6,     9,     6,   -10,    -2,    13,    20,    19,     7,    11,   -17,    -8,    -1,    12,    10,     4,    14,    -1,    -5,     1,   -30,   -17,     8,    16,   -13,   -21,    -2,     8,    12,     3,    -1,    -7,    -4,     1,    29,    30,    10,    -4,   -12,    10,    10,    23,    29,    11,     6,     3,   -20,   -16,   -21,   -17,    41,    21,     1,    10,    11,   -22,     5,    11,     0,    -4,     5,     6,    14,    13,     8,     9,    -6,    -6,   -13,    -1,    16,    -9,    10,    15,     4,     3,   -15,   -23,    23,    44,     0,     3,   -13,    -9,     5,     3,   -16,    -8,   -11,     3,    12,    -5,   -16,    -4,     6,     2,    -2,   -12,     3,    -4,    29,    42,   -31,    -5,   -15,   -31,   -19,    22,    -2,    -6,     0,   -17,   -22,   -21,   -24,   -13,    16,    18,    -8,   -37,   -26,   -21,   -16,    -3,   -15,     9,    10,    14,    11,    30,   -26,     5,    -8,   -23,   -11,    16,    -2,    14,    -8,   -13,    -9,   -31,   -16,    -3,    14,     0,   -43,   -40,   -24,   -18,    -5,   -10,    -7,    -9,    24,     8,   -20,    17,   -23,     2,    -3,    -4,     5,   -22,    -2,   -28,   -35,   -20,   -22,    -7,    16,    17,    11,    12,     1,   -15,   -24,   -10,   -13,     5,     2,    11,    -1,   -18,   -53,   -58,   -32,    -4,    -1,     1,   -12,   -26,   -14,   -24,   -21,   -12,    29,    28,    24,    35,    18,     1,    10,    -2,   -12,     4,   -10,    11,    25,    14,     4,   -35,   -47,   -44,     3,    -8,    -4,    -8,   -18,   -24,    -2,     9,   -12,    12,    33,    34,    40,    31,    21,     3,    11,    -3,    -9,     0,    18,    21,    20,    -7,   -21,   -19,     3,   -24,   -11,    -6,    -2,   -12,    -5,   -29,    -5,    25,    24,    27,    43,    50,    26,    21,    29,    11,     5,     7,     2,    15,    14,    18,     9,    10,   -24,   -21,    34,   -39,   -13,    -4,     0,   -15,   -14,   -22,   -15,    -7,    20,    10,    33,    40,    35,    12,    -3,    -3,    -2,    18,    37,    33,     8,    23,    14,     1,    -2,     0,    17,   -51,   -18,    -4,    -6,   -24,   -14,     4,   -24,   -28,     0,     3,     4,    14,     4,    -9,   -16,    -6,    22,     2,     6,    13,    11,     4,    -5,    -6,     8,    10,   -12,    -5,   -22,    -4,    -9,   -25,   -38,   -19,   -25,    -9,   -18,   -15,    -2,   -10,   -19,   -19,    -6,    17,    -4,     0,   -18,     4,   -10,   -31,   -28,   -10,    15,    -7,   -30,    -3,    -9,     2,     2,   -13,   -46,   -22,   -38,   -33,   -34,   -30,   -26,   -16,   -18,     3,    19,    22,     8,    18,    -9,   -10,   -21,   -17,    -2,    12,     5,   -15,   -37,   -22,   -15,    -4,     0,   -21,   -43,   -24,   -22,   -20,    -5,     1,   -24,   -13,   -13,    16,    20,    34,    22,    11,     6,   -16,     2,    10,     6,     2,    -1,   -34,   -30,   -28,    -2,   -10,   -11,   -26,    -8,   -19,     0,     4,    -4,     0,    -2,   -13,    23,    55,    22,    16,    31,    20,    18,    -3,     1,     7,   -19,   -12,    -1,   -19,   -15,   -29,    -4,   -10,    -9,   -13,     1,    21,    10,    -4,   -12,   -15,     3,     4,    27,    14,     9,    41,    33,    11,    -4,    -4,   -17,    10,   -13,     9,    13,   -12,   -28,   -27,    -7,    -4,    -2,    -7,    -3,    11,     5,   -11,   -23,   -13,    21,    25,     3,    18,    41,    29,    21,    12,   -15,    -5,     0,    18,     3,    14,    18,   -40,   -33,   -18,    -1,     1,     3,   -14,   -11,    -8,   -16,   -18,   -25,   -17,     3,    -4,     9,    34,    45,    30,     3,    -7,   -18,     6,    38,    30,     7,   -28,   -14,   -46,   -23,   -11,    -1,    -2,     0,   -14,    -3,   -50,   -34,    -2,   -15,   -32,   -33,    -5,    22,    20,    28,    10,     6,   -31,   -12,     3,     6,   -17,   -45,   -44,   -28,   -24,    -9,   -17,    -4,     4,     0,     2,   -20,   -18,   -20,   -32,   -24,    26,    15,   -18,    -9,    -6,    11,    -4,   -41,   -20,   -14,   -27,   -28,   -54,   -42,   -22,   -16,    -5,    -1,     1,    -3,     0,    -2,     1,     1,     0,    -8,    -6,    -1,   -26,   -36,   -20,    -6,    -6,   -23,   -43,   -30,   -32,   -27,   -16,    -9,    -3,    -1,    -8,    -3,     4,     4,    -1,    -3),
		    89 => (    0,    -4,     3,     3,    -4,     1,     4,    -2,     2,     0,     1,     1,    -3,     2,     2,    -4,     5,    -4,     0,     1,    -1,     0,     0,     3,     2,     5,     2,    -2,     3,     2,     5,     4,     3,    -1,     1,    -2,    -1,     3,    -1,   -12,   -25,   -16,    -1,    -2,    -7,    -2,   -18,   -14,     2,    -7,    -6,     0,     5,     0,     3,     2,     3,     2,    -4,   -21,   -10,     0,    -2,    -8,    -6,    -1,    -6,   -19,    -1,    -6,   -28,   -11,    -9,    -7,   -10,   -11,   -14,    -7,    -7,    -2,    -6,     0,     0,    -5,    -1,     5,     4,   -12,   -20,   -23,   -19,   -24,    -6,   -10,    -3,   -15,   -13,   -20,   -28,   -24,   -20,   -21,   -33,   -21,   -14,   -13,   -12,    -4,    -3,    -5,     1,     4,    -1,     4,    -3,    -4,   -13,    -5,   -27,     4,   -16,    -8,   -10,   -23,   -38,   -30,   -19,   -17,    -8,    -8,   -19,   -32,   -37,   -18,   -10,    -9,    -3,   -25,    -5,     4,    -2,     2,     2,   -11,     1,    -3,    -6,   -10,   -11,   -15,   -35,   -13,   -14,   -13,    -1,    -4,     2,   -14,    -8,   -17,    -2,    -6,   -20,   -13,    -3,    -9,   -11,    -3,     1,    -1,    -5,   -14,     0,    -6,   -21,   -20,   -46,   -22,   -16,   -18,   -10,    11,    33,    19,    11,    14,     0,     3,    10,    -1,   -16,   -18,    -9,   -16,    -7,   -10,     2,     0,   -11,     0,   -14,   -27,   -35,   -33,   -48,    -3,    -9,    13,    14,    -1,    -9,    14,    -2,    -1,   -10,    -2,    -3,    -6,   -17,   -15,   -27,   -11,    -2,    -8,   -15,   -13,    -5,   -16,    -5,   -31,   -23,   -48,   -17,   -21,    11,    -1,   -13,    -1,    -1,   -41,   -16,    -2,    -5,    -5,     3,   -17,   -12,   -26,   -39,   -11,    -7,     0,     2,    -2,    -8,   -13,   -30,   -37,   -23,   -35,     1,    10,    -2,    13,    -7,    -8,     6,   -20,   -20,    -8,    22,     8,     6,   -20,   -15,    -8,   -15,   -37,    -3,   -16,     4,    -9,   -16,     1,    -5,   -11,   -18,    10,     9,     4,   -23,   -16,   -36,   -28,   -15,   -19,   -35,   -22,    21,     2,    -6,   -28,   -11,     1,   -18,    -4,    -5,   -13,     1,   -33,    -3,    14,    -3,   -14,   -13,    -3,     9,    -7,   -16,   -44,   -26,    -4,   -10,   -17,   -20,     1,   -13,     0,    -2,   -10,    -6,    14,   -22,   -10,    -4,   -14,    -5,    -6,     4,    12,     7,     7,     4,    -3,    17,   -10,   -18,   -36,    -9,   -23,   -38,   -24,   -14,   -10,   -27,    -5,     1,    13,    -1,     5,   -43,   -18,    -4,    -7,    -4,   -21,   -16,    22,    20,     9,     5,     1,    -6,   -29,   -17,   -20,   -33,   -26,   -10,    -7,     8,   -25,   -27,    -4,    -4,    15,     0,   -14,   -30,   -19,    -7,    -3,    -5,   -16,   -24,    -2,    12,     8,     7,     5,    22,   -28,   -13,   -43,   -31,   -20,   -14,     9,     4,   -15,    13,    13,     1,     3,     7,   -34,   -21,   -12,     7,    -4,     0,    -3,   -22,    -6,     2,     1,    15,    10,    12,   -22,   -10,   -41,   -35,   -33,   -18,   -15,   -17,   -27,    10,     9,    21,     8,     4,   -51,   -36,    -9,     4,    -2,     4,    -2,   -24,   -18,    12,   -14,    23,    -2,     3,   -10,    13,    -9,     1,    -9,   -19,   -25,   -30,   -15,    25,    10,    14,   -11,    -7,   -39,   -16,   -18,    -3,     2,     2,    -3,   -18,   -16,    17,   -17,     0,    20,   -18,    -1,    -4,    -5,    -6,   -25,   -10,    -2,     2,     0,     9,     7,    11,   -12,    -8,   -23,    -6,    -8,   -15,    -6,     0,     3,   -19,   -10,    17,    14,    12,    -3,   -12,    -3,    25,    10,    16,     4,     8,   -10,   -14,    12,    17,     6,   -10,     6,    11,   -18,   -36,    -1,   -19,   -14,    -3,    -1,   -12,    -7,     7,    33,    25,    39,   -11,     4,    23,    50,    12,    -6,   -15,    -3,    -3,     2,    22,   -15,    -5,   -10,    -5,   -20,   -12,     9,   -20,    -3,     2,    -6,    -8,    -9,    -2,    14,     7,    -5,     5,     9,    -3,    -1,    -3,   -15,   -34,   -15,   -11,     9,    24,   -11,    -8,     2,    -5,    -7,    27,    11,   -19,     0,     2,     3,   -19,   -12,   -28,    -8,     4,    18,    10,     2,    -2,    -6,   -14,   -13,   -12,    -1,     3,    -2,    12,     4,     7,   -18,     0,     2,    33,    -7,   -38,     5,    -3,     3,    -7,   -10,   -17,   -16,   -20,   -20,    -2,    -3,   -13,   -21,    -9,   -24,    15,     5,    -6,    -5,    -1,     3,     7,    -3,    11,    -6,    26,     6,   -30,     1,    -2,    -2,    -4,     6,   -17,   -19,   -17,   -24,   -24,   -42,   -45,   -41,   -34,    -7,     9,    21,   -17,    -7,   -18,    14,     4,    11,    34,    -3,    29,    10,   -18,    -1,     2,     0,    -9,     2,    -2,    -4,    -9,    -6,   -15,   -20,   -39,   -36,    -8,    28,    -6,    -1,     0,    -9,     5,    12,    20,    24,    32,    22,    24,     9,    -2,     3,    -2,    -3,    17,   -12,   -11,     5,    -4,   -13,   -12,   -19,    -1,     6,    19,    27,    -3,   -16,   -20,   -26,    -7,    31,    38,    24,    39,    18,    15,    -8,    -9,     2,     1,     2,     2,     6,    11,     2,    -1,     4,    -2,    -2,    -1,    -3,    -9,   -19,   -11,   -34,   -44,   -23,    -5,     4,    29,    17,    12,    15,    -2,     0,     4,     5,    -1,    -3,     0,     4,    -8,    -2,    -1,     1,     1,     1,     4,     4,    -3,    -2,   -13,    -6,   -17,   -28,   -20,   -19,   -12,   -16,     2,    -6,     2,     0,     1,     3),
		    90 => (   -5,     2,    -3,     2,     2,    -2,    -4,     2,    -1,    -2,     3,     2,     1,     4,     1,    -4,    -3,     4,    -5,     4,     1,    -1,     1,     1,    -4,     4,     2,    -4,    -4,     0,    -3,     5,     0,     2,    -3,    -3,    -3,     0,    -4,    -4,     4,     4,    -6,    -4,    -1,     3,     1,     3,    -1,     1,    -5,    -1,     5,     1,     0,    -2,     3,    -4,     1,     5,    -1,     1,   -11,    -6,    -7,   -11,   -10,    -6,    -9,   -13,    -9,    -5,    -2,     3,    -1,    -5,    -2,     0,    -3,    -7,    -5,     2,     1,     0,     0,    -4,     1,     5,    -6,     1,    -6,     0,     3,    -4,    -6,   -10,   -18,    -8,    -5,    -6,     5,    11,    10,     1,     0,     1,    -5,    -9,     5,     4,    -1,     0,     4,    -2,     4,    -7,    -6,   -18,   -13,     7,     4,     1,    -2,   -14,    -9,   -10,    -7,    -6,    13,    17,     7,    15,    15,     1,    -3,    -6,    -1,    -4,    -6,     3,     5,     2,    -4,     3,    -1,    -5,     4,   -16,    -6,    -9,    -9,    -4,     2,     3,    -7,    -6,     1,    -7,     1,    20,    20,     2,    -6,    -5,    -5,    -5,    -4,   -14,     5,    -2,    -8,    -7,    -5,   -12,     4,     7,     3,   -10,    -8,    -3,    -6,   -11,    -5,    -9,    11,     4,     1,     9,    14,     9,    -6,    -6,    -7,   -21,    -5,     1,     2,    -6,   -10,   -11,    -2,     6,    16,     3,    -8,     8,     7,     3,     7,     5,     0,    19,     5,    11,    23,     7,     1,     5,    14,    -1,    -4,     0,   -12,     1,     1,    -4,    11,   -10,     8,     9,     6,    13,     6,   -12,    -9,     3,    11,   -10,    -3,    -8,     1,     8,     3,     7,    18,    16,     9,    10,    -7,    -5,   -11,    -7,    -5,     0,     5,    -2,    23,     3,    -6,    -1,     7,     8,    -6,   -24,   -26,   -21,   -19,   -20,   -10,    -4,    -2,     0,     2,    21,    12,    -5,     6,    -7,    -1,    -4,     3,     2,     2,     1,    -2,    19,    17,    15,    13,     2,   -23,   -19,   -22,   -15,   -11,     2,   -22,   -15,   -15,    -8,   -10,   -12,    15,     4,    -5,    -8,   -11,    -1,     4,    15,     2,    -5,    12,    20,     8,   -11,     2,   -21,   -24,   -33,   -26,     1,     5,     7,   -12,   -14,   -22,   -31,   -26,   -15,     1,     3,    17,     1,    -2,    -2,    -3,    -2,     3,    -5,    14,     9,     6,    -8,    -3,   -17,   -28,   -33,   -21,     1,    -4,    -8,   -31,   -36,   -22,   -23,   -24,   -10,    -1,    -6,    10,     8,    -4,     5,     5,    -3,     1,     2,    23,     3,    21,   -10,   -12,   -25,   -37,   -38,   -18,   -10,    -4,   -13,   -28,   -23,   -27,   -26,   -25,   -12,     2,    11,    11,     4,     1,    -8,     3,    -1,    -1,   -15,    26,    16,    -6,   -19,   -27,   -31,   -27,   -24,   -23,   -18,   -11,   -26,   -23,   -20,   -22,   -23,   -23,   -11,   -15,    -6,   -12,     8,    -8,    -3,    -4,     3,    -1,     2,    23,    11,    -4,   -14,   -18,   -27,   -22,   -23,   -13,   -13,   -13,    -4,   -10,   -19,   -17,   -20,   -22,   -10,     3,    -1,    -8,     2,    -6,     0,     3,     2,    -9,    -1,    13,    18,    13,    -3,    -9,   -13,   -16,   -14,   -17,   -13,    12,   -10,   -10,   -30,   -29,   -28,   -12,   -20,    -5,    20,     0,     8,   -12,     6,     3,    -3,    -9,    11,    20,    15,    16,    16,   -10,   -14,     3,    -1,   -10,   -12,    -8,   -16,   -31,   -30,   -30,   -26,   -17,     1,    12,    -2,    -4,     7,   -27,     5,     2,    -2,    -5,    -2,    29,     9,     8,    15,    -4,    -4,    -1,   -11,    -5,    -9,   -24,   -11,   -24,   -25,   -35,   -20,   -10,    10,     2,     6,     2,    -5,    -6,    -3,     4,     1,     5,    -1,    19,     2,     4,     8,    -4,     2,     6,    -4,     0,    -8,    -8,   -12,   -18,    -7,    -8,    -3,    12,     0,     2,    -9,     2,   -17,    -9,     2,    -5,     0,     4,     0,    14,    -7,    14,     8,     3,   -13,    -8,     5,    -9,     1,     6,    -1,    10,    12,   -14,    -4,     3,    -3,     8,    -6,    -2,   -12,    -2,     0,     2,     1,    -6,     0,     1,   -16,     2,    19,     1,     1,    -4,     9,    -9,     0,    -2,    -1,   -10,     3,     2,     9,     7,     3,   -11,    -1,    -9,    -1,     4,     5,     5,    -2,    -3,    -8,   -11,    -6,   -14,    15,     5,    -5,     3,     7,    -7,     2,    -5,   -11,    10,    11,    -2,     4,     4,    -8,    -5,    -7,   -12,     1,     6,     6,     5,    -1,    -1,   -10,    -6,    -7,     7,    13,    -5,    -9,    -3,     0,     5,   -11,    -4,    -2,   -12,    -2,    -8,     5,    -1,     1,     0,   -12,   -16,   -13,   -12,    -2,    -3,    -3,    -5,    -4,    -8,    -4,    18,    14,     9,   -10,    -2,    -3,   -10,     5,    11,     9,     3,     6,     8,    -7,    -9,     1,    -3,    -6,     0,     0,    -3,     4,    -4,     1,     2,     0,    -6,    -4,    11,    20,    20,     5,     1,     0,    -8,    -7,   -14,     1,    -1,    -9,   -22,   -29,   -26,   -18,   -17,   -11,    -3,    -4,    -2,    -1,     3,     4,     3,     0,    -1,   -11,   -17,     0,    -5,    -1,    -6,    -2,     2,   -11,   -11,    -8,   -13,   -39,   -21,   -21,   -22,   -15,    -6,   -16,     0,    -4,     3,    -3,     4,     0,    -3,     0,     2,    -2,     0,    -2,     1,    -4,     0,    -2,     4,    -7,    -6,    -2,    -1,    -1,     0,    -5,     2,   -10,   -13,   -12,    -1,    -2,     0,    -5),
		    91 => (   -2,    -1,     3,    -2,     3,    -2,    -3,    -1,     3,     2,    -1,     2,     4,    -3,    -1,     5,     5,     4,     4,    -2,    -4,    -1,     2,     4,     2,     4,     4,    -3,    -1,     2,    -1,     3,    -2,     5,    -1,     0,     2,    -1,    -2,    -3,    -2,    -9,    26,    13,    15,   -16,    -5,    -1,    -3,    -2,    -3,     0,    -3,     1,     0,     3,    -2,     4,    -3,     3,     4,    -5,     2,     4,   -16,   -17,   -12,   -14,    -5,     9,     9,    18,    42,    25,    23,     8,    13,   -27,   -20,   -26,    -2,     0,    -5,    -1,     0,    -3,    32,    15,    -3,   -16,   -29,    17,     5,     4,   -22,   -36,   -16,    -1,    -3,     2,     8,     1,     3,   -22,    -7,   -16,   -14,   -17,   -13,    -2,    -1,    -2,     3,    -2,    31,    29,    25,     2,    -8,    10,    21,    18,    10,     3,   -23,     5,    -8,     9,    -5,    -2,    -2,   -23,   -24,   -12,    23,    18,    16,   -11,    -8,   -13,    -1,    -5,    12,     8,    34,    29,     5,     5,    20,     3,    -5,    -4,   -10,   -11,   -23,    -6,    -6,    -8,   -12,    -9,   -27,     9,    23,    30,    24,   -20,   -11,   -17,    -5,    -4,   -15,     1,    34,    13,    11,    -3,   -21,   -16,    -6,    -8,    10,   -12,    -7,   -16,   -21,   -15,   -11,   -39,   -12,    15,    26,    24,     8,    -1,    -7,    -7,     4,    -1,   -17,   -20,   -18,   -14,   -21,    12,   -38,    -8,    35,    26,    22,    -5,     6,   -14,   -31,   -16,    -8,   -26,    -8,    19,    26,    29,     6,   -14,   -19,    -7,    -4,     1,   -22,   -15,   -18,   -18,   -17,    24,   -31,    -8,    32,    -2,    21,    -1,    -9,   -11,   -15,   -25,   -23,   -23,    12,    14,    14,     4,     4,   -10,   -22,    -9,     0,    -1,   -20,     0,   -15,   -20,   -12,    29,   -10,     5,    14,    -1,   -17,   -21,   -17,   -13,   -22,   -40,   -23,   -33,     4,     2,    12,    10,     3,    -5,   -19,   -10,    -3,    -3,   -14,    -1,   -14,   -10,   -20,    10,     7,   -13,    22,     3,     2,    -1,    -5,   -13,   -33,   -29,    -7,    -8,     0,     2,    12,    19,   -12,    -2,     4,     9,    -4,     3,    -2,     0,     1,   -15,   -27,    12,   -20,    -8,    -2,   -12,    -6,   -13,    14,     1,   -26,    -9,    -6,    -8,    -7,   -14,    17,    10,   -11,     3,     0,    24,    -5,     4,   -15,     0,     4,    -9,   -12,   -14,   -26,   -22,     2,     0,    -7,   -15,     7,    -8,    -8,    -6,    -4,    -8,    -9,   -15,     1,     6,   -19,     7,    14,    27,     3,    -2,   -11,    -1,    -6,   -11,    -3,    -4,     2,    -6,    -8,   -12,     5,   -11,     1,     3,   -14,    -9,   -23,   -10,   -16,   -20,   -18,   -40,   -19,    18,     5,     4,    -1,     4,     6,     6,    -8,   -16,     5,    -8,   -10,   -17,   -34,   -46,   -16,    14,    10,    11,     1,    -5,    -7,   -31,   -23,   -27,   -30,   -17,   -11,   -22,    -1,     1,     3,     2,    -2,    -2,   -11,   -34,   -17,   -17,   -23,   -35,   -52,   -44,   -16,     9,    19,   -15,   -21,     8,     3,   -25,   -29,   -14,   -28,   -15,   -36,   -32,   -26,    -7,     2,    -4,     0,    -2,   -11,    -8,   -16,   -17,   -24,    -5,   -21,   -14,   -23,    -7,    24,     6,   -11,     7,     5,    -8,    -7,    -3,     0,   -13,    23,   -33,   -25,    -7,     5,    -1,    -2,    -7,    -4,    -4,    -7,   -11,     4,     1,    12,     4,   -17,    -6,    15,    -4,    11,   -10,     9,     4,    16,    14,    13,    -4,     0,   -25,   -18,   -17,     3,    -5,    -3,   -18,   -11,     2,   -21,    -1,    13,    26,    15,   -23,   -27,   -19,     8,     4,     4,    17,     4,     7,   -16,    -6,     7,     1,     6,    -1,   -16,     1,    -5,     0,    10,   -17,   -10,    -3,    29,    32,    41,    37,    30,     4,   -30,    -2,    -5,    13,    20,     3,     6,   -14,    -2,     1,    19,    43,    14,    13,   -16,    -7,     4,     1,    -2,    -9,    10,    20,    29,    34,    22,    20,    17,    -1,   -12,    -3,    11,     0,    12,     2,     3,     6,    27,    24,    30,    17,    10,     1,   -12,    -3,     8,    10,    -4,    -3,   -10,   -21,   -12,    -1,    -3,   -11,   -12,   -23,    -6,     4,   -16,     2,   -20,   -12,     2,    11,    10,    -4,    14,     5,    -2,    15,    -8,    -1,    14,     6,   -13,    -9,    -9,    17,    -3,   -10,   -27,   -23,   -21,   -27,     4,     3,    -2,     8,   -21,    -8,    -3,    -2,     2,    -1,   -23,   -16,    -5,     0,     5,    -4,    -5,    -4,    -4,   -11,     5,    21,    26,    11,    -3,    -4,     6,     2,    22,     5,   -17,   -17,   -16,    12,   -10,    -7,    19,     2,   -10,   -15,   -13,   -18,    23,     0,     5,     2,     4,    -6,     1,     0,     0,    -9,    -9,    -9,     5,     5,    -6,     1,   -16,   -34,   -15,   -18,   -11,   -29,    -3,   -26,   -10,   -10,   -23,    15,    21,     3,    -4,    -1,    -1,   -10,    -8,   -12,    -3,   -10,   -14,    -8,   -15,    -5,    -1,    18,    19,   -12,   -27,   -19,   -19,   -20,   -35,   -24,   -11,    -8,     3,     1,    -2,     1,    -3,    -2,     2,    -8,    -8,   -22,   -21,   -15,    -8,    -7,    -5,    -1,    -6,   -15,   -20,   -15,   -13,   -19,    -3,    -4,    -7,    -8,    -5,    -3,     4,     3,     2,     2,     2,    -4,     1,     3,    -4,     1,    -4,     0,    -3,     4,    -9,   -15,     4,    -4,    -5,     1,    -3,     3,    -3,    -4,     0,     0,     0,    -1,     0,     2,     1,    -2),
		    92 => (    4,     5,     5,     4,     2,     0,    -3,    -4,    -1,    -4,     5,    -5,    -5,    -6,     9,     9,     5,    -3,    -4,    -2,     1,     0,    -4,    -2,     2,     1,    -3,     2,    -3,     3,    -1,     2,    -2,     4,    -5,     6,    -8,   -16,   -22,   -32,    -6,    -9,    -4,    13,    18,     1,   -14,   -39,   -25,   -27,   -18,    -4,     5,    -4,     0,     3,     3,    -3,    -2,   -12,   -13,     1,     5,     2,     2,    33,    32,    37,     3,    10,    28,    46,    38,    17,   -17,   -35,   -19,    -8,   -19,    -6,    -2,     1,     5,     4,    -3,    -1,     2,   -26,   -32,    14,    20,    26,    -1,   -22,   -34,   -44,   -57,     0,    -6,     0,     3,   -18,   -43,   -28,   -24,    -5,     2,   -27,   -30,    -2,    -5,     1,    -3,    -2,    -8,   -21,     0,    11,    47,    37,    27,    46,    13,   -11,   -16,   -17,   -11,     6,   -14,    -4,     6,    -9,    -7,   -21,     3,   -21,   -36,    -3,   -24,    -8,     2,    -3,   -19,   -11,     0,   -20,   -17,     4,    28,     9,    22,     0,     7,     7,    11,     4,    -2,     4,    12,    16,     8,    25,    -9,   -15,   -31,    10,   -43,   -11,    -2,    -2,     3,     1,    10,    -5,    -4,    -6,    20,    -3,     5,   -21,     5,   -17,     1,     0,    12,     7,    18,     8,    -2,     9,    -4,   -13,   -54,    -7,   -39,   -10,    -5,    -4,    15,     1,    19,    43,    12,     6,    13,    -4,   -29,   -15,    -2,     6,    -9,     7,    15,   -14,     4,    -6,     5,    24,    21,   -38,     8,    23,   -25,   -17,   -22,    26,    17,     6,    -4,    36,    14,    -8,    11,     8,    -9,     9,     8,     2,    -3,   -20,   -13,    -5,   -17,     5,     2,   -16,     1,    22,    -7,   -14,   -41,   -12,     3,   -18,     5,    20,   -25,     3,     2,   -12,     1,   -11,     0,    12,    15,    13,   -10,     0,    -8,    -4,     0,    -9,    -2,    -7,    20,    -4,   -18,   -55,    -7,    -9,     5,     2,   -10,    10,   -12,    25,    39,     5,     5,   -13,    23,    -9,     2,     2,    -7,     1,   -10,    26,   -14,   -16,    -4,     6,   -11,   -36,   -21,   -16,   -13,   -17,    -2,   -20,     3,     2,    -8,    11,    19,    14,     5,    12,    15,    -5,   -19,   -26,    -6,   -21,    -4,   -16,    -1,     7,     8,    -3,   -26,   -20,     9,    10,   -13,   -23,    -2,   -11,   -38,     0,   -13,     3,    35,    17,    -1,    24,    -5,   -26,   -15,   -12,   -27,   -20,   -22,   -13,    15,    28,   -10,    24,    21,   -21,    25,     6,    -1,    -6,    -4,   -22,   -14,    -4,    -5,    16,    58,    18,    -9,     3,    -6,    -4,    -7,     6,   -23,   -17,   -21,    -7,    10,    18,    -5,     6,    21,    44,    34,    36,    38,    -6,     3,    -2,    -8,     4,    17,    21,    36,    39,   -22,    14,     4,   -32,   -15,   -21,   -16,   -10,    -8,    -2,    -3,    15,   -29,    13,    37,    66,    54,    28,    24,    11,     0,   -15,    29,    32,    -1,     9,    18,    16,    23,     5,   -11,    -6,    -8,   -18,    -5,    -1,    -7,   -17,    -6,   -14,     8,    22,    21,    19,    -4,    21,    45,    36,    -2,    -2,    37,    34,   -21,   -17,     4,    35,    15,    36,    16,     3,    14,    -3,   -10,    -8,    -5,   -16,   -10,     7,    -9,    70,    57,    35,     7,    40,    48,    27,     0,    -7,    34,    24,    -7,   -13,     7,    -6,    -6,    -5,     4,     1,     2,    -2,    10,    -6,   -11,    -2,    -4,    -5,    21,    73,    41,    16,    12,    19,    19,    17,    -3,     0,     5,    13,    -8,    -6,     3,   -15,     8,    -9,   -14,     2,     6,    -2,   -23,   -12,   -18,   -24,    -3,    18,    64,    56,    43,    31,    24,    21,    -6,     9,     2,   -20,     7,    -9,    -1,    -2,   -12,     0,    11,     8,    12,    17,   -10,   -12,     4,    14,   -11,   -27,    11,    36,    40,    54,    38,    15,    -1,   -12,     8,    27,    -5,   -11,    33,   -17,    -6,    -1,    -2,     1,    -1,    14,    23,    26,     1,     0,   -20,     3,   -22,    -6,    13,    43,    53,    65,    26,    21,    10,     5,     4,    -4,    -3,    -2,    32,   -13,    20,    -6,     6,     0,    23,    37,    21,     1,    11,    10,   -21,    -1,    -5,   -21,    46,    74,    54,    47,    61,     9,   -10,     6,    -7,    -4,     0,     0,   -11,   -23,    -8,     9,   -17,    -1,    20,    19,     7,    10,   -14,    -1,   -14,    -9,     3,    16,    62,    62,    56,    44,    42,    18,   -24,    10,    -4,    -3,    -4,     3,     1,   -30,    -2,    10,    15,     6,     8,    35,    16,     9,     6,     6,   -12,   -10,    40,    75,    60,    43,    59,    54,    40,    25,   -20,     1,     1,    -4,     3,     0,   -25,   -10,   -19,   -35,    15,   -14,    -1,    17,    19,     9,   -31,   -49,    -8,     6,    46,    64,    85,    60,    35,    47,    35,    -9,    12,     4,    12,    -1,     4,    -1,   -10,    -5,   -29,   -54,    19,   -16,   -16,   -21,   -31,   -28,   -38,   -38,     6,     9,     7,    32,    53,    14,     3,     9,   -21,   -20,   -11,     0,     9,    -4,     5,     4,     4,    -4,    -8,   -15,   -34,   -51,   -24,   -56,   -67,   -51,   -46,   -68,   -67,   -53,   -53,   -50,   -41,   -65,   -19,   -11,   -24,     3,     1,     0,     2,     1,     2,     4,    -5,     4,    -8,    -7,    -9,    -8,    -6,    -6,   -25,   -30,   -22,   -26,   -29,   -14,   -15,   -13,    -9,   -11,    -7,    -9,   -11,     2,    -4,     2,     3,     4),
		    93 => (   -1,     0,    -3,     2,    -3,    -4,     2,     2,     3,    -2,     2,    -1,    -3,    -6,     1,    -3,     3,    -3,    -5,     4,     4,     5,     1,    -3,     2,    -4,    -1,     3,     4,    -5,    -1,    -1,     4,     1,    -1,    -2,     4,    -5,    -5,    -2,    -3,    -6,    -8,    -8,   -10,   -12,    -3,    -1,    -5,     1,     1,    -5,     2,     3,    -5,     2,     0,    -5,     0,    -1,    -2,    -5,    -1,     0,   -20,   -25,    29,     7,   -10,   -19,   -32,   -19,   -19,   -13,   -17,   -11,   -34,   -27,   -32,   -19,    -3,    -1,     2,    -5,    -2,    -1,    -2,    -3,     0,    -8,     5,    13,   -18,   -29,   -39,   -31,   -37,   -47,   -59,   -31,   -24,   -30,   -39,   -26,   -25,   -18,   -10,   -25,    -9,    -7,     2,     1,    -4,     1,     3,     1,    10,    28,    33,   -13,    -8,   -39,    -7,    -9,   -11,   -29,   -47,   -44,   -44,   -40,   -38,   -40,   -30,    -9,   -14,   -12,    -9,   -19,     0,     5,     4,    -3,     1,     6,    13,    28,     2,   -10,    -4,    12,    24,    18,    18,    -9,   -15,    -8,   -14,   -12,   -29,   -41,   -26,   -24,   -25,   -10,    -6,   -26,    -9,     5,     2,    -1,     2,    17,     9,   -17,     8,    21,     0,    17,    -9,    13,     6,   -13,   -18,   -22,   -29,   -26,   -18,   -36,   -30,   -23,   -24,   -23,   -18,    -3,   -15,     2,    -2,    10,    -3,    15,     3,    -4,    21,     7,    14,    -4,    -5,   -22,    -2,     3,    -7,    12,   -21,   -30,   -42,   -47,   -29,   -28,   -21,   -24,   -17,    -4,   -12,    -6,     4,     4,   -16,     9,     0,    -2,    -7,   -20,    -6,    -5,   -24,     0,    27,    29,    32,    21,    -6,   -41,   -49,   -51,   -39,   -17,   -21,   -24,   -16,    -9,    -9,     3,    -3,   -13,   -13,     3,    -7,     9,   -16,   -11,   -20,    -7,   -10,    19,    25,    28,    33,     3,   -21,   -57,   -53,   -53,   -35,   -19,   -15,    -7,   -12,   -16,   -13,    -4,    -1,   -22,    -9,    27,     3,    14,     0,   -11,   -19,     1,     3,    12,    20,    17,     4,   -18,   -28,   -59,   -64,   -50,   -41,   -37,   -20,    -1,    -9,   -11,    -6,     0,    -2,   -32,    -1,    34,    20,     4,    -5,    -1,    -7,    10,    15,     9,    15,    -1,   -17,   -20,   -21,   -28,   -23,   -33,   -25,   -35,   -27,   -10,    -2,   -23,   -15,     0,     1,   -25,   -29,    24,    -8,    -2,   -23,   -15,    12,     9,    26,    21,    19,     4,     3,     2,   -21,   -20,     8,     0,    -2,    14,    27,    19,   -19,   -15,   -10,    -4,     1,    -9,   -23,    26,    16,     5,    -2,   -10,    11,    19,    19,    16,    16,    13,     6,   -11,    -3,    -4,     8,    -2,    -7,     8,    15,    24,    23,   -20,   -13,     1,    -5,    10,    -3,    12,   -23,   -15,   -14,   -10,     5,    17,     9,    -4,    -4,     1,   -12,    -4,     7,   -13,    -2,    21,    -3,     3,     3,    43,    16,   -26,   -10,    -6,    -2,    12,     2,     7,   -25,   -21,   -16,    -2,    11,     3,   -10,   -19,   -16,   -16,    -3,   -17,     2,     2,    -1,    15,    28,    19,    17,    16,     4,   -21,    -3,    -1,     4,     4,    -1,     2,   -25,   -39,   -16,   -26,     6,    22,   -18,   -21,   -20,   -36,   -43,   -14,   -18,   -17,    -1,     8,    24,    24,    23,     2,    -4,   -17,   -16,    -8,     4,     1,    -5,    19,    -8,   -19,   -15,   -31,   -13,   -15,   -37,   -20,   -21,   -22,   -40,   -40,   -20,   -21,   -32,    14,    11,    35,    18,    12,    -3,   -14,    -7,    -3,    -4,    -3,     4,     2,     2,   -11,   -25,   -17,    -1,   -12,   -40,   -17,    -8,   -20,   -17,   -32,   -16,    -2,    -7,     2,    12,    17,    12,     1,     6,   -13,    -7,   -16,     5,     0,    -7,   -10,   -13,    -9,   -11,    10,    -3,    -7,   -18,   -11,     5,    11,     4,    -8,     5,    15,    -7,     0,     3,     9,     5,   -11,     8,    -3,   -21,   -11,     5,     1,   -10,   -21,   -15,   -18,   -24,     0,     9,    10,    -8,     6,     7,    12,    17,    18,    24,    -1,   -11,    -7,    14,    14,     5,    -2,    11,    -8,    -6,    -4,    -4,    -2,     0,     2,    12,    -4,   -31,   -23,   -13,    -8,   -15,   -13,   -19,    -8,     4,     1,     3,    -8,   -17,    -2,     0,   -20,    -7,     7,   -11,    -1,   -10,    -2,     1,    -1,     0,    -2,     1,    -4,   -28,   -27,   -27,   -24,   -15,   -21,     0,    -2,   -20,    -7,   -20,   -20,    -8,    -7,    -7,    -8,    -5,     8,   -14,   -10,     2,     3,     3,     2,     7,   -14,    -4,    -6,    -5,     0,   -11,   -11,   -15,     1,    10,    -7,   -14,    -6,   -16,   -12,   -26,   -11,   -13,   -13,   -10,   -21,    -6,    -9,     0,    -1,     3,     1,    10,    -7,   -14,   -11,    11,    16,     9,     0,     1,    36,     6,   -14,    -4,    -7,   -18,   -26,   -16,    -6,   -17,     2,    -5,   -27,   -13,    -9,     2,     1,     4,     1,     2,   -20,    -2,    -8,     3,    10,     4,    -1,    -8,   -10,    -6,    13,     8,    -9,   -16,   -14,     1,    -5,   -35,   -23,   -22,   -31,    -1,    -2,     2,     4,     1,     4,    -1,   -10,    -9,   -12,   -11,   -13,   -25,   -23,    -9,   -21,   -15,     0,   -27,   -11,     2,     1,   -15,   -13,   -13,    -5,   -23,    -3,     4,     1,    -1,     4,     0,    -2,    -2,    -3,     2,    -3,    -3,    -1,    -3,   -11,    -7,   -12,   -12,   -18,   -13,   -24,    -3,     2,     1,   -18,    -9,   -12,    -7,     4,     1,    -1,     5,     2),
		    94 => (   -2,    -5,     2,    -2,     2,     4,     1,    -1,     2,     3,     5,    -3,    -8,    -3,    -9,    -6,    -2,    -3,    -3,    -5,     3,     2,     0,     4,    -3,     1,    -1,    -5,     4,     4,     0,     3,     1,     0,    -9,   -19,    -4,   -18,   -18,   -20,   -21,   -18,    -4,   -25,   -23,   -12,     1,     0,   -21,    -6,    -9,    -2,    -5,    -1,     0,     1,     2,    -2,     2,   -26,   -39,    -9,   -19,   -27,   -15,   -20,   -35,   -55,   -37,   -24,   -35,   -15,    -4,   -12,   -25,   -23,   -25,    -4,   -18,   -16,   -24,   -12,    -5,     0,    -1,    -4,    -1,   -29,   -48,   -11,   -36,   -34,   -18,   -27,   -33,   -15,   -19,   -42,   -28,   -19,    14,   -19,   -28,     0,    -6,     3,     5,    10,   -26,   -18,     2,     5,     4,     3,   -13,   -24,     4,   -14,   -29,     3,     3,   -10,   -29,    -3,    14,   -16,   -14,   -40,   -14,   -22,   -22,    23,    16,    13,    -2,   -15,   -28,     6,    -9,    -1,    -2,     1,   -13,   -27,   -28,   -14,   -20,    -2,     9,     6,    29,    -9,    -8,   -17,   -30,   -39,   -15,     6,    47,     9,     3,     8,   -16,   -17,   -28,    11,   -18,     3,     2,     0,    -5,    -5,   -15,   -15,    -4,     3,    -7,    -5,   -34,   -15,   -17,    -4,   -44,   -70,   -12,     4,    20,    27,    42,    41,   -19,   -12,   -20,   -16,    -5,   -14,     5,   -10,   -20,     0,   -17,    -3,    -6,    26,    -6,   -18,   -27,     5,    19,   -12,   -55,   -49,    -7,    11,    19,    15,    12,    12,   -14,   -15,   -29,   -24,    -9,   -15,   -20,   -23,    19,    -2,   -10,     0,     9,    14,   -16,   -25,   -20,    10,     1,   -22,   -34,   -26,   -25,    40,     5,    14,     1,   -23,   -25,   -33,   -28,   -12,   -23,   -11,    -1,   -21,    14,   -10,   -13,   -18,     3,    -4,   -11,    -8,   -31,    -3,    -9,    -7,   -21,   -35,    -3,    25,    11,    -6,     1,    19,     6,   -26,   -25,    -7,    -6,   -10,    -1,   -15,    17,    24,    -3,   -17,   -24,     2,     4,   -16,    11,     0,    -8,    -4,   -24,   -50,   -12,    17,     5,    -7,   -13,    16,   -19,   -41,   -37,    -6,    -1,    -9,     3,   -32,   -10,    19,   -21,     0,    -6,   -10,    13,    -1,     9,    15,     7,   -12,   -48,   -37,     3,    19,     2,    -3,   -17,   -35,   -33,   -34,   -53,   -21,    -6,   -22,     3,   -16,     8,    -2,   -18,     0,    22,     7,     1,    -4,    23,     9,    13,   -35,   -37,   -36,     1,     4,     6,    -6,   -22,   -30,   -31,     4,    11,     7,   -14,   -21,     1,   -16,    -6,    -6,    -8,     2,    24,     5,     1,     7,    15,    14,    -7,   -33,   -39,   -30,   -12,    10,    13,   -15,   -23,     5,    19,    16,   -16,   -10,   -25,     4,     2,     1,   -29,    -7,    32,    19,     0,    11,    -7,    26,    31,    23,    -4,   -10,   -10,   -22,    -2,     3,     7,     6,     6,    19,    -2,     4,    -8,   -23,   -20,    -1,     1,    -3,    43,    -1,    26,     8,    -6,    -7,     3,     6,    21,    14,    14,     3,   -16,   -25,    -8,    -3,    -6,    14,    -4,    14,    36,   -10,   -32,   -37,   -14,     4,    -1,    -4,     2,   -24,   -13,   -22,     8,     1,   -11,    -4,    -5,   -34,   -20,   -12,   -21,    -8,    -6,     3,     9,    -8,    19,     6,    -3,   -38,   -10,   -19,   -25,   -11,    -3,     4,    11,   -35,     1,    -5,     1,    12,    15,    -6,     0,    -5,   -37,    -5,     1,    13,    -4,     8,    11,   -10,     5,    14,   -19,   -13,   -26,    15,    -4,   -16,   -11,     3,    11,   -20,     7,    15,    11,    20,    -1,    -6,   -11,   -14,   -36,    -7,    10,    24,    -4,     9,     6,    10,    21,     3,   -30,    -6,   -24,   -19,    -8,    -3,     2,    -4,   -21,     2,    -6,     5,    23,     0,     4,     4,    -3,   -41,   -41,   -12,    -6,    26,     4,   -16,    18,    12,    12,    19,   -19,   -14,   -23,   -32,    -1,    -4,    -2,     2,   -11,    -6,     5,   -13,     1,     9,    -1,   -16,   -29,    -7,    -4,     0,     2,     5,     1,    12,    16,    16,    14,    20,   -22,    -7,    -2,   -11,    -2,    -1,    -4,     2,   -25,    -5,     4,    -7,     6,     9,     8,   -23,   -22,   -23,    -5,    -1,    -1,     6,   -11,    15,    10,     4,    15,    19,    16,   -12,    17,    -4,   -15,    -3,     4,     4,    -2,   -26,   -38,    14,     6,    -6,   -25,   -38,   -58,   -27,   -19,     0,    -4,    -8,   -11,   -17,     7,    14,    19,    23,     7,    -8,    -3,    31,     9,    -2,     0,     0,    -2,   -16,   -27,   -20,    -4,   -10,    -5,   -38,   -50,   -27,   -22,   -16,    -4,    -1,    13,   -21,     0,    13,    23,    36,   -21,   -15,     3,     9,     7,    -3,     4,     3,    -3,    -5,   -12,    -3,     0,    -4,   -15,   -24,   -29,   -27,   -14,    -5,   -24,   -13,     2,    -9,     1,    -8,     5,    -6,   -27,    -3,   -23,   -15,   -10,     1,    -3,     4,   -13,    -4,   -14,    -2,    -6,     2,   -11,   -25,   -35,   -13,     1,   -14,   -43,    -1,     6,    -6,   -25,   -46,   -23,   -32,   -39,   -18,   -26,   -19,   -13,     3,     0,    -3,     0,    -5,   -20,     1,    -3,    -6,    -8,   -24,   -43,    -4,   -14,   -28,   -44,   -28,   -46,   -35,   -34,   -32,   -48,   -36,   -40,    -5,    -4,     4,    -2,     3,     4,    -4,     4,     3,    -5,     2,    -5,   -12,    -8,   -14,   -25,   -21,   -20,   -11,   -19,     3,   -27,   -35,   -24,   -18,   -20,   -13,   -22,    -8,     3,     0,     2,    -3),
		    95 => (   -2,     2,     3,    -1,    -2,     2,     4,     0,     4,     5,    -2,    -3,     3,    -2,    -1,     1,    -1,    -4,     0,     2,    -3,    -5,    -3,     2,    -4,     4,     1,    -4,     5,     0,    -3,     2,    -2,     4,    -1,     3,    -2,     4,    -5,    -3,    -1,     2,    -4,    -7,    -9,   -12,    -3,    -2,    -2,    -2,     4,     3,    -2,    -5,     0,     3,    -1,    -1,    -3,     3,     4,    -4,    -7,   -11,   -12,   -19,   -17,   -16,   -21,   -13,    -9,    11,    -3,    -3,    -3,    10,    15,     7,     6,    20,    -6,    -4,     0,    -3,     0,     0,    -9,     5,    -2,    -5,   -20,   -28,    -7,     1,    19,     5,    19,    28,    38,    13,   -10,   -20,    29,    -7,    -7,     9,   -11,   -14,   -15,     4,     8,    -2,     3,    -3,   -12,     1,   -15,   -16,    15,    -1,   -27,    22,     1,    17,    19,   -19,   -20,    -8,     6,   -12,     7,    22,   -18,     6,    20,    24,    43,    41,    12,   -11,     3,     4,    -9,     3,     0,     4,   -12,   -23,     3,    30,    29,     2,   -23,   -26,   -17,    -8,    13,     2,     9,     3,     7,    20,    21,    20,    30,    26,    24,    -9,    -2,    -5,    -5,    -6,    11,     7,   -18,    -7,    27,     5,     9,   -25,   -22,    -4,    10,    28,    11,    25,    18,    -7,     7,    15,    27,    -6,    16,    14,    25,     1,     0,    -1,    -1,   -17,    -2,    -4,   -12,    15,    17,    22,    18,    -2,   -25,   -12,    26,    24,    38,    29,    10,     7,     9,     7,    -9,   -18,   -13,    18,    18,     7,     0,    -3,   -28,   -21,   -24,   -12,    -1,     7,    34,    24,    22,   -16,   -11,   -23,    -5,     7,    -9,     4,     8,   -15,    -6,   -25,   -14,   -14,   -13,   -18,    29,     5,    -3,    -7,   -27,   -26,   -14,    -8,     2,     4,    17,    19,    11,    17,   -35,   -44,   -52,   -62,   -69,   -89,   -49,   -66,   -64,   -60,   -39,   -30,   -28,   -18,    29,    15,     4,    -3,    -9,   -20,    -9,    -3,   -11,     3,    14,    13,     7,    -8,   -33,   -43,   -51,   -37,   -36,   -75,   -82,   -72,   -86,   -82,   -76,   -35,   -19,   -11,     9,    18,    -3,    -2,    -3,    -4,    -2,   -11,    -1,    -5,    11,     7,   -16,    -7,   -11,   -15,     0,    11,    13,     1,   -21,   -23,   -42,   -47,   -55,   -45,   -35,    -8,     1,     5,     0,    -2,     1,    15,     2,    14,    17,     6,    23,     3,    18,     3,   -10,   -12,   -12,     9,    10,     8,     9,    -9,     2,     5,   -21,   -13,   -23,   -18,    -1,     2,    -2,     3,     1,     7,    18,     8,   -13,   -12,    -5,     9,     1,    12,   -11,   -13,   -20,   -21,    -2,    -2,     5,     3,     1,     1,     4,    16,    -6,   -11,   -14,   -23,     1,    -8,    -7,     2,    25,    10,    22,     1,    -5,    15,     0,    -8,    -8,   -22,   -16,     3,    -4,   -17,   -10,   -20,    -3,    -6,    14,     6,    40,   -19,   -26,   -14,     1,     9,    -6,   -33,   -21,   -28,    11,   -23,     0,    -7,    16,    14,    -9,   -12,   -13,   -17,    -8,   -35,   -19,     1,     5,   -11,    -3,    -4,    34,     0,   -21,   -22,    -5,    -5,    -3,   -18,   -35,   -28,   -16,    -8,   -13,     5,    12,     0,    -7,   -19,    -4,    -6,    -5,   -15,   -35,   -15,    -7,     5,     7,     4,    -1,   -19,   -38,   -34,    -3,    -7,   -14,    19,     0,   -18,     9,     4,   -14,    -6,     3,     3,    -2,   -13,   -24,   -33,   -16,   -19,    -8,    12,     8,     8,    10,     3,     3,    -3,   -37,   -35,    -3,     1,    15,    26,   -11,     7,    -7,    -1,    -4,   -23,     2,    -9,   -18,   -28,   -52,   -28,   -23,   -22,    -5,     1,     0,    20,   -16,   -18,    -4,    -2,   -40,   -34,     4,     1,    29,    26,    12,     2,   -13,   -27,   -43,   -24,   -13,   -32,   -15,   -52,   -27,   -35,   -29,     6,     8,    15,    22,    10,     3,   -14,    25,     1,    -7,   -24,    -2,    -3,    15,    19,    19,    -5,   -18,   -16,   -13,    -4,    -9,   -10,   -10,     5,    -9,    13,     5,    18,    12,    11,     0,     5,     1,    -6,   -12,    -4,   -27,     3,    -4,    -3,    -8,     9,    18,    -3,     5,     1,   -18,   -32,     1,    -9,    -6,    -1,   -18,    21,     8,    26,     6,    -7,     0,    13,    16,    25,     9,    27,    -4,     1,    -4,     2,   -19,     8,    -7,     8,     1,    -6,    -8,   -17,   -20,    -7,   -10,    -9,   -16,    18,    19,     5,     5,    -4,     4,     2,     6,    42,     9,    41,    38,    -1,     0,    -5,    14,    14,    -1,     2,    -5,   -11,    16,     4,    -9,    -2,    -6,    -2,     5,   -11,   -11,   -11,   -12,   -17,    21,     6,    21,    19,    12,    29,    47,    -5,    -3,    -3,     1,    19,    26,    13,    20,   -12,    -7,    16,    -7,   -19,    -3,    14,     9,    23,   -20,    -3,    -3,     4,     4,    10,    -8,   -28,    -6,   -11,    -5,     1,    -5,     2,     4,    24,   -21,   -13,    31,    17,    28,    32,    22,    -5,    31,    22,    23,    18,   -16,    -1,    17,    27,    24,    20,    37,    22,    16,    -4,     3,     0,    -4,    -5,    -2,    -2,    -5,    -8,    -7,    -5,     1,     2,     0,     6,     2,    27,    14,     4,   -41,   -18,    -9,     5,   -24,   -15,     5,   -11,    -7,     3,     5,    -3,     2,    -2,     1,     2,     3,    -4,     0,     1,    -4,     4,     1,    -2,    -2,     2,   -10,    -7,    -4,    -1,    -2,    -8,   -19,   -25,   -21,     0,     1,     3,    -2,    -3),
		    96 => (   -2,     3,    -3,     2,    -4,    -1,    -4,    -4,     4,     2,    -3,    -5,    20,    21,    -5,     0,     4,    -4,     0,     4,     2,     1,     2,     2,     2,     4,     3,    -3,     1,     4,    -1,     2,     3,    10,    10,    19,    30,    19,    15,    10,    28,    44,   -14,     9,    19,    26,    25,     7,    22,    11,    11,     7,     3,     2,     3,    -4,    -1,     2,     2,    -2,    28,    31,    21,    22,    12,    14,    23,    33,    51,    36,    19,    17,    22,    25,     8,     1,     6,    -6,    -6,    -7,     8,     6,     4,     1,    -2,     3,    -4,    40,     1,     5,    35,    42,    23,    15,    25,     4,    11,    38,    25,    15,    -7,   -23,   -16,    -3,    10,   -16,    -7,    -7,    -3,    -6,     0,     4,    -2,     1,    -7,    47,     3,    36,    28,     0,    -3,     6,     7,     6,    20,     4,    -1,   -13,   -19,    -5,    -9,   -13,   -40,   -22,   -30,   -31,   -30,   -22,    -3,     7,     0,     1,    -6,    -9,    14,    11,    -2,   -12,   -17,     5,     9,     1,    24,     3,   -32,    -2,   -34,   -11,   -12,   -26,   -44,   -45,   -52,   -36,   -20,   -14,     9,     8,     3,    -5,    -4,   -24,    11,    -7,   -15,   -32,   -28,    25,    11,    18,    14,     2,   -11,   -35,   -25,   -29,   -59,   -59,   -40,   -59,   -54,   -51,   -25,    -7,     4,   -18,    -2,     0,    -3,   -30,    14,     7,   -25,   -34,    -2,    -2,    14,    12,     6,     1,   -20,   -39,   -54,   -56,   -70,   -47,   -33,    -9,   -56,   -56,   -41,   -16,     8,   -23,    -3,     1,     2,   -27,    19,     0,   -12,   -10,    17,    12,     3,    -1,    -9,     0,   -49,   -81,   -58,   -33,   -35,     1,     3,    12,   -17,   -30,   -39,   -35,     3,   -25,     0,    -6,     0,    -8,    21,    -5,   -20,    -6,    12,    -4,    -5,     7,     0,   -54,   -35,   -27,    -8,    -2,    -4,    28,    32,    26,    15,     8,    -1,   -30,   -23,   -12,    -2,    -7,    -2,    -9,    10,     9,   -13,    -1,    13,   -14,     6,    -6,    -8,   -60,   -38,     2,     8,    27,    22,    12,    14,    10,    -5,    -4,     9,   -12,   -31,   -36,     3,     5,    -5,   -16,    18,    15,   -20,     7,     4,    -9,   -11,   -15,   -25,   -52,   -27,    -1,    16,    13,    13,    14,    17,    -1,     0,    -6,     4,     3,   -15,   -19,    -2,     0,   -10,   -28,     6,    -3,    -6,     0,     7,    -6,   -12,   -11,   -28,   -15,    17,   -15,    19,    -8,    13,    18,    18,     9,    20,    20,    23,    11,   -23,   -22,    -2,    -1,   -10,   -27,    -9,    17,     9,   -12,     0,    -6,     5,   -26,   -36,   -10,    -3,    -1,    13,    -1,   -23,    14,     2,    14,    14,    31,    25,     8,   -19,     4,     2,    -1,    -6,   -23,   -16,     7,    23,    -8,    17,    -5,     8,     3,   -18,    -1,     3,    12,     5,     1,    21,   -15,     9,     6,    21,    27,     5,    45,    -5,     1,    -4,     1,    -9,   -16,   -20,    -7,    20,    -3,     2,     4,     0,    -2,    -6,    15,    15,     5,    -6,    -8,     5,   -13,     8,    14,    -5,    -4,     9,    32,    -1,   -29,     1,    -1,   -11,   -22,   -10,     4,    16,     3,    -8,     2,    13,    22,   -13,    -4,    13,     0,     5,    -2,   -25,     7,   -12,    -4,   -13,     5,    22,    31,    -1,   -18,    -4,     2,     4,   -20,   -13,   -11,    -1,    -5,    14,   -14,     0,   -13,    -8,     6,    19,    14,    -9,   -18,   -16,     0,   -27,    -6,   -11,     1,    34,    30,    -3,   -17,     5,     4,    -2,   -21,    12,   -12,   -26,    12,    -1,   -13,   -37,   -22,   -16,    -1,    10,    -6,    -6,     3,    -5,    -7,    -5,    -9,     5,    19,    18,     5,   -11,   -10,     1,    -5,    -1,    -8,    20,   -17,   -13,     6,    10,     1,    -1,   -26,   -25,   -12,    22,    18,    16,    -8,   -27,   -11,     0,    -7,    -8,    -1,     1,    17,   -13,     2,     2,    -5,     1,   -14,    20,     1,   -28,    -7,   -24,    -6,     5,   -18,   -26,   -11,    11,    41,    21,     9,    21,   -13,    15,   -11,   -19,   -22,   -12,    13,     3,     0,     3,    -2,    -4,    -8,     5,    -4,    -2,     9,   -18,    -9,   -12,   -19,   -24,     6,    16,    13,     5,    12,   -15,   -26,     4,   -18,   -10,   -21,   -25,    -3,     6,     3,     4,     1,    -5,    -7,    -9,    -1,     9,   -26,   -45,   -30,   -21,   -37,   -19,     4,    -3,   -15,   -21,   -10,   -18,   -27,   -14,   -38,   -41,   -43,   -45,   -11,     9,     1,     0,    -4,     1,    -6,   -11,    -3,    -5,   -14,   -19,   -37,   -51,   -39,   -29,    -6,    -6,   -34,   -64,   -66,   -56,   -34,    -9,   -31,   -34,   -22,   -38,    -1,    -3,    -3,     3,    -3,    -2,    -1,    -5,    -1,     1,    -8,    -8,    -2,    -2,     8,     1,   -17,   -29,   -28,   -40,   -20,   -32,   -39,   -12,    -9,   -10,     0,    -3,    -4,    -1,     1,     4,     4,    -5,    -2,     2,     0,    -6,   -10,    -9,    -7,    -5,     1,    -4,     0,    -2,    -5,     0,    -2,    -4,   -11,   -28,   -12,   -19,   -16,    -5,     4,    -2,     3,     2,     5,     0,    -3,    -3,     0,     4,    -6,    -5,    -4,    -5,   -13,    -6,    -2,   -10,    -7,    -5,    -5,    -6,     2,    -8,    -2,     2,    -2,     2,     1,    -1,    -3,     1,     0,     2,    -4,    -5,     1,     4,     0,     5,    -4,   -10,    -3,     4,     2,    -2,     1,    -1,    -1,     2,    -4,    -2,     2,     2,     3,    -4,    -4,     0,    -5),
		    97 => (   -1,     2,     4,    -5,     5,    -2,     5,     2,    -3,    -1,     0,     0,    -1,     2,    -5,    -1,     3,     5,     1,     4,     1,    -1,    -5,     3,    -4,     1,    -1,    -1,     2,     3,     1,     4,    -3,    -4,    -5,     4,    -4,    -1,    -3,   -18,   -10,   -11,     3,    -9,   -23,   -33,    -1,    -7,    -1,    -3,    -1,     1,    -4,    -1,    -3,    -2,     5,    -1,    -4,    -5,   -10,    -2,    -4,    -8,    -5,   -19,   -20,   -39,    -6,    -3,    -8,   -16,   -10,     0,    -2,     0,    -9,    -8,   -13,   -14,    -1,    -2,     0,     0,    -1,    -3,     4,    -8,    -3,   -25,   -23,   -51,   -45,   -38,   -45,   -55,   -48,   -55,   -29,   -13,   -11,   -10,     0,   -16,   -22,   -23,   -38,   -10,    -8,   -10,    -3,     1,     2,    -1,    -6,    -7,   -28,   -37,   -39,   -43,   -66,   -69,   -64,   -35,   -36,   -35,   -33,   -22,   -47,   -36,   -25,   -23,   -27,   -15,   -29,   -54,   -54,   -30,   -10,     4,     1,     1,     3,   -34,   -56,    11,   -26,    -9,     7,    11,   -18,   -12,     2,    16,    22,    -4,    21,     8,     1,   -25,   -45,   -28,   -18,   -61,   -42,   -52,   -25,    -1,    -1,    -1,    20,    20,    17,   -15,   -13,   -11,   -15,     2,    -5,     1,    10,     3,     9,    19,    -5,   -12,    -5,     6,    25,    18,    18,   -23,   -41,   -32,   -30,   -19,    -4,    24,    25,     9,    19,   -22,   -10,     5,    -6,    -1,    -9,     7,    11,     6,     9,   -12,   -11,    37,     2,    -9,     2,    -2,    -5,    -9,    -1,   -34,   -44,   -22,   -23,    50,    12,    -4,    12,     0,   -15,     7,    11,    21,    18,    11,     2,    -8,   -13,    -1,    -6,    14,    23,     6,    15,     0,   -13,   -14,   -17,   -50,   -59,   -18,     5,    25,    -8,     5,    15,    12,    14,     4,    16,    31,    29,     5,   -23,   -11,    11,    10,     2,    15,    18,    -1,    20,    -1,    11,   -13,   -23,    -4,    -2,    51,     2,    20,    14,     0,    15,    14,    -4,    17,    28,    14,    15,   -19,   -33,    -9,    15,    33,    16,     0,    12,     8,    23,     0,    -7,   -19,   -19,    13,     1,    44,    -4,     4,    33,     8,   -10,    -3,    -3,     9,    16,    12,   -16,   -17,    13,    25,    45,    29,    20,     0,    16,   -11,     9,   -14,     1,    12,     7,   -37,   -21,    28,     0,    14,    31,     8,   -16,   -14,    -3,    -3,    12,     3,     8,    25,    21,    22,    44,    40,    25,    14,     2,   -23,    -7,    -1,    33,     1,    11,    23,    18,    25,     1,     7,    31,     0,   -25,   -15,     7,    -3,     1,     8,     1,    17,    22,    15,    51,    32,    22,     9,   -21,   -19,   -35,   -12,     5,   -10,     2,    23,    -7,   -20,    -6,    12,    13,   -21,   -32,    -3,    -6,   -18,    -2,     4,   -11,     7,     3,     7,    29,     6,     8,    13,   -10,   -10,   -16,   -30,    -9,     6,    20,   -21,   -26,    -1,    -3,    -1,     7,   -20,   -25,    -5,     3,    -9,   -35,   -31,   -13,    -8,   -13,     2,    -8,   -15,     0,    12,    29,    -6,     5,     4,    27,    19,    18,     8,   -11,   -15,     1,    -7,    -2,   -16,    -8,    -2,     1,    -5,     0,    20,    14,   -13,   -32,   -18,   -16,    -6,   -10,    35,    53,    41,    11,    34,    21,    32,    24,   -22,   -21,   -18,     2,    -7,    -6,   -10,     0,     4,     1,   -17,    -1,    -1,     0,   -22,   -38,   -13,     1,     1,    25,    36,    46,     9,    25,    16,    31,    26,     3,    16,    -6,   -27,     6,     2,    10,   -10,    -2,    18,    17,   -10,   -17,   -22,   -10,   -19,   -21,   -14,    -9,     3,     7,    52,    29,    16,     8,     5,    18,     7,     2,     6,     2,   -18,    -5,    10,     3,    -3,     7,    11,    11,     5,    11,   -20,   -11,   -11,   -19,   -27,   -12,   -14,    29,    54,    19,    17,     3,     9,     3,    -2,    15,    -5,   -20,    -6,     2,    12,    -5,   -13,   -33,     6,     2,    12,    10,     3,    -7,    -8,   -13,     0,     0,    10,     2,    11,    -3,    -2,    -2,    -2,   -13,   -12,    13,   -13,   -23,     3,    -1,     2,    -4,   -11,   -22,    18,    16,    18,    11,    22,    20,     3,     6,     5,    -9,    11,     3,   -17,   -25,   -19,   -11,     8,   -10,    -7,   -22,   -18,    -6,     3,    -2,    -2,   -13,   -22,   -24,    11,    31,    14,     3,     3,    10,    -6,    10,     7,    -6,   -22,    -2,   -27,   -21,   -23,   -26,   -19,   -36,   -35,   -22,     3,   -23,    -4,    -4,     5,   -10,   -40,   -20,    16,    29,    19,    10,    -2,    22,    -1,    -8,    -1,   -39,   -32,   -14,   -30,   -36,   -30,   -20,   -20,   -42,   -38,   -13,     3,   -18,     3,     0,     2,     0,    -6,    -2,    21,    10,    18,    -1,     1,     0,     6,    -3,     1,   -23,   -27,   -18,   -15,   -42,   -38,   -32,    -9,   -35,   -39,   -22,   -19,    -3,     4,    -3,    -4,   -13,    24,    -2,    -1,     2,     6,   -17,    10,     9,    -5,    -7,     5,   -36,   -31,     2,   -23,   -30,   -42,   -26,    -7,    -2,   -27,   -11,    -5,    -3,    -1,    -4,    -2,    -3,   -26,   -18,   -25,   -14,   -13,     4,    28,    -4,    -8,    -2,    -2,     2,     5,    -7,   -25,    -6,    -6,     0,    11,    -2,    -1,    -4,     0,     4,     2,    -1,     5,    -4,     1,    11,    14,     0,   -13,    -9,     0,    -1,   -20,    -6,   -12,   -22,     6,     2,    28,    11,   -12,     0,    15,    -2,    19,    -3,     0,    -2,    -4),
		    98 => (    3,    -3,    -3,    -1,     3,    -2,     1,     5,     1,    -1,     2,    -3,     3,    -4,     0,    -5,    -5,    -2,     2,     3,     1,    -4,    -2,    -2,    -1,     1,     0,     0,     1,     4,     2,     5,    -4,     1,     5,     3,     2,     3,     0,     3,    -4,    -7,    -7,   -18,   -17,   -18,    -7,     5,    -6,    -4,     0,    -5,    -2,    -3,    -3,     3,     2,     5,    -5,    -1,     0,    -1,     3,    -2,   -10,   -28,   -39,   -36,   -13,    -2,    -8,   -25,   -25,    -9,    -4,     1,    -6,    -9,   -14,   -10,     0,     0,     0,     1,     4,     5,    -6,    -3,    -6,   -15,   -11,   -48,    16,    23,    30,    12,    29,    34,    22,    12,     3,    11,    -9,   -22,   -18,   -29,   -17,    -2,    -6,    -8,    -5,    -2,     1,    -6,     4,    -5,   -31,   -35,    -7,     8,    10,    14,    -9,   -22,     3,    -9,    -5,    -8,    -4,     2,    -4,     9,     1,     8,   -31,   -17,    -7,    -1,     2,    -7,    -1,    -3,    -1,   -25,   -31,   -54,   -16,    10,    13,   -13,    -1,     5,   -28,   -16,    13,    -3,     6,    19,    11,     1,    15,    -1,   -12,   -19,   -16,    -6,     7,    -5,     4,    -2,   -29,   -14,   -12,   -16,     1,    42,    22,    13,    14,     6,     2,     7,    10,    17,    12,     1,   -16,    14,   -12,    -4,   -16,    -5,   -15,   -13,     1,    -2,    -4,   -19,   -11,   -24,    -8,    -2,    24,    35,   -20,    -8,     8,   -16,    -5,   -17,   -12,   -12,   -17,    -4,     1,     9,    -6,   -23,   -12,   -19,    -8,   -10,    -6,    -7,    -6,   -11,   -20,   -13,   -31,   -29,     9,    36,   -13,    -9,    19,    11,   -12,   -24,   -25,   -11,   -38,     5,     0,     5,    -7,   -10,    -5,   -25,     1,    10,    12,    -2,     3,    -3,    -8,    -6,   -38,   -29,    -5,   -11,   -13,     3,    23,    27,    12,   -14,   -18,   -10,    -4,    18,   -21,    -4,     1,    12,    -5,   -12,    -7,     5,   -32,   -30,     3,    -8,   -15,   -16,   -18,   -37,    10,   -17,   -47,   -10,    14,    50,    47,    31,    11,    -4,     3,     7,     7,   -25,    22,    12,     3,   -20,   -34,   -40,   -33,   -33,    -1,    -5,    -5,   -22,   -14,   -14,     2,    -4,   -18,    -3,   -36,     2,    24,    39,    28,     0,    -9,   -21,    -7,    -8,    -6,    -6,   -16,   -16,   -37,   -27,    -8,   -12,     1,     2,    -9,    -5,    -8,   -19,   -10,   -27,   -40,   -41,   -48,   -47,     3,     3,    10,    31,     7,    -2,    10,    11,     3,     8,     7,    -3,    -5,   -21,   -15,   -11,    -4,    -2,   -10,    -3,   -13,    -7,    -4,   -23,   -39,   -55,   -43,   -32,   -25,    -2,    -1,    19,     8,    -8,    -3,   -13,   -26,     1,     8,   -28,   -26,   -20,   -18,    -5,    -3,    -3,     1,   -24,   -14,     5,    -1,   -15,   -20,   -29,    -5,    13,     6,     5,    -5,   -16,     0,     3,     1,   -22,   -11,    13,    -8,   -28,   -28,   -16,   -32,   -16,    -5,     4,   -15,   -18,   -23,   -11,   -15,     1,    -7,     5,     0,    11,    -6,   -20,   -13,    -6,    15,   -10,   -20,     2,    -1,    12,   -24,   -18,   -19,   -17,   -36,   -13,    -1,    -5,   -10,    -9,   -18,    -2,    18,    14,     4,    25,     5,     1,   -20,    -5,   -31,     1,   -31,    21,   -16,    19,    19,     9,   -12,    -6,   -11,    -9,   -44,   -17,     4,    -2,   -14,   -34,    10,     4,   -10,    18,    16,     3,   -12,    -3,    -9,   -37,   -33,    -9,   -24,    -8,     8,    24,     6,    28,    22,     0,   -18,   -15,    -8,   -21,    -5,    -3,    -7,   -12,    31,     0,     9,    22,    -5,   -20,   -13,     7,   -14,   -34,   -14,   -12,   -43,   -15,     9,    15,    14,    13,    11,     8,   -29,   -16,    -1,   -13,    -1,   -10,   -19,    21,    23,    30,    23,    10,   -23,   -13,     3,     8,   -33,   -20,   -23,    -6,   -14,    -2,   -12,     0,     8,    13,     2,   -18,   -26,   -11,   -38,   -13,    -4,    -2,   -16,     4,    20,    11,    15,    10,    -9,   -29,    -6,     5,   -24,    -5,    -4,     6,    14,   -13,   -14,   -10,    16,    13,     7,   -16,   -14,    -3,   -33,    -5,   -13,    -7,   -19,   -19,     5,    -2,     2,    -3,   -15,     1,   -12,    -2,     5,   -13,    14,    -9,   -10,   -19,   -31,     6,    14,    18,    -5,   -13,   -19,   -11,   -28,    -5,   -13,    -9,   -17,   -22,   -19,     3,    28,    21,   -17,   -11,     5,     8,    14,   -20,    -5,   -25,   -16,    -8,   -15,    -8,     4,   -10,   -29,   -10,     2,    -3,   -18,    -2,    -4,     4,    -5,    -9,   -28,    18,     5,    22,     6,   -19,   -10,   -18,     4,    -3,    -1,    -8,   -10,   -21,    -8,    -2,   -14,   -38,   -17,    -7,     2,    14,   -26,    -3,    -5,    -3,   -11,    -7,   -22,   -23,    11,     9,     6,    -1,   -18,   -15,    -3,     1,    12,    15,    24,   -15,     3,    -2,    -1,   -15,   -15,    -4,   -21,    -3,    -7,    -2,     1,     3,    -3,    -2,    -5,   -15,     0,    -9,   -22,   -15,   -24,   -27,   -23,   -28,   -27,   -30,   -22,   -14,    -6,    -1,     0,   -12,    -5,    -5,    -6,    -2,    -5,     4,    -2,    -5,    -3,   -10,    -8,    -5,    -3,    -6,    -7,    -7,    -9,    -5,   -20,   -23,   -29,   -16,   -13,   -10,    -9,   -19,   -32,   -32,   -18,     2,     0,    -4,     5,    -1,    -4,    -2,     4,     0,    -8,    -6,   -10,    -5,    -6,    -7,    -3,    -4,     0,   -18,    -6,    -4,    -7,    -8,    -8,    -6,     2,    -3,     4,    -3,    -2,    -3,    -4,     1),
		    99 => (    1,     3,    -1,    -1,    -5,    -4,    -4,    -4,    -4,    -4,    -1,    -2,     1,    -3,     2,     1,    -1,    -3,     4,     2,     0,     5,    -2,    -5,    -3,     2,     1,    -3,    -4,     0,    -5,     2,     2,     4,     3,     1,    -2,    -2,    -8,   -10,   -14,   -14,     3,    -4,     2,    -3,    -7,     0,     0,    -2,    -7,    -3,    -1,    -1,     2,    -2,     0,     3,    -3,    -4,    -3,     2,    -2,    -4,    -1,    -6,     0,    -8,     0,     3,   -11,     2,     2,     2,    -4,     1,    -7,    -8,   -10,    -2,     1,     1,    -5,    -1,     3,     0,     1,   -11,    -5,    -8,    -7,    -5,   -17,   -14,    -8,    -1,     4,    -6,    -6,     1,    -3,    -7,    -8,    -9,   -17,    -4,   -15,    -9,   -17,   -11,    -2,    -5,     0,     1,    -2,    -5,    -7,    -7,   -26,    -2,     2,     1,     1,    -7,   -21,   -20,   -10,   -22,   -13,   -22,   -11,   -27,   -38,    -4,    -4,    -2,     2,   -24,    -8,    -3,     4,     3,    -4,   -10,    -3,     2,    -1,    -7,    -7,   -11,    -6,   -16,   -21,   -27,   -32,   -38,   -23,    -7,    -4,    11,   -15,   -12,   -13,    -6,    -3,    -7,   -11,     3,    -3,     3,    -2,   -11,    -3,   -11,   -16,   -14,   -24,    -7,   -14,    -1,    -4,    -3,    -1,     1,   -14,   -26,    -9,   -16,   -20,   -15,   -15,    -9,    -6,    -1,    -9,   -13,     2,    -3,    -6,   -10,    -9,   -16,   -29,   -37,   -37,   -19,   -14,     5,     0,    12,     3,     7,    12,   -19,    -7,   -19,   -17,   -31,   -16,    11,   -11,    -3,    -4,    -9,   -18,   -15,    -7,   -10,   -20,   -25,   -29,   -40,   -26,   -21,     1,     5,     6,    -8,     3,     1,    19,   -18,    -7,     6,    -4,    -1,   -18,     0,    -3,   -22,    -5,     0,     0,   -18,   -14,   -18,   -23,   -15,   -27,    -8,     4,    -9,     2,     8,    11,     7,     8,    31,     8,   -10,     4,    20,     4,     0,     0,    -4,   -10,   -16,   -10,    -9,    -5,   -22,   -15,     0,   -12,   -17,   -24,   -11,     5,   -17,   -24,    11,    12,     7,    20,     3,    14,   -10,    20,    15,    -5,     2,    -5,   -18,   -17,   -17,    -7,   -13,    -1,   -40,    26,     1,    -7,   -10,   -12,    -1,     0,   -11,   -30,     1,     6,    16,    10,    -2,   -15,   -20,    -1,     3,     3,    -6,     0,   -10,   -26,   -24,    -5,    -8,    -1,   -18,     9,    22,    19,     2,    10,     0,   -13,   -39,   -26,    -4,    -8,   -12,     2,    -1,    -7,    -1,    -5,    10,     0,    14,    -3,    -5,   -25,   -13,   -19,    -2,     3,   -20,    -7,    13,    12,     6,    12,    -3,   -14,   -47,   -13,    -6,   -33,   -31,   -19,     4,    -1,   -18,     4,     3,   -10,    18,     5,   -11,   -30,   -18,    -9,     1,    -2,   -13,   -17,    16,    14,    14,    -2,    -4,   -32,   -28,    -9,    -6,   -21,   -23,   -26,    -6,    -7,   -16,    -1,     4,    11,    12,    -8,   -22,   -25,   -14,     1,    -1,    -3,     2,   -24,    15,    23,     6,     7,     0,   -19,   -33,    -7,   -16,   -21,    -4,    -3,     2,     0,   -28,     3,    -4,    -5,     9,     9,   -24,   -29,   -16,     1,    -9,     2,    -7,   -15,    15,    29,    19,    34,    11,     4,     7,     5,   -20,     3,     1,     3,     0,   -30,   -20,   -14,   -20,     1,    -4,    20,    13,   -24,    -3,   -13,    -4,     1,    -5,   -39,    -3,    -3,    -1,    12,    19,    28,    21,    17,    24,    15,    -3,    -6,   -18,   -23,   -26,    -4,   -14,   -10,    -4,    17,    -6,   -24,    -9,   -17,   -16,    -4,     1,   -38,    11,   -11,   -19,    -4,     9,    -2,    -4,    24,     5,    -2,   -29,    -8,     0,    -9,    -8,    -2,   -25,    -4,   -10,    15,    14,   -11,    -3,   -21,   -11,    -4,    -6,   -21,    16,     1,   -22,   -19,   -13,   -28,   -24,    -9,    -9,     2,   -31,     9,     0,   -14,   -14,   -10,   -32,     1,   -19,    -5,    19,    22,    15,   -18,    -3,    -5,     0,    -8,    16,    12,    -4,   -15,   -19,   -28,   -17,   -23,   -13,   -36,   -26,    11,     9,   -15,   -27,   -10,   -15,     5,    -1,    -6,    19,    22,    40,   -20,    -4,     1,     4,   -14,     6,     7,    -4,   -12,   -13,   -16,   -26,   -17,    -6,    -5,   -17,    15,   -12,   -50,   -14,    -5,   -10,    -7,    15,   -16,     1,    10,    24,   -25,    -3,    -2,     4,   -16,   -12,   -21,    -8,   -11,   -18,   -10,   -16,    -9,   -16,    -3,    -3,    25,   -29,   -33,    -4,    -1,    -9,     0,     2,    -4,     4,    -9,   -23,    -6,    -2,     1,    -1,   -13,   -12,   -12,    -4,    -6,    -9,    -9,    -3,   -12,    -3,     0,     1,     8,   -14,     4,     9,    -2,   -10,    19,    -1,    25,    10,    -1,   -10,    -6,    -2,     2,    -4,   -11,    -3,   -17,    -9,     1,     7,   -19,   -20,   -11,    -6,     2,    -5,     7,     8,    15,    -9,    -3,    -3,    17,    11,    15,    10,     2,    -5,    -5,     3,     0,    -4,    27,   -19,     0,    14,     5,     0,   -25,   -10,    -9,    -1,    -8,   -18,    15,    12,     7,    -4,    -8,    10,    20,    13,    15,     2,    -8,    -6,    -3,    -4,     0,     2,     4,    29,    15,    13,    13,    -2,     3,    17,   -14,    -5,    -7,   -22,     1,     7,    -3,    -4,    -2,    13,    21,    32,    17,     1,     8,     3,     5,    -2,    -1,    -2,    -4,     0,   -10,    -6,     9,    21,    17,    15,     0,     4,    -6,   -16,    -3,    -6,    -5,    -3,   -13,    -9,    -7,    -4,    10,   -11,     5,    -4,     0,     0)
        );

 ---------------------------------INFO-
 -- COEF =43.138084

 -- MIN =-127.99999
 -- MAX =84.78604

 -- SUMMIN =-9094.42
 -- SUMMAX =6612.154
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
