----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (   -3,     0,    -1,    -5,    -6,     8,     1,     0,     5,    -6,    -2,     9,    -1,   -16,   -14,     3,    -9,     7,     4,     2,   -10,    -8,    -4,     6,    10,    10,    -2,    -9,    -7,    -7,    -1,     3,     2,    -8,     6,     3,    -1,     1,    -5,     7,    13,     9,   -14,     9,    27,    11,    -4,    -8,    -9,     7,    -2,     3,     3,    -1,     4,    -8,     6,    10,     1,    10,    26,     2,   -14,     1,   -16,   -43,    -5,    -8,    -4,   -25,   -23,   -37,    -5,    -8,   -15,    -6,    -6,    -6,   -22,   -17,   -15,   -18,     2,    -6,     4,    -9,    -3,    20,    -2,    14,    10,   -31,   -21,   -17,   -28,   -21,   -38,   -25,   -37,   -40,   -12,    26,     1,   -32,   -23,   -16,   -23,   -14,     9,     6,    -6,     6,    -6,     5,     2,    -3,   -14,   -35,     7,   -24,   -53,   -26,   -26,   -41,   -67,    -6,    -2,   -19,    -8,   -36,   -26,   -22,    -4,   -13,   -20,   -14,     5,   -10,   -19,     3,     2,     7,   -19,    -5,    -1,   -13,    -9,    -4,   -15,   -10,   -33,   -60,   -37,   -52,     8,    24,    -2,   -24,     2,   -34,   -43,     2,    -7,    -6,   -11,   -45,   -13,   -10,    -9,     9,   -20,   -14,   -13,    -1,   -11,   -10,   -20,   -20,   -18,   -64,   -46,   -19,    -6,   -21,    27,    19,     4,   -39,   -35,   -21,     5,   -44,   -19,   -41,   -11,    25,     1,   -19,   -17,   -17,     5,    -8,   -12,     7,   -15,   -18,   -42,   -66,   -64,   -23,    -2,     1,    43,    23,   -40,    -1,   -37,   -32,    13,   -23,   -37,   -14,   -40,    26,    31,   -52,    27,    18,    -6,    -9,   -12,    -2,    -7,   -35,   -22,   -63,   -13,   -12,    15,   -22,    10,    47,   -20,     8,   -41,   -50,   -11,   -28,   -15,   -51,   -18,   -13,   -12,    -9,    47,    -5,    -4,    -5,   -32,    -5,   -24,   -60,   -24,    -7,   -13,    16,   -11,   -16,    31,     8,     1,   -31,   -76,    -7,    -5,   -18,   -23,   -41,     1,     8,   -11,    -9,    11,    19,   -19,   -25,   -11,    16,    -1,    -6,   -20,   -13,    -9,    -3,   -47,   -50,   -17,   -35,    10,   -33,   -34,   -13,   -30,   -37,   -16,   -13,   -36,     4,     5,    45,   -19,     9,   -25,    -4,    -8,    -4,   -16,   -12,   -30,     3,    19,   -16,   -18,     4,   -26,     8,    60,   -43,   -34,     6,   -31,   -49,   -18,   -28,   -19,    -8,    -4,    14,     8,     0,    -2,     9,     3,    -1,   -49,    -1,     6,   -11,    23,   -10,   -20,   -51,     6,    29,    50,   -10,     2,    31,     0,   -51,   -33,   -32,   -26,     7,    -2,    22,    23,   -10,    -1,     5,    22,   -29,   -27,     3,   -10,   -37,    13,   -35,   -92,   -73,    -6,    25,    44,    13,    -7,    34,   -16,   -29,   -23,   -13,   -40,     2,    -4,    -1,     1,   -13,    -9,    18,   -22,   -30,   -25,    -6,    11,    17,    40,    -6,   -63,   -67,    -3,     8,    20,    15,   -36,     2,    -4,   -18,   -25,     7,   -32,    -2,     1,    -8,   -19,   -16,     8,   -33,    -1,   -50,   -25,   -41,    -9,    17,    54,    11,   -83,   -27,    -9,    11,    -5,   -13,   -37,    30,   -28,   -22,     3,   -21,   -25,    -4,    -8,     2,    -9,   -25,     7,     2,   -58,   -17,   -37,   -44,   -24,    24,    25,   -27,  -100,    -3,   -10,    66,   -19,   -11,   -28,   -24,     0,   -24,   -26,   -19,   -56,    24,     0,     4,   -34,   -17,   -44,   -13,   -29,   -28,   -32,   -79,     9,    12,    32,   -23,   -73,   -26,    -1,    33,    12,     0,    18,   -23,   -11,    13,   -23,   -30,   -55,    20,     1,     4,   -15,    11,   -15,   -25,   -11,    -6,   -25,   -41,    29,    29,   -26,   -41,   -83,    -9,    -4,     4,   -12,     2,     0,    -8,    10,   -20,    -1,    -4,   -25,   -13,     8,    18,     4,    12,     5,   -22,   -10,   -41,   -30,     9,    22,    26,     0,   -45,   -47,    33,    10,   -27,   -21,     0,   -38,   -16,   -17,   -15,     3,   -72,   -14,    -9,    -4,     1,    -9,   -18,     8,    -9,   -26,   -50,   -41,    12,     4,   -27,   -31,    -9,   -10,     8,    12,   -25,    -1,   -44,   -27,   -32,    -9,    -7,   -11,   -14,     7,    10,     2,    -4,   -23,   -26,   -11,   -13,     2,   -32,   -19,   -12,     9,   -11,     0,    -8,    -8,    20,   -10,   -10,   -27,   -39,   -39,   -21,     7,     3,   -37,     3,    15,    14,    -2,     4,   -19,   -58,     6,     3,    12,     3,   -19,    13,     6,    20,    -7,   -43,    33,    27,    30,   -60,   -25,   -32,   -28,   -20,     6,    -8,    -2,   -10,    14,     5,     3,     4,   -22,   -43,   -19,     8,   -16,    -4,   -19,   -43,    25,    14,    20,    27,   -30,   -28,   -33,   -71,     0,   -43,   -28,   -14,    20,    -3,   -16,   -40,   -22,    -8,     9,    -9,   -10,     2,   -25,    26,    12,     8,   -44,   -51,   -32,   -34,     6,    51,    11,     9,   -45,   -16,   -10,   -33,   -30,    17,   -19,   -24,    -2,    -6,    -9,     4,     2,     8,     3,    -7,   -72,   -28,   -27,   -25,   -12,   -26,   -43,   -49,   -73,   -68,   -84,   -35,   -21,   -25,   -27,   -20,   -36,   -14,   -24,   -18,    -2,     2,    -4,    -1,     1,     6,    -8,    -4,    -7,   -34,   -52,     5,    -3,   -33,   -18,    -9,   -27,   -21,   -25,   -24,   -13,   -37,   -55,   -23,   -39,   -24,   -10,     0,    -9,    -6,    -7,     1,     4,   -10,    -2,    -9,    -2,     6,     3,    -3,    -5,   -10,     6,    -4,     5,   -24,     6,     0,   -15,     1,     9,     2,    -6,   -13,   -13,   -20,    -4,     1,   -10,     7),
		     1 => (   -2,    -5,    -3,    10,     2,    -4,     1,    -3,     8,    -8,     3,    -7,    -5,    -9,     4,     7,     1,     4,    -7,     4,   -10,    -5,     9,    -5,    -1,     4,    -8,     7,    10,    10,     9,     8,   -10,     9,     2,     4,   -10,    -5,    -5,    -9,   -16,   -10,    33,    25,    -1,   -16,   -10,     7,    -9,    -8,    -1,    -5,    -7,     7,    -5,     9,     6,     2,    -1,     8,     3,    -3,     8,     5,   -28,   -28,     1,    -8,    -8,    -9,   -16,   -34,   -39,   -45,   -57,     6,    18,   -50,   -15,    -3,    -9,   -14,     4,     9,     7,    -8,    61,    43,    -3,     7,     9,    49,    40,    26,    27,    14,     6,   -75,   -77,   -77,   -66,   -18,   -20,    -6,     8,   -39,    18,     3,   -27,    -3,     6,     7,    -1,    -2,    41,    35,    19,   -11,    -8,     1,    -1,    -8,   -29,   -70,   -68,   -83,     8,    34,     3,     7,    12,    17,    10,    17,   -20,   -83,   -43,   -70,   -41,   -39,     2,   -10,    41,    56,    18,     4,   -19,   -20,   -96,   -42,   -35,   -61,   -81,   -46,    -6,    57,    -4,    -6,    -2,    21,    23,   -24,   -35,   -80,   -59,   -43,   -42,   -34,    -3,    -4,    -1,    22,    19,   -17,    -2,     8,   -78,     5,     7,   -60,   -62,   -31,   -45,   -17,    -4,    19,    -2,    23,   -23,   -26,   -14,   -83,   -58,   -23,    -3,   -13,    -7,    -2,   -18,    18,    10,     2,   -17,   -32,   -86,   -19,   -45,   -70,   -52,    -9,    33,    15,    16,    -6,    39,    -9,   -31,   -22,    -1,   -53,   -57,   -23,   -25,   -18,     0,   -13,   -13,   -12,    -8,   -12,   -28,   -31,   -61,   -53,   -26,   -98,   -90,     2,    23,    18,    34,    21,    12,   -20,   -34,   -17,   -29,   -50,   -58,   -31,   -32,    -6,     7,    -2,   -13,    15,   -12,     1,   -46,   -23,   -17,   -28,   -69,  -129,   -31,    -7,   -16,     1,    41,     7,   -41,   -27,   -58,   -23,   -14,   -31,   -54,   -28,     2,   -31,     1,    12,    -6,   -13,    -5,    -5,   -40,   -52,   -34,   -46,    -7,   -65,   -51,   -25,     9,    47,    40,    -6,   -40,   -36,   -53,   -20,   -19,   -25,   -56,   -62,    -3,    66,     2,    -1,    10,    17,    19,     4,   -26,   -31,   -51,   -84,   -44,   -71,   -20,   -29,    -1,    59,     4,   -53,   -30,   -17,   -19,     9,   -16,   -34,   -62,   -57,    -3,    57,     2,     2,   -19,    45,    11,   -12,   -16,   -12,   -81,   -69,   -39,   -38,     3,   -18,    40,    -8,    23,   -82,   -88,   -30,    39,    53,    53,    36,   -15,     1,    -8,    34,     3,    -9,    -2,    13,    22,   -16,   -20,    -7,   -40,   -92,   -41,   -21,   -14,    11,    46,   -19,    16,   -76,   -87,     7,    35,     4,    -4,   -67,   -38,     3,    19,     6,    -7,     7,    21,    21,    26,   -49,   -30,   -20,   -10,   -58,   -40,    15,    -7,   -32,    46,     2,   -35,   -75,    -5,    46,    52,    65,    37,   -19,   -30,    63,    60,     1,     7,     3,    24,    58,    24,    -6,   -14,    -6,    34,     4,   -14,    35,     2,   -20,   -17,   -48,   -36,   -60,   -22,   -49,    -7,    69,    28,   -36,   -82,    20,    12,    -7,     5,     9,     7,   -25,   -19,    -5,    13,     3,    35,    22,    18,    40,    17,    18,   -32,   -15,   -13,   -71,   -60,   -64,    -7,    52,    34,    64,    79,   -20,   -14,    -4,     6,    -5,    12,   -29,    10,     4,    31,    11,    24,     8,    10,    17,    -6,    13,    13,   -17,   -31,   -24,    14,    28,    36,    61,    67,    75,    46,    -3,   -12,   -27,   -23,    -5,    -2,   -18,   -19,   -25,   -29,   -13,    11,   -32,     9,   -15,    -6,    24,   -36,   -77,   -59,    14,    39,    44,    27,     5,     5,    -2,    21,    41,     6,    29,    -4,    -9,    33,    32,   -38,    31,    38,    11,     3,   -33,    -7,    18,    16,    21,   -46,   -56,   -85,   -14,    26,    -7,    -7,   -14,   -44,     4,    42,    54,    11,    27,    -2,    -6,    33,    11,     0,    54,    22,   -34,    -1,   -13,   -37,    14,    -2,    21,   -24,   -64,   -72,   -18,   -19,    -7,    41,   -45,   -26,     1,    21,    19,    23,    -1,    41,    27,   -12,    -3,     1,   -45,   -72,   -24,     3,   -15,     3,   -13,    20,   -30,    -1,   -16,   -62,   -65,   -54,   -19,    24,    15,    14,    19,    28,    28,     6,     5,    31,    35,     5,    -1,     4,   -38,   -86,   -16,    -3,   -22,    16,   -23,    -6,   -10,    25,   -28,   -21,   -53,     5,    38,    61,    22,    39,    28,    35,    52,    82,    10,    -8,    -8,   -10,     3,   -29,    -6,   -28,   -35,    34,   -21,    -9,    20,    -1,     5,    17,    -7,    10,    10,    18,    49,    60,     4,    -5,   -13,    25,    40,    79,    -5,     0,     3,    -7,   -11,   -25,   -45,   -13,   -39,   -23,   -39,   -68,   -20,   -32,   -77,    28,    25,   -10,    11,     8,   100,    67,    11,    -6,    10,   -17,    13,    20,    -2,     6,     7,    -1,    -3,     1,    -4,    -7,   -10,   -33,    20,   -67,   -36,   -53,   -44,   -46,   -73,   -28,   -43,   -28,   -31,   -39,   -34,   -21,   -17,   -13,     3,   -10,     8,    -4,    -7,    -4,    -7,   -17,   -34,   -43,   -21,   -26,   -33,    13,    -6,   -53,   -50,   -67,   -70,   -55,   -38,    -9,   -19,   -10,    -9,    -2,     5,   -10,     5,    -8,     2,    -4,    -2,   -10,     6,     9,     3,    -5,    -5,    -6,    -8,   -10,   -14,     7,     6,    13,    -3,    -6,    -3,   -10,    -9,    -1,     5,    -7,     8,     9,     2,     5,     7),
		     2 => (    0,    -8,     4,    -9,    -8,     4,     6,     4,    -1,     7,     2,    -9,    -1,     2,     1,     4,     2,   -10,    -3,     1,     1,     5,    -1,     4,     2,    -7,    -3,    -5,    -1,     5,     0,    -2,     8,     6,    -7,     8,   -20,   -29,   -19,   -16,    -9,   -44,   -32,   -11,    -2,    11,    -2,    -9,   -12,    -7,    -7,   -18,     4,     5,     9,     7,     3,    -8,     2,   -26,   -30,     1,     7,   -52,   -13,   -22,   -22,   -37,   -20,   -99,   -29,    -5,   -15,   -23,   -42,   -51,   -39,    -8,   -23,     4,    12,    22,     6,     8,    -4,     8,   -15,   -41,   -39,    -1,    44,   -18,    -6,    41,    43,     6,   -43,   -55,   -32,   -56,   -52,   -19,    27,   -17,   -58,   -34,    -6,   -22,   -28,    13,    -7,    -9,    -8,    10,    -3,    24,   -14,   -27,    -5,    43,     9,    -4,   -42,   -31,   -27,   -63,   -65,   -42,    16,    16,     4,   -21,    22,    31,    -8,   -48,     7,     6,   -26,   -10,     0,     8,   -14,     7,    52,    11,    -2,    -2,    -9,   -17,   -48,   -67,   -72,   -69,   -54,   -26,   -10,     6,    32,    35,    25,    42,    10,   -36,   -30,     3,   -28,    -6,     9,    10,    17,     5,     9,   -11,   -14,    25,    13,   -17,   -17,   -27,   -12,   -70,   -54,   -46,   -27,    42,    16,    29,   -11,    12,     7,   -57,   -49,    48,   -29,    -5,     5,     7,    42,     2,    -2,   -26,    -4,    28,    -3,    10,     0,    20,    14,    30,   -25,   -26,   -21,   -17,   -53,   -13,    18,    12,     5,   -94,   -11,    68,   -34,    -5,   -53,    48,    45,   -29,   -19,    17,    -2,   -16,   -27,   -54,     5,    36,     1,    16,    22,   -64,   -81,   -29,   -34,     8,    22,    -8,    -4,    10,    11,    34,   -50,   -12,     1,   -23,    50,   -24,   -44,    -9,   -10,     1,   -34,   -24,    16,   -19,   -32,     4,    16,    10,   -25,   -21,    -8,    40,    12,    19,    15,    -9,    -9,   -48,    35,   -17,    -9,   -18,    42,   -53,   -28,    27,    25,    36,    -4,    -1,    12,     3,    23,    52,    96,    30,   -35,   -19,     5,    45,    15,    22,     8,   -44,   -24,   -35,    23,   -26,     7,   -39,   -28,   -36,    25,     7,    24,    51,    45,    25,   -26,   -20,   -54,   -18,     4,     3,     0,   -45,    -4,    27,    -1,    13,     9,   -45,    -1,   -14,    14,   -41,    -8,     3,   -81,   -22,    42,    31,    27,    27,    -2,    13,     3,   -60,   -69,   -36,   -29,   -26,   -35,   -32,   -27,    12,    21,     4,    -4,   -72,   -12,    10,    59,    -3,    -2,     3,    -5,    32,   -11,   -37,   -51,   -53,   -96,   -28,   -22,     0,   -36,   -66,   -40,   -50,   -28,    -3,    -6,    -8,   -20,   -38,   -16,   -15,    24,    34,    90,    12,    -8,    -3,   -14,     4,   -51,   -72,   -25,   -34,   -59,   -69,   -54,    18,    23,   -45,   -66,   -25,    23,    15,   -13,   -25,   -65,   -44,     9,    15,     1,    35,    67,    23,     6,   -13,     7,    13,    17,   -15,   -36,   -81,   -39,   -46,    16,     8,    37,    19,    -2,    19,   -20,    21,    21,     2,   -13,     0,     6,    13,    18,    15,    25,    39,    -5,     4,     6,    22,    37,    15,   -23,     4,   -17,   -11,     9,    14,    23,     0,    43,    50,    44,    69,    -4,   -49,   -86,   -49,   -21,   -13,   -19,    13,    44,    36,     7,   -14,    27,    33,     3,    26,    -3,   -28,    -4,   -15,    25,   -18,    49,    -3,     4,     2,    14,   -10,   -25,   -41,   -21,    -8,     7,   -10,     5,    -5,    39,    58,     5,     2,   -33,    65,    38,    66,    45,    -4,   -26,   -11,    -7,   -30,   -14,    20,    17,    40,    21,    -4,   -11,   -15,     2,   -15,     1,    -5,    58,     9,    52,    93,     7,    -8,    -8,    57,    74,    34,    30,    10,    -6,   -17,    47,    24,    23,    -9,    -9,    16,    27,    22,    -6,   -41,   -22,    -4,    31,    19,    64,    36,    68,    72,    -6,     8,    12,    30,    38,    39,    45,    33,    12,     2,    -4,     0,   -30,     0,     0,    38,    24,   -17,   -12,    -3,   -23,    -1,   -18,    31,    60,    16,    67,   -10,    -3,    15,     8,    -6,    38,    56,   -11,   -19,   -13,   -12,   -19,   -33,   -33,   -75,   -36,    11,     6,    28,    64,    50,    26,   -45,    -3,    39,    45,    42,    58,     2,     0,    -8,    28,    16,    47,     1,   -38,   -45,   -32,   -27,   -39,   -51,   -62,   -81,   -34,     4,   -11,    30,    27,    11,   -27,   -11,    -9,    11,    38,   -27,   -35,     0,   -10,     1,    17,    19,    24,     7,    -6,   -17,    -9,   -38,   -51,   -47,   -71,   -56,   -43,     9,   -66,  -118,   -39,     4,    -6,     6,   -30,   -36,    -9,    18,   -11,    -6,     8,     9,   -25,    18,   -30,   -39,   -10,   -24,    -9,   -75,   -81,   -72,   -68,   -78,   -37,   -33,   -89,  -132,   -69,    20,     8,    19,   -29,   -14,    27,     1,    -4,    -8,    -2,     3,    -6,   -20,   -39,   -56,   -56,   -46,   -55,   -64,   -68,   -37,   -24,   -62,    12,   -20,   -51,   -47,   -99,   -88,   -44,     6,   -33,   -40,   -16,     7,     8,    -1,     3,    -8,    -3,     4,   -31,   -33,   -32,   -36,   -25,   -80,   -41,   -15,   -20,   -34,   -18,   -49,   -46,   -60,   -77,   -84,   -59,   -52,   -52,    -1,   -10,     7,    10,    -1,     6,     7,     3,     4,     1,    -8,     1,     0,    -7,    -6,   -35,   -25,    -5,   -28,   -22,   -24,   -22,   -14,   -16,   -21,   -60,   -65,   -23,     0,     3,    -3,     6,    -3),
		     3 => (   -2,    -9,     0,    10,     0,    -7,     6,     8,     9,     0,    -8,    -7,    -5,   -11,    -1,    -1,    10,     8,     8,     4,    -3,     0,     3,     7,     7,    10,    -5,    -6,     5,     4,     7,     2,     9,    -5,    -7,    -4,    -9,    -6,     2,    -6,   -16,    -4,    -9,   -19,   -25,   -22,     6,     4,     7,     6,     1,     0,     0,    -8,    -8,    -7,    -5,     8,   -10,     8,    -5,     9,   -13,   -11,   -10,   -37,   -40,   -12,   -34,   -43,   -27,   -32,   -55,   -68,   -58,   -31,   -84,   -72,   -81,   -25,    -6,     1,     2,     7,     9,    -7,     6,   -10,    -9,   -24,   -13,   -29,   -29,   -29,   -44,   -32,    -4,   -10,   -38,   -39,     6,    46,    28,   -21,   -11,   -19,   -58,   -75,   -36,    -7,    -4,    -5,     2,    10,   -10,    16,    45,    20,     2,    27,    35,    55,    45,    -5,     2,    21,    37,     8,   -34,   -11,    28,     2,    -9,   -68,   -30,  -128,   -83,    -6,   -23,     4,     5,     2,     4,   -15,    16,   -23,   -29,   -41,    12,   -34,    18,    17,     3,    -5,    -7,     2,     0,    18,    32,    13,    12,    33,    14,   -18,   -30,   -23,   -23,    -2,     7,     8,     5,    -7,   -26,   -11,    -6,    -1,    24,     2,     7,    -6,    17,    62,    25,    -2,    -7,     1,     3,    38,   -40,   -23,     7,    -1,    -2,   -34,   -42,    -6,     5,    16,     0,   -38,   -20,    51,     4,    -5,     9,    -1,    23,    41,     9,   -22,    11,    26,    39,    -4,    -7,     2,    41,   -11,   -30,   -64,   -38,   -56,   -38,    -9,     7,    -4,     8,    60,    27,    15,   -28,    31,    -8,   -50,    31,    19,    44,    13,     0,   -19,   -11,    14,    -5,     4,    22,    27,   -12,  -100,  -114,   -31,   -47,    -9,   -10,   -27,    74,    61,    13,   -66,   -20,    -8,   -27,    -8,   -42,   -33,   -77,   -95,  -147,   -65,    15,     5,    15,    23,    28,    13,     7,   -72,  -147,   -61,   -65,     3,     2,   -17,    98,    42,   -36,   -73,   -84,  -118,   -99,  -107,   -99,  -175,  -144,  -130,   -54,   -16,     4,   -18,   -12,     8,     8,    35,    21,   -27,  -132,   -36,   -36,   -11,     2,   -13,   -13,   -25,   -54,   -75,  -115,   -83,  -117,  -156,  -109,   -93,   -46,    36,    52,    53,     6,    19,     0,    26,    64,    43,    30,   -73,   -66,   -58,   -24,     0,    -8,    -3,   -37,   -54,    16,   -20,   -17,   -51,   -24,   -50,   -21,     7,    54,    50,    35,   -15,     4,   -18,    28,   -48,   -10,    -6,   -16,   -23,     3,    -9,   -12,    -9,     4,     0,   -50,     9,    61,    38,    -2,   -26,     6,   -22,    13,    44,    24,    35,   -17,    -4,    -3,   -37,   -43,   -63,   -41,    -6,   -20,    -2,   -39,   -40,   -18,   -11,   -13,    12,    -4,    -1,     9,    54,   -20,   -36,    54,    17,    -5,    18,    18,    19,    -4,     5,    -3,   -11,    -5,   -28,   -50,   -13,   -39,   -47,   -56,  -100,   -29,   -16,   -17,    29,    39,   -14,    33,   -11,   -69,   -89,   -54,   -35,     7,    15,     0,    43,    39,   -11,   -12,     6,   -10,     3,   -17,    -5,   -55,    -6,   -40,   -33,    78,     1,    -6,     4,    35,    42,    24,    -1,  -109,   -81,  -117,   -68,   -37,     7,    -9,    25,   -14,   -25,     5,     2,    -1,    21,    10,    27,   -42,   -24,   -63,   -34,    28,    -7,     0,    15,    49,    -6,   -50,   -15,   -75,   -26,   -84,  -154,  -187,   -76,   -84,   -83,   -46,   -32,    21,    19,    21,     1,   -13,    23,     6,   -33,   -63,   -64,   -28,   -11,   -19,    13,    66,    17,   -38,    29,    10,    47,    -6,   -21,   -64,   -44,   -94,   -89,   -36,    16,   -16,     0,   -13,    19,    34,    25,    -5,   -82,  -115,   -41,   -27,   -23,    -8,   -11,   -45,    76,    11,    12,    21,     8,    23,   -20,   -19,   -42,   -33,    20,    -2,    -2,    -9,   -12,    -2,    -2,   -10,   -22,   -38,   -52,   -85,   -35,   -31,   -17,    -9,     6,   -80,    59,    51,     3,    -3,     0,    30,     4,    22,    18,    18,    18,   -17,   -30,    -3,     2,   -16,   -15,    -3,   -36,   -60,   -77,   -70,   -20,   -17,    -4,   -20,     9,   -11,    28,    60,    -3,   -23,    15,    47,     2,    32,    14,     6,   -27,   -21,   -35,   -42,    12,    -7,   -50,   -23,   -22,   -41,   -83,   -65,   -24,     0,     5,    -5,   -17,    -6,    25,    18,    28,   -19,   -34,    -9,   -27,    -3,    -7,   -30,   -21,   -29,   -16,    -9,    25,   -46,    -8,   -49,   -56,   -81,   -78,   -64,   -28,    -7,    -6,   -10,     6,    44,    41,     7,    54,   -34,    10,   -25,    -7,   -18,    10,   -12,     0,    17,    -4,    59,    -4,     0,    54,   -27,   -64,  -109,   -82,   -36,   -56,    -5,     0,    -2,     0,    -7,    18,   -22,   -25,     7,   -19,   -21,    13,   -15,   -24,   -23,   -51,   -14,   -34,   -29,   -49,   -20,   -62,   -66,   -55,   -65,   -26,   -33,    -5,     4,     0,    -2,     3,     3,   -39,   -15,    -6,   -30,   -50,   -33,    -6,    15,   -48,    -3,    -9,   -26,   -73,   -74,   -67,   -25,   -17,     1,   -24,   -60,   -39,     4,   -14,     6,     2,    -6,    -8,    -2,   -30,   -10,     7,   -28,   -51,   -73,   -81,   -30,   -50,    19,    49,    31,     5,   -33,   -40,   -25,   -31,   -52,   -33,   -42,    -6,     7,    -5,     5,    -7,     6,     5,     6,     2,    -4,    -2,   -11,     1,     1,   -23,    -4,   -15,     2,   -12,   -29,    -3,   -31,   -27,     4,    -6,   -21,    -6,    -8,    -6,    -2,     6,    -6,    -1),
		     4 => (    4,    -4,     3,     2,    -5,     9,     7,    -7,    -4,    -3,    -8,     0,   -14,   -15,   -18,    -6,    -6,    -9,    -2,     7,     4,    -1,     5,    -1,   -10,    -6,    -6,    -3,     8,    -2,     3,    -9,    -2,     2,   -28,   -36,   -13,   -15,   -35,   -13,   -38,   -66,   -29,   -30,   -35,   -26,   -10,     4,   -24,   -13,   -22,   -28,     4,     3,     9,    -4,     5,     2,    -6,     7,   -35,   -10,   -37,   -43,   -64,   -28,   -31,   -69,   -42,   -44,   -26,   -25,   -60,   -49,   -47,   -11,   -60,   -54,   -48,   -41,   -12,   -35,     9,    -6,    -7,     2,    -4,   -28,   -72,   -35,   -53,   -31,   -33,   -43,   -23,   -45,   -49,   -42,   -41,   -45,   -72,   -86,   -42,    -9,     5,    -7,   -19,   -12,   -40,   -26,    -7,    -5,    -7,    -5,   -18,   -66,   -10,    11,    50,    14,   -21,   -62,   -41,   -21,   -18,   -57,   -97,   -76,   -44,   -70,   -39,    77,    36,    10,    47,   -27,   -33,   -17,   -30,    -8,    -7,    -4,   -33,   -25,    -6,    11,    43,   -16,   -10,   -21,   -19,   -19,   -14,   -84,   -98,    11,   -41,    14,   -33,    11,     6,     8,     9,   -57,   -24,   -17,   -17,    -8,     6,    -2,    -3,    -8,   -25,   -22,    47,   -40,    18,    31,     8,   -33,   -66,  -139,  -128,   -71,   -18,    11,    48,     0,    -1,     9,   -44,   -58,   -64,   -17,    -2,   -24,     6,   -39,    -9,     7,   -12,   -17,    22,    -3,    10,    12,    18,    18,   -61,  -110,  -153,   -62,   -25,    73,    49,    51,    19,    -8,   -39,   -56,   -55,    -3,   -15,   -57,   -36,   -86,     7,    -8,    20,    19,    29,    -9,    18,    48,    -8,   -17,     7,  -120,  -108,   -47,    67,    45,    27,   -17,   -39,    21,    -6,   -22,   -33,     6,   -52,   -77,    -6,   -57,    10,     9,    54,    24,   -65,   -12,    36,     5,    26,    31,    44,   -59,   -84,    -5,    97,    16,     9,     0,   -48,   -17,   -21,     5,   -58,    12,   -49,   -39,     9,   -30,    -1,    24,    18,    -7,  -115,   -29,    16,    40,    -9,    19,    40,   -62,   -68,    45,    45,     7,    34,    26,   -30,   -60,   -38,   -73,   -75,    16,    -3,   -25,     2,   -44,    15,     9,    28,     8,   -42,    -9,    16,    12,    26,    27,     7,   -92,   -94,     8,    24,    -2,    13,   -21,   -56,   -57,   -27,   -53,   -22,    15,   -19,   -58,     7,   -27,    20,    27,    28,    30,     8,     8,   -39,   -25,    23,     1,     9,   -26,   -62,    28,     3,     5,    -2,     9,   -38,     1,    40,    86,    84,    68,   -65,   -45,    -1,   -21,   -39,    -1,    46,    17,   -13,    -2,   -12,    22,    41,    -1,    -5,    -7,   -22,   -27,    16,    -5,    28,     3,    11,    43,    80,    40,    11,    -6,   -62,     2,    -7,    -6,   -40,     4,    22,    64,    10,    41,    19,    -7,    -5,   -12,   -20,   -11,   -44,     4,   -17,    11,    17,    39,     5,    57,    46,   -10,    25,   -23,   -36,    -4,     7,    10,    11,   -11,    51,    -5,    -5,    41,    -1,     5,     1,    13,     6,    36,    26,    36,    27,    13,    16,    39,    -2,   -11,    18,   -35,   -48,   -50,    20,    -8,    -9,    -7,   -57,    31,    52,   -27,   -32,    45,     3,   -16,     7,     3,    -7,    13,    38,    33,    -3,   -23,    26,     0,    -7,    17,   -38,   -52,    -7,   -16,   -23,     2,     0,    -7,    51,    37,    79,    -1,   -50,    10,   -31,     7,   -46,   -33,   -16,   -23,    10,   -33,   -44,   -43,    -7,   -73,   -26,    13,   -22,   -30,     2,   -12,     7,     6,   -37,    -6,    38,    45,    56,   -40,   -46,   -50,   -28,   -11,   -31,   -43,   -26,   -19,   -23,   -73,   -52,   -25,   -48,   -52,   -19,     7,     8,   -13,   -19,   -28,     8,    -2,    -4,     1,   -13,    19,    -6,   -62,   -11,   -68,   -37,   -13,    -8,    -5,   -39,    -3,    10,    -8,   -48,    18,   -37,   -12,   -19,    52,    17,     3,   -24,   -39,    -9,     0,     0,     0,   -12,   -41,   -93,   -60,   -55,   -13,   -44,   -53,   -33,    40,    15,    -6,    11,    -7,    -9,   -11,    29,     2,   -25,   -16,    -3,    -8,    -6,   -81,   -12,    -9,   -28,   -26,   -16,   -53,   -35,   -58,   -44,   -41,   -16,   -45,   -19,     6,     7,   -15,    24,   -43,    12,   -32,   -17,   -28,   -42,   -64,   -16,    17,     5,   -68,   -38,    -5,   -12,   -24,    -9,   -27,   -12,     0,     4,   -51,    11,   -70,   -50,     3,     7,   -24,    -9,   -25,    -4,   -22,   -14,   -44,   -37,   -56,     9,    29,    -4,     7,    17,    -6,    -8,   -10,   -14,   -28,     0,   -20,    31,    29,     7,   -85,    -9,   -28,   -29,   -26,   -20,   -30,     2,     3,    39,   -40,   -50,    -9,   -22,    15,   -24,    18,     4,    -6,    -7,     9,    -5,     6,   -70,   -19,   -29,   -19,    -5,   -16,   -40,   -18,   -35,   -26,    60,    -9,    38,    35,    49,   -45,    -6,     8,    -7,    -4,   -59,     3,   -17,    -5,     4,    -6,    -5,    -9,    -5,   -43,  -115,   -67,   -48,   -32,   -47,   -44,   -43,     8,    17,   -38,    -4,    18,     4,   -24,    -8,    27,   -31,    14,   -27,   -12,   -13,    10,    -7,    -4,     7,   -14,   -18,    -8,   -31,   -51,    12,   -11,   -60,  -102,   -88,   -68,   -31,   -51,   -89,   -22,   -55,   -70,   -90,   -85,   -70,   -16,   -26,    -2,     9,    -6,    10,     0,    -4,    -3,    -5,     5,   -31,   -26,   -35,   -39,   -31,   -66,   -36,   -28,   -76,   -22,   -33,   -44,   -34,   -48,   -58,   -51,   -40,   -13,    -6,    -1,     2,     8),
		     5 => (    6,    -3,    -4,     5,     9,     1,     3,     4,    -5,     8,     7,    -1,    -3,     3,     0,     9,    -6,    -7,     4,     9,    -9,    -3,     3,    -2,     5,    10,     5,     8,     9,     4,     9,    -7,     6,    -9,     2,     2,     7,     9,     6,    -7,   -20,   -19,   -20,   -18,   -13,   -21,    -7,    -5,   -12,    -3,    -3,     0,    -9,     7,    -8,    10,     9,    -6,    -2,   -10,   -10,    -7,     5,     6,   -11,    -4,   -35,   -71,   -64,   -88,   -31,    33,    30,    38,    56,    45,    57,    44,    42,    48,   -22,   -12,     3,   -10,     7,     7,    -5,    15,    38,    -9,   -23,   -18,   -15,   -50,   -57,   -44,   -18,   -44,    36,   -17,   -66,   -51,    -6,   -12,    18,    28,   -19,    -8,    26,    22,    30,    10,     4,   -15,   -19,     5,   -50,   -50,   -63,   -75,  -105,   -34,   -80,   -53,   -52,     1,    54,     3,    19,    -2,    -1,    -6,    10,    29,    39,    44,    55,   108,    29,    -9,    -1,    -8,   -11,    -8,   -46,   -44,   -91,   -90,  -108,   -57,    -8,    -4,    19,     1,     7,   -13,    16,    40,    23,     6,    77,    65,    36,    65,    70,   101,    48,   -15,     4,    -1,    19,   -15,   -47,   -83,   -83,   -51,   -26,   -48,   -13,     8,    49,     4,     0,     5,    21,    36,    76,    10,    63,     0,     6,    61,    22,    49,    33,     9,    -3,     9,    -7,   -27,   -40,   -55,   -24,    -5,   -16,     3,    -1,    46,    30,    11,   -18,   -26,     9,    27,    34,     3,    34,    -1,   -36,    -7,   -21,    21,    24,    17,    -9,   -12,   -30,   -25,   -32,   -21,   -51,   -24,   -39,   -54,    19,    55,    31,   -40,   -36,   -61,  -122,   -67,   -63,  -162,   -76,   -88,   -61,   -24,   -14,    -7,    18,     4,     0,   -16,   -61,   -69,   -62,    -9,   -59,   -67,   -57,   -30,   -28,   -16,   -21,   -35,   -67,  -153,  -191,  -220,  -238,  -230,  -161,  -123,  -112,   -62,   -38,   -31,     2,    11,     5,   -12,    -4,   -35,    -6,   -19,   -37,   -23,    -5,   -24,   -29,     6,   -30,     5,   -48,   -15,     4,   -47,  -138,  -142,  -139,  -114,  -108,   -74,   -41,     1,     6,     6,    -6,    -3,    -5,   -23,    -7,   -24,   -41,   -42,   -33,   -39,   -31,   -18,   -18,     0,   -22,   -20,    17,     5,    20,   -23,   -69,  -115,   -84,   -38,   -44,    -8,    14,   -19,     5,    -7,     0,   -22,    -5,   -19,   -18,   -34,   -20,   -34,   -16,    16,    15,    13,    14,     5,    10,   -22,   -21,     1,   -21,   -40,   -61,   -43,   -17,   -15,     0,   -28,    -3,     0,    -7,    -9,    -4,    17,   -26,     6,   -43,    16,    32,    58,    24,   -12,    23,     5,    -4,   -12,   -30,     9,     4,    22,   -25,   -16,   -34,     2,    -5,   -16,    17,    -9,    -5,     6,    34,   -33,   -57,   -48,   -10,   -16,    35,     5,     2,   -20,     8,   -38,    32,     6,     5,   -35,     1,     6,    -1,     1,   -14,   -10,   -17,   -16,    -2,   -28,   -18,   -14,    30,   -35,   -56,   -41,   -49,   -26,   -25,   -14,    21,   -24,   -46,   -12,   -36,    20,   -13,    -9,   -27,     9,    -5,    12,     9,    -8,    -9,    -5,    -1,     7,   -25,     9,    -1,   -50,   -53,   -79,   -81,  -131,  -104,   -64,    12,     8,   -35,    15,    12,    67,   -14,    21,    14,    17,    23,   -33,   -42,   -27,   -28,   -28,    -6,   -20,   -54,    13,   -25,   -31,   -38,   -80,   -38,  -101,  -138,   -46,   -57,   -74,   -58,    16,   -18,   -27,    58,    30,    35,    23,   -16,   -24,   -61,   -31,   -11,   -19,    -2,   -14,     3,    29,     2,   -26,   -42,   -11,    32,   -20,    -6,   -37,  -103,   -54,    -5,   -24,    13,     1,    39,   -19,    -4,    16,    -4,   -20,   -59,     8,   -50,   -39,     1,    -2,    42,    -4,     7,   -34,    -7,   -14,    22,    35,    10,    32,    23,    14,    20,   -10,    20,    -8,    16,    14,    14,   -19,     1,   -33,   -53,     4,   -15,   -20,    -7,    -5,    28,    14,    99,    -4,    11,    -3,    51,    36,     4,    14,   -38,    42,    38,    15,     5,    -2,   -19,    29,    21,   -26,    33,   -58,   -39,   -25,    -9,     3,     4,   -12,   -27,   -14,    63,    51,     1,   -11,    11,     3,    18,    33,    17,    22,    -9,    15,    19,   -23,   -35,    22,    35,    40,    35,     5,   -20,   -31,    -2,    -7,     7,     3,   -38,     9,   -29,   -17,   -29,   -16,   -22,   -16,    51,     9,    25,   -23,    -3,   -21,     4,   -11,    15,     6,    49,   -19,   -19,   -24,   -35,   -30,    -2,     3,     2,    -7,    19,    25,   -31,   -27,    11,     5,    54,    29,     8,   -45,   -18,   -18,    -2,    56,    -9,   -56,   -48,   -39,   -48,   -39,     5,    17,   -79,   -82,    11,    -2,   -10,    -2,   -35,    -3,    45,    37,   110,    53,    -9,    33,    66,     0,    18,    12,    40,   -34,   -53,   -26,   -42,   -49,    -9,    28,    36,    -7,     2,   -24,   -27,     7,    -8,    -2,    -4,    43,   -20,    -4,    38,    53,    14,    44,    36,    30,    15,     7,   -27,   -12,   -23,   -54,    12,    26,     7,    12,    27,     6,    -5,     4,    -4,    -6,    -5,     7,     9,     0,   -21,   -23,   -13,    -5,     3,   -10,    23,    20,    17,   -16,   -21,   -12,    -8,   -12,   -13,    -6,     9,     5,    17,    -9,     4,     3,     6,    -1,    -1,    -3,     6,    -8,    -3,     1,   -10,     5,    -2,    -9,    10,    -4,     2,     9,   -11,     3,   -10,    -9,   -15,   -18,   -15,   -15,   -14,     9,     4,     0,     7,    -7),
		     6 => (   -6,    -4,     5,     6,     6,    -9,    -6,    -7,     4,     6,     3,     6,    24,    13,    -2,     2,     3,    -2,    -7,     2,    -1,     5,    -6,    -4,     4,    -5,     7,    -3,     9,     8,    -8,    -9,     5,     3,    16,    20,    36,    50,    43,    19,    45,    31,   -15,     2,    20,    41,     3,    33,    38,    33,    29,    39,    10,     6,    -6,     6,     7,     5,    14,    30,    43,    25,    31,    34,     8,    -7,   -27,    36,    57,    26,    27,    71,    40,    18,    25,    -9,   -13,    -3,     7,    -3,    14,    16,    -3,    -9,     5,    -4,    -2,    88,    49,   -11,    42,    59,   -12,    10,   -27,    16,    16,    39,    19,   -17,   -15,     2,   -33,    -4,    29,    -1,    -6,   -14,   -13,     1,     7,   -10,    -1,     6,   -30,    42,    -4,    23,    24,   -19,     5,     1,    18,    27,   -31,    -6,    -8,   -42,   -25,   -27,   -33,    53,    44,    20,   -25,   -52,   -27,   -30,    -6,    19,    -7,     5,     7,   -15,    -1,   -59,   -46,   -19,   -32,    36,     1,   -27,    22,    31,   -15,   -20,   -48,    12,    16,    29,    12,    -1,   -28,   -45,   -31,   -14,    10,    21,    -7,   -10,    12,   -44,   -40,   -77,   -61,   -10,   -30,     1,   -48,    35,    50,     8,    -7,   -15,   -15,   -38,    16,    -4,   -43,    -4,   -52,   -68,   -14,   -19,    29,    -9,    -2,   -10,     4,   -42,   -37,   -95,   -61,   -30,   -13,   -14,    10,    56,    40,     4,    24,   -32,   -40,   -36,   -95,   -76,   -75,   -43,   -65,   -81,   -49,   -33,    19,   -49,     3,    -3,    10,   -44,   -33,  -104,   -14,   -18,   -46,    27,    13,   -10,    43,     7,   -35,   -70,   -66,  -112,  -101,   -98,   -66,   -75,  -125,   -95,   -81,   -57,   -17,   -44,     8,    -7,   -19,   -27,   -24,  -110,    -5,     8,    -9,   -33,   -27,     4,   -20,   -45,   -42,   -85,   -80,  -114,  -115,  -100,   -60,  -109,  -102,   -73,   -19,   -21,   -26,   -16,    -8,     3,   -14,   -30,   -52,   -99,   -59,     4,    25,     0,   -29,    -3,    23,   -34,  -100,   -93,   -22,    28,    -3,   -49,   -34,   -27,   -47,   -20,   -16,    30,   -36,   -43,     6,     0,     7,   -59,   -44,   -17,   -43,    -1,    33,   -24,    -6,    10,    21,   -80,   -73,   -19,    23,    31,    26,   -29,     0,   -67,   -33,   -47,   -45,    -8,   -59,   -31,     7,   -10,    10,   -33,   -41,   -46,   -24,    39,    25,    -8,   -29,     2,   -28,  -107,   -32,    -7,    41,    16,    -2,    30,    34,    -6,   -23,   -31,    46,   -15,   -35,   -33,     3,     1,   -25,   -19,   -70,   -59,     1,    50,    24,   -61,   -45,     2,   -21,   -46,   -36,     5,    -9,   -11,    -5,    40,    62,    28,   -11,    17,    11,   -16,   -35,    26,     2,     4,    -6,   -47,   -81,   -31,    42,    28,    13,   -16,    18,    47,   -11,   -13,    22,   -10,    19,   -31,    29,    25,    14,    32,    42,    14,   -11,     5,   -23,    -7,     4,    -2,   -11,   -41,   -60,     1,    60,    35,   -10,    -1,   -11,    63,     8,   -29,    42,   -16,     3,   -18,    24,     6,     6,    24,    50,    22,     0,    16,   -50,   -65,    -9,    -9,   -11,   -33,   -23,    35,    72,    -9,   -12,   -55,    31,    53,    -9,   -35,    52,   -10,   -12,     1,   -10,   -10,    19,    44,    29,     5,    12,    -1,   -62,   -55,    10,     0,     2,   -22,    -3,   -22,    32,    17,   -30,   -31,    -2,    22,    11,   -10,     7,    -6,   -13,   -32,    16,   -22,   -32,    38,    44,     5,    54,    48,   -25,   -51,     5,     0,     9,   -36,     0,   -18,    14,    32,     0,   -43,     5,    -6,    40,    14,    28,   -41,   -17,   -38,   -12,    20,   -12,    48,    17,    37,    33,    65,   -33,   -54,    -8,    -2,    -5,   -37,    28,   -55,   -42,    19,    -7,   -26,   -34,     7,    29,    26,    41,    34,     5,     3,   -28,    14,   -30,   -18,   -41,    35,    15,    43,   -15,    -4,     6,   -13,     1,   -37,    18,   -24,   -41,    -1,   -58,   -24,   -16,     0,   -21,     4,    55,    59,    13,     5,    43,   -12,   -14,   -17,    17,    32,    43,    54,    -3,     5,    -4,     2,     0,    -4,     3,   -16,     9,    -4,   -48,   -58,    -9,   -40,   -64,   -49,    38,    39,   -14,    16,    -5,     9,    28,   -29,    31,    54,    20,    11,    20,     3,     8,     6,    -8,   -17,   -17,   -22,    27,   -65,  -116,  -116,    -9,   -29,   -35,   -33,   -42,   -24,   -63,   -40,    22,   -42,   -42,   -41,    14,   -20,   -95,   -62,    19,    -7,    -7,    -6,    -9,    -1,   -33,     0,   -30,   -38,   -49,   -22,    57,    15,   -89,   -69,   -79,   -87,   -87,  -105,   -98,   -22,   -26,   -63,   -52,   -75,   -87,   -28,   -28,     1,     6,     3,    -6,    -6,    -9,   -11,   -15,    -4,   -16,   -17,   -32,    -1,   -22,   -49,   -78,   -56,   -35,   -52,   -59,   -96,   -42,   -44,   -20,   -29,   -47,   -32,     3,    -2,     0,    -4,     8,    -7,    -3,     6,   -12,   -16,     4,   -18,    -7,    17,    24,     7,    -2,    -4,     1,   -15,    -2,   -28,   -44,   -33,   -29,   -48,    -4,    -6,     1,     1,    -7,     5,    -5,     3,    -3,    -7,    -4,   -10,    -5,     0,     4,   -12,    -5,   -13,     1,     2,     4,     0,    -4,    -6,   -13,   -11,    -8,     3,     7,     5,    -5,     1,     2,    -3,     1,     9,    -6,    -2,   -10,    -6,     4,     1,     3,    -5,    -3,     8,    -1,     5,     7,    -4,    -3,     7,    -5,     1,   -11,     5,     1,    -5,     5,    -2),
		     7 => (    3,     2,    -7,    -2,    10,    -9,    -9,    10,     1,     7,     3,     3,    -4,    -5,     2,    -3,    -6,     4,    -3,     5,     3,    -2,     7,     9,     0,    -9,    -4,     6,    -2,     3,    -4,     0,     2,    -9,     3,     2,    -5,     8,   -13,   -23,    -8,   -21,   -25,   -25,   -42,   -44,   -27,    -9,    -4,    11,    14,    -6,     9,     1,    -8,     3,    -1,    -8,     5,    -5,    -6,    -9,     2,   -16,   -23,    -7,   -47,   -84,   -40,   -23,   -18,   -12,   -22,   -11,     0,    -4,   -20,    -4,    -9,    16,     4,   -11,     5,    -3,     7,     2,     1,   -10,    -2,   -32,   -49,   -39,   -47,    -7,    -9,   -31,   -57,   -72,   -37,   -32,   -32,   -16,     0,   -23,   -14,   -11,   -27,   -17,    -4,     2,    10,    -8,     7,    -3,    -9,    -3,   -18,   -20,   -20,   -61,   -80,   -40,   -82,   -23,     9,    -6,   -43,   -64,   -75,   -83,   -57,   -44,   -33,   -25,   -53,   -75,   -52,   -46,   -31,     0,     2,    -4,    -1,   -62,   -18,    43,    66,    37,    60,    19,   -31,    12,    11,    17,    35,    20,     9,   -12,   -46,   -61,   -99,   -66,   -59,   -90,  -135,   -92,   -26,     9,    -8,     5,   -13,   -44,    -6,    31,    32,    31,    14,    -4,    32,     0,    48,    21,    22,   -25,   -37,   -24,   -46,     0,     1,   -20,   -52,   -51,  -103,   -54,   -57,   -19,    -4,    25,     0,    14,    13,    30,    15,    -3,    -3,   -33,     8,   -29,    23,   -13,   -33,   -57,   -28,   -34,   -51,   -47,   -10,   -42,    11,    16,   -17,   -59,   -65,   -24,   -29,    57,    29,     4,    51,    66,     0,    32,     9,    20,    10,   -37,   -24,   -18,   -24,    20,    15,    11,    -5,    -8,     4,     2,    -7,   -26,     1,   -87,   -80,   -29,     0,    42,    10,    29,    46,    61,    19,    13,    70,    21,   -34,   -43,   -33,    -3,    -8,    12,   -23,     0,    23,    -9,    22,    22,    25,   -20,   -29,    -2,    61,    82,     7,    -6,     6,   -19,    23,    -8,    33,    42,    37,    -2,    -4,     9,   -25,    -5,   -19,   -11,   -11,    25,    40,    17,    29,    21,    14,   -10,     0,    40,    26,    71,     0,   -25,    14,    41,    -4,   -18,    51,    76,    49,    39,     4,    -1,     2,     9,     9,    -8,   -24,    47,   -25,    47,    24,   -17,   -29,   -37,   -19,   -58,   -16,    54,     1,     9,     9,   -28,   -46,   -79,    -4,    -3,     8,     2,   -32,   -26,   -25,   -58,   -35,    -8,   -22,   -41,     4,     1,    -3,    -8,   -26,   -17,   -11,    10,    41,    66,    -9,    16,    41,   -51,   -54,   -61,   -22,   -21,   -46,   -59,   -67,   -63,   -97,  -104,   -14,    -9,    -2,   -14,    40,    16,    25,   -16,    13,    58,    24,    25,   -46,   -41,   -16,   -15,   -14,   -45,   -40,   -67,   -47,   -67,  -107,   -84,   -75,   -76,   -89,   -50,     9,     5,    21,    -6,    24,    40,    52,   -26,     9,   -10,   -30,   -73,   -52,   -11,    -2,     1,   -23,    -6,   -73,   -33,   -30,   -91,   -48,   -35,    -4,   -10,    15,    -2,    28,    33,   -18,    19,    13,   -14,    54,     8,    28,   -12,   -19,   -91,   -36,   -16,    -8,   -16,   -18,   -15,   -49,   -44,   -45,   -61,     4,    37,    36,    34,    38,    23,    25,   -34,   -27,    -3,   -10,    13,    -2,    16,    28,   -31,  -102,  -100,   -43,   -27,    -6,    -9,    -3,   -33,   -31,   -39,   -57,   -70,    -1,    10,   -42,    -2,     3,    18,    20,   -33,   -23,   -46,    15,    24,     9,   -14,    17,   -25,   -40,     7,   -10,   -20,    12,   -11,    48,   -24,   -48,   -78,   -86,   -55,   -34,   -91,   -61,   -10,    48,    51,   -48,   -47,   -37,   -14,    -9,   -41,   -31,   -46,   -23,   -42,   -37,   -21,    32,   -16,    -6,    18,     7,   -15,   -39,   -97,   -51,   -56,   -45,    15,   -29,   -27,    -2,   -13,   -31,   -26,   -10,   -47,   -29,   -20,   -24,   -42,   -35,   -45,   -78,   -10,   -40,     0,     7,   -12,     2,   -19,   -54,   -10,     6,    25,   -21,   -12,   -10,    -7,    12,    13,   -44,   -54,   -43,   -69,   -68,   -51,   -19,     3,    18,    -3,   -34,   -16,   -65,    -6,   -12,   -10,    -4,   -56,   -40,    42,    49,   -27,    16,     0,   -14,   -30,   -15,    16,   -97,   -64,   -88,   -94,   -55,   -61,   -50,    -8,   -13,   -45,   -37,   -10,   -16,   -14,   -22,   -17,   -15,   -86,    29,    45,    42,    52,    64,    19,    19,     2,   -22,   -38,   -63,   -60,   -65,   -52,   -72,   -52,   -55,     7,    15,   -95,   -54,    -7,   -20,     2,     0,     8,   -24,   -99,    25,    -5,    33,    84,     5,     1,   -13,    22,   -32,   -22,   -61,   -28,   -69,  -114,   -89,   -82,   -78,    -7,     1,   -43,   -32,    -4,   -47,     1,   -10,     0,    20,    -6,    41,    61,    42,    15,    51,     9,   -19,    15,   -15,    20,   -36,   -29,   -97,  -100,   -82,   -51,   -70,     5,   -19,   -75,   -11,   -28,    -7,     8,    -8,    -3,   -17,    38,   -40,     8,    -2,    18,   -22,   -45,    -8,    26,   -11,   -54,   -70,   -54,   -65,   -37,   -24,   -35,   -89,    -8,   -13,   -58,    10,     1,   -11,    -9,     9,     5,    -4,   -45,   -52,   -57,   -14,    28,    48,    18,   -27,    -2,    15,    31,   -35,   -12,    -3,   -20,    10,    -4,   -27,    27,    39,    18,   -14,     1,     7,    -8,    -1,    -3,     1,     7,    42,    39,    -9,    -4,   -11,     1,    26,    19,   -18,    58,    39,     3,    15,     8,     9,    -8,    12,    46,    35,    41,    -3,     6,     1,     2),
		     8 => (   -4,     3,     1,     4,    -4,     6,    -7,     1,     8,    -5,    -3,     8,    -2,    -1,    -1,    -7,    -8,    -6,    -4,    -4,    -9,    -6,    -5,    -7,     0,    -1,    -3,     6,     5,    -5,    -6,     7,     3,     8,     8,    -8,     7,    10,     1,     3,    -1,   -12,    -8,   -11,   -28,   -23,   -13,     6,    -6,     1,     6,     5,     0,     8,     7,    -4,     4,    -7,    -8,     8,    -9,     8,    -4,    -3,   -10,   -28,   -72,   -63,   -17,   -16,   -10,   -30,   -40,    31,    47,    16,   -30,   -30,   -28,   -30,   -10,   -15,     8,    -2,    -3,    -9,   -22,   -20,   -17,   -29,   -18,   -56,    39,    30,   -17,   -46,   -42,   -31,   -30,    12,     9,     8,    64,    32,     1,   -22,    41,    56,    -1,   -14,   -20,     9,     1,    -6,   -20,   -30,   -55,   -73,    -1,    30,    -7,   -44,   -38,    23,   -13,    -2,    12,    15,    19,     6,   -10,     2,   -23,     0,    23,   -25,   -44,    33,    38,    -1,    -5,    -5,   -15,   -32,   -33,   -54,     2,    -4,   -54,   -29,   -18,     0,    -6,    21,    -5,    16,   -19,   -55,   -67,    39,    -7,    39,     4,   -18,   -19,    -5,   -19,   -15,     5,     0,   -32,   -57,   -41,     7,    -8,   -25,   -44,   -20,    10,   -21,   -17,   -19,   -47,     0,   -29,   -29,   -29,    18,     2,   -16,   -15,   -42,   -37,   -27,    -6,    -5,     6,   -44,   -13,   -21,    -4,    -5,   -21,   -22,    -5,    -8,   -34,    -8,   -24,   -54,   -32,    14,   -11,   -39,   -27,     7,     3,   -10,   -40,   -33,   -34,    -3,    12,    28,   -19,   -33,    -9,    -6,   -22,    -3,   -38,   -17,     6,    19,   -48,   -37,   -24,    -7,   -20,   -19,   -32,   -43,   -25,     6,     9,    16,   -53,   -60,   -19,     4,    61,    30,    -4,   -13,   -32,     4,   -15,   -17,   -32,    14,    -2,   -21,   -49,    -6,   -17,   -31,   -46,   -43,   -22,   -23,   -49,    23,    10,   -53,   -57,   -49,   -41,    -2,    21,   -31,     8,   -14,   -28,     0,   -13,    10,   -27,   -27,    -8,     2,    22,    62,   -19,   -25,    15,     6,     6,     5,    15,    27,     3,   -19,   -40,   -62,   -28,   -36,     8,    13,    -1,   -12,   -13,   -31,   -21,    25,    15,     0,    15,    38,    21,     6,   -25,   -43,   -17,   -12,    19,   -10,     4,   -37,   -40,    41,   -26,   -26,   -13,   -79,    -5,   -40,    -5,     3,   -29,    -2,    29,    39,    26,    -8,    11,    35,    26,   -37,   -23,   -41,   -33,   -44,   -25,   -17,    -1,   -43,    -5,    21,    23,    35,    11,   -69,   -72,   -54,    10,    -4,   -37,   -58,     8,    22,   -14,   -53,    26,    79,    30,    24,    -9,   -27,   -37,    -4,     4,   -63,   -19,     2,    20,    48,    36,    36,    -6,   -61,   -94,    12,     0,     3,    -2,   -71,   -33,   -11,   -21,   -58,    12,     9,    -7,     1,    10,    -3,   -24,   -23,   -85,   -37,    28,    41,    41,    33,   -17,   -54,   -77,   -57,   -91,     1,   -10,     3,   -16,    19,     9,   -37,   -30,   -27,     4,    -6,    22,    34,    -3,    -4,   -32,   -70,   -26,   -14,   -28,    10,   -12,   -48,   -57,   -29,   -22,     0,   -46,   -36,     4,    -5,    -8,    36,    -6,   -31,   -35,   -32,   -80,   -53,   -16,    20,    25,   -28,   -21,   -18,    -3,    -9,    -5,   -30,    -7,    11,   -27,    -9,     6,    -9,   -52,   -28,     4,    -6,   -19,    26,   -24,   -35,   -44,   -25,   -69,  -125,   -49,    13,    37,    -6,    -6,     7,     7,   -21,   -52,   -47,     8,   -22,   -24,   -23,   -19,   -10,     6,   -15,   -11,     4,   -22,   -26,   -15,   -28,   -37,   -38,   -24,   -42,    -2,    -3,    21,    14,   -22,    26,    19,   -15,   -14,   -16,     4,   -30,   -15,   -31,   -13,    -5,    -9,   -23,     5,    -5,   -18,   -14,    -8,   -25,   -50,   -61,    17,    19,    -2,   -14,    25,    16,   -12,    35,   -29,    -7,     0,     2,   -35,   -29,   -24,   -21,     1,    -2,   -31,   -35,     8,    -5,   -15,     0,   -22,   -18,   -58,   -64,   -14,    16,   -12,   -13,   -11,    20,   -28,     6,   -45,   -46,   -16,    -3,   -60,   -24,    -6,     3,     1,    -1,   -23,    -1,   -17,    -8,   -19,    -1,   -26,   -32,   -46,   -10,   -37,   -33,   -20,    15,    53,    16,    19,     8,   -24,   -23,   -16,   -19,   -33,   -27,   -16,   -15,   -24,   -12,   -29,   -10,   -16,   -23,   -10,   -15,   -21,   -63,   -72,   -40,   -26,   -25,   -57,   -27,    30,    23,    24,   -38,    -4,     3,    -2,     2,   -15,     1,    -2,    -3,   -15,   -11,   -28,    -2,    -7,     1,   -24,    -7,    -8,   -33,   -61,   -80,   -27,    -5,   -29,    -2,   -29,   -12,   -41,   -17,     8,   -28,   -24,     2,    19,    20,     6,   -12,     1,    -2,   -32,    -1,     9,    -5,    -5,    -7,   -14,   -23,   -22,   -38,   -29,   -28,   -70,   -23,   -30,   -32,   -16,    26,    21,   -21,    34,    19,     3,    -5,   -14,   -16,   -54,   -38,   -14,     8,    -3,     7,   -14,    -5,   -13,   -35,   -24,   -13,   -24,   -26,   -40,   -50,    -8,    14,   -12,    23,    -5,    -6,    21,    20,     8,   -40,   -14,   -16,    -1,   -16,    -6,     5,     3,    -5,    -4,   -14,   -11,   -24,   -38,   -13,   -11,   -19,   -29,   -61,   -73,   -59,   -61,   -90,     1,    -8,   -10,   -75,   -68,   -38,   -27,    10,    -9,    -5,     9,    -6,     2,    -4,    -6,     3,   -14,    -4,   -12,    -6,    -2,   -19,    -5,   -22,     6,   -19,    -1,    -2,     0,     5,    -2,    -4,    -2,     4,   -10,    -5,     5,     8,    -3,     5),
		     9 => (   -3,    -5,     6,    -6,    -5,    -9,    -6,     8,     5,     1,    -8,    -1,     2,     0,     9,    10,    -4,    -1,   -10,     5,    -1,    -6,     5,     4,    10,   -10,    -2,     1,    10,    -5,     8,     7,    -8,     5,   -11,    -5,     9,    -2,    -5,    -5,   -27,   -15,    -4,    -2,   -10,   -10,   -18,     7,     1,   -13,    -6,   -10,    -2,    -3,    -4,    -4,    -1,     1,     7,    -5,     4,     8,    -1,    -1,    -7,   -11,   -14,    -2,    -3,    -4,   -27,    -5,   -12,    -4,    -9,    -2,   -25,    11,   -10,   -12,   -10,     9,     0,    -5,    -1,     0,     6,   -17,    -2,   -16,   -12,    -2,   -32,   -14,   -20,   -44,   -28,   -10,   -24,   -25,   -27,   -12,    25,   -14,   -25,   -33,   -26,     2,   -14,   -11,     1,    -5,     0,    -8,     0,   -16,   -15,     5,   -43,   -11,   -12,    -5,   -18,   -22,   -59,   -78,   -88,   -85,   -46,    -5,    31,   -42,   -64,   -45,   -33,   -29,   -26,   -57,   -40,     4,    -1,     5,    -9,   -13,     3,    -9,   -18,   -22,   -57,   -33,   -50,   -15,   -16,    19,   -22,   -34,   -70,   -75,   -72,   -62,     8,   -32,   -41,   -47,   -30,   -26,   -63,     4,    -9,   -13,     1,   -14,    17,   -26,    -9,   -61,   -48,   -47,   -63,   -23,   -29,   -47,   -16,   -18,   -18,   -46,     3,   -31,    15,    28,     1,   -19,   -28,   -34,   -43,   -39,    -4,   -15,   -23,   -21,   -32,   -54,   -57,   -69,   -80,  -111,   -90,   -71,   -34,   -28,   -36,   -67,    21,    14,    -6,    -9,    84,    32,    31,    23,   -14,   -40,   -16,   -26,   -33,   -11,     8,     0,   -39,   -30,   -37,   -51,   -60,   -86,   -28,   -56,   -25,   -12,   -54,   -21,     7,    31,    33,     3,     5,    -5,    -4,    35,    13,   -25,   -37,   -19,    -8,   -18,    49,    -5,   -21,   -35,   -20,    -9,   -66,   -13,   -14,   -23,   -28,   -53,    10,    41,     7,     3,    -9,    27,   -34,     6,    16,    -1,    29,    27,   -80,   -38,     0,   -12,   -33,   -28,    -4,   -24,   -45,   -56,   -21,    -2,    -9,    17,   -24,    17,   -10,   -38,   -38,   -31,   -73,   -66,   -32,   -14,   -26,    -7,    45,    96,   -34,   -58,     9,   -81,   -18,   -13,   -22,   -37,   -33,   -11,    47,    24,    32,   -12,     9,   -15,   -42,   -71,   -80,   -92,   -41,   -16,    24,    -9,    23,    10,    67,    90,    -7,   -51,     4,    -8,     7,   -48,    21,   -23,   -42,    -4,    21,    11,    37,   -18,   -54,   -38,   -68,   -47,   -21,   -71,     0,    -1,    44,   -13,    29,    36,   -14,   -69,   -59,   -58,    -8,   -15,   -21,   -35,    23,   -30,    -3,    14,     7,    23,    52,     5,     5,     9,   -30,    27,    50,     3,    -2,    54,    19,    57,     9,   -20,   -46,   -30,   -33,     4,     1,   -15,     4,   -32,    26,   -28,    -3,   -23,    51,    53,    46,     0,    21,    25,    21,    32,     5,     7,    -3,    25,   -16,   -57,   -23,   -71,   -65,   -13,     8,     2,    -6,     7,   -58,   -38,    27,   -29,   -41,   -33,    10,   -26,     7,    24,    25,    55,     2,    15,    -7,     2,    32,    13,   -46,   -56,   -77,   -60,   -48,   -10,    51,   -10,   -11,   -15,   -38,   -33,    18,   -19,    -6,    -2,   -27,   -13,    13,    19,   -18,    10,   -39,   -44,     1,    22,    11,    -6,   -68,   -24,   -22,   -72,   -35,    -3,    -9,    -4,     5,   -11,   -32,    -9,   -27,   -31,   -21,    29,   -28,   -49,   -35,   -25,   -18,    -9,   -25,   -11,    -2,    35,    27,   -27,   -35,   -16,   -36,   -71,   -30,    39,    -4,   -15,    -1,     7,   -33,   -14,   -66,   -48,     0,    25,   -32,   -53,   -11,    14,   -20,   -12,    22,   -25,    -6,   -15,    16,     4,   -31,   -24,    -5,   -27,   -17,    47,   -27,   -27,    -2,    -9,   -37,   -24,   -71,   -59,   -26,   -23,   -43,   -65,   -41,   -53,    -6,   -28,    -5,   -34,   -38,   -25,   -11,     2,   -67,   -31,    -5,   -13,    15,    55,   -36,   -25,     6,    -1,    25,   -20,   -51,   -30,   -89,   -69,    21,   -27,   -59,   -10,    34,    24,   -12,   -39,   -13,    -4,     2,   -14,   -38,   -33,   -25,    -6,    13,    47,   -10,    -7,    -2,    -8,    -9,   -26,   -54,   -26,   -62,   -46,    16,    22,     4,   -23,   -11,   -29,   -24,   -75,     3,   -18,   -17,    14,   -35,   -27,   -37,   -16,    11,    39,   -39,    -4,     7,     6,   -32,   -52,   -63,   -51,   -81,   -27,    16,    27,    30,    21,   -11,   -34,   -54,   -39,   -24,   -15,   -58,     2,     9,   -34,   -17,     3,    15,    -4,   -22,    -8,     1,     6,   -29,   -37,   -79,   -39,   -51,     8,    44,    32,    10,   -33,   -10,   -50,   -51,   -13,     3,    -7,   -11,   -10,    11,    -3,     6,   -32,   -11,    16,   -20,     7,     7,     8,   -16,   -27,   -37,     0,     4,    25,    10,    32,    11,   -12,     1,   -51,    10,   -36,   -32,    -1,   -27,    19,     4,    -2,    17,     1,    -6,    -5,   -13,    -1,   -10,     8,    32,   -14,    14,    -6,   -17,    -3,    20,    11,    32,    -4,    27,    -1,   -30,   -28,     9,    41,    25,     7,   -14,   -20,   -25,    22,     5,    -5,    -5,     3,     8,    10,     1,    54,    25,   -10,    31,    27,   -21,     3,    16,    48,     8,    39,    31,    18,    55,    69,    37,    26,    52,     8,   -21,    15,   -11,     2,     3,    -9,    -6,     5,     9,    -5,   -15,   -10,    14,    55,    47,    33,    32,    67,    35,    30,    25,    25,    13,    24,    39,    51,   -19,   -24,   -13,   -13,    10,    -3,    -9,    -3),
		    10 => (    5,     8,     3,    -9,     4,    -4,    -8,     2,     7,    -5,     4,    -2,    -8,     1,     1,     2,     3,    -4,    -7,    -5,     2,    -4,     0,     5,    -9,    -1,     0,     5,    -1,    -9,    -7,    -9,     6,     9,    -4,     5,     9,   -11,   -11,    10,    23,     3,   -17,    32,    41,    45,     1,     7,     7,    -1,     1,    -5,    -2,     1,    -5,     6,     9,    10,   -12,    37,    34,   -10,    -9,     7,   -13,   -17,   -30,    -4,    -1,   -22,   -11,   -47,    -6,   -55,   -46,   -50,   -40,   -14,   -46,   -28,   -22,    -7,   -10,     9,     9,     5,     5,    -2,   -11,    -1,   -13,    -3,    18,   -30,   -78,   -47,     4,    11,    -7,   -39,   -32,   -63,    -7,    -2,     4,   -37,   -38,   -21,    -4,     7,   -70,     0,     7,     7,   -10,   -15,    11,   -51,   -34,   -42,   -28,   -52,   -55,   -45,   -80,   -84,   -17,    15,   -40,    11,   -18,     1,    -7,     3,    15,    12,   -36,   -54,   -58,    -7,    -7,   -10,   -23,    -8,     8,   -60,   -29,   -59,   -18,    -1,   -70,   -29,   -51,   -33,    -5,   -10,   -25,    -2,   -25,    -6,   -70,   -33,    35,     3,   -56,   -37,   -48,   -36,     3,     5,   -40,    -5,   -11,    -5,   -25,   -25,     8,    -7,   -22,     3,   -20,     3,     2,   -23,   -15,     0,     9,     5,   -32,    24,    44,   -26,   -56,   -56,    -3,    -8,    -1,   -48,   -26,   -16,   -10,     5,    -7,   -41,    -7,   -20,    -6,     7,    -8,   -21,   -17,     8,   -27,     6,    28,    10,   -55,    -3,   -19,   -25,   -80,   -57,   -40,    22,    86,   -68,    34,    16,   -11,   -15,   -13,   -46,   -25,   -23,     1,    -3,    13,   -78,    12,    33,    -1,    45,    31,   -40,   -56,   -13,   -25,   -26,   -81,   -32,   -60,    -9,     6,   -14,    52,    -6,   -11,    11,   -31,    10,    18,   -19,     9,    -6,     2,     0,   -21,   -25,    34,    17,    29,   -13,    30,   -15,   -36,   -35,   -33,   -74,   -64,    -1,    -3,     4,    31,    17,    -7,    -4,   -10,   -16,   -14,    -7,    11,    -5,    -1,   -15,     8,   -67,   -23,    23,    -4,    -2,   -16,   -34,     4,   -10,   -48,   -44,   -52,    -4,    -7,   102,   -34,   -35,   -39,     9,    15,   -32,   -65,   -55,    -7,     5,   -14,    15,   -42,   -73,   -58,   -11,    18,    27,    -4,   -60,   -62,   -46,   -62,   -59,   -35,     5,     2,    14,   -16,   -44,    38,    42,    11,   -25,   -91,    -9,    15,     7,    34,    -4,   -58,   -77,   -33,     6,    34,    44,    13,   -48,   -58,   -23,   -48,   -62,   -23,    -8,    -7,    23,    28,   -36,    73,    36,    22,     5,   -34,    29,    15,    -9,     5,   -40,   -96,  -131,   -50,     3,    11,    47,    66,   -41,   -22,    26,     6,    -4,   -39,   -15,     7,     5,   -10,   -49,     3,    43,   -34,     9,    24,    25,    11,    54,    43,   -11,   -69,   -54,   -43,   -32,    25,    65,    57,   -44,    -1,    38,    -4,   -23,   -21,   -13,     8,    -7,   -34,   -60,   -39,   -23,   -23,    -9,    20,     7,    25,    47,    97,   -37,   -98,   -50,   -18,    -3,    53,   -12,    23,   -53,    -4,    23,   -13,   -15,   -79,   -14,     8,     5,   -28,   -36,   -27,   -10,   -40,   -42,    30,    -9,   -15,    23,    29,   -71,  -103,   -10,    16,    20,    22,    19,   -41,   -70,   -47,   -15,   -33,   -45,   -68,    64,     6,   -15,   -33,   -44,   -10,   -29,   -55,   -18,    11,   -14,     2,    -1,    15,   -58,   -56,    -6,    20,    16,   -17,    16,    -6,   -67,   -27,   -31,   -32,   -40,   -40,   100,    -3,   -14,   -37,   -37,   -35,   -70,   -44,   -24,     3,   -12,    16,     8,   -40,   -50,   -34,     4,    51,    15,     9,   -22,   -33,   -42,     0,   -34,   -17,   -29,   -49,   -24,     2,    29,     0,   -27,   -39,   -41,   -61,   -24,    37,     7,    -3,     8,    -8,     9,   -21,   -18,   -47,   -26,    33,   -17,   -17,     3,   -30,   -35,    -5,   -53,   -30,   -11,   -10,    36,   -14,   -33,   -10,   -40,   -70,   -31,    14,     7,    26,    29,    36,    22,    -6,   -63,   -47,   -10,   -32,     4,   -18,    14,   -36,   -11,   -42,     4,    24,     7,     7,     3,   -19,   -43,   -49,   -24,   -44,   -30,     2,    10,    53,     5,    47,    20,   -31,   -30,   -26,   -27,     6,    24,     2,   -21,   -38,    -7,     0,    11,   124,    29,     7,    -9,   -40,   -66,   -55,   -29,   -50,   -37,   -21,    33,    -3,    -2,     3,   -53,    12,    24,    25,   -31,   -57,   -11,   -51,   -42,   -29,   -18,    -6,    20,    69,    28,    -9,     6,    -4,   -44,   -52,   -83,   -35,   -28,   -32,    36,    69,    23,    13,   -13,    -6,   -34,     6,   -21,     0,   -11,   -51,   -41,   -12,   -14,     0,     2,   -56,     1,    -5,    -2,   -15,     0,    27,    19,   -54,   -69,   -75,   -57,   -50,   -30,    -8,   -36,   -48,   -29,   -35,   -15,    25,   -64,   -39,   -35,   -24,    -8,     8,    11,     6,     5,    10,    -2,   -12,     0,   -39,   -33,   -37,   -57,   -16,   -28,   -73,   -85,  -141,  -136,  -140,  -109,   -63,   -52,   -53,   -51,   -64,   -51,   -28,   -23,     3,    -3,    -4,     4,     9,    -9,     4,     7,   -25,   -37,   -90,   -27,   -36,   -69,   -45,   -51,   -36,   -37,   -14,   -49,   -47,   -50,   -67,   -58,   -51,   -42,   -20,   -22,     1,     5,     5,     4,    -3,    -7,    -9,     9,    -4,     6,    -9,   -16,   -20,     1,    -4,    -4,    -1,   -11,   -12,   -13,    -7,     0,    -9,    -2,     4,   -11,    -2,   -10,     4,    -7,    -7,     2),
		    11 => (    1,     2,    -8,   -10,     8,    -9,     9,     6,    -1,     5,     9,   -10,    -6,    -7,     8,    -9,     2,     7,    -5,    -2,     1,    -7,     3,    -7,     7,    -2,     8,    -7,     1,    -3,    -8,    10,     0,    -9,     1,     5,     9,     0,     1,   -10,    -5,   -18,     1,   -14,   -19,   -16,    -2,    -8,     2,    -7,    -6,     7,    -7,     9,    -4,    -7,    -9,   -10,    -7,    -9,    -9,     1,     7,     3,   -17,    -8,    13,     9,     2,    -7,   -11,   -32,   -74,   -89,   -72,    18,    23,   -30,   -14,   -24,    -9,    -8,     2,     3,     5,   -10,    26,     4,    -5,    -9,   -10,    33,    30,    41,    32,     8,     7,    -1,     9,   -46,   -75,   -56,    -7,   -25,   -24,   -41,    11,    31,   -29,     0,    -1,     9,    -5,     7,    23,    20,     9,    20,    29,    26,   -10,     2,   -28,   -23,   -21,   -27,   -30,   -59,   -45,   -22,     8,    18,    40,    -1,    -1,   -16,   -46,   -35,   -51,   -43,    -3,    -5,     2,    44,    34,    34,    -7,     2,   -52,   -29,   -43,   -47,   -21,   -15,   -89,   -96,   -62,     7,    19,    10,    -2,    39,    32,    14,     8,   -31,   -37,    -3,    -2,    -1,    -6,    39,    69,   -11,   -26,    -5,   -58,    36,    29,    -3,   -88,  -101,  -128,  -105,   -50,   -32,    -1,   -11,   -12,     7,     0,     7,   -27,   -42,   -29,   -19,     5,   -15,   -24,     2,   -29,   -34,   -26,   -33,   -67,     0,    42,     3,   -56,   -80,   -89,   -70,   -23,   -13,    26,     0,     5,    -6,    -6,    11,   -56,   -83,   -50,   -14,    -1,   -36,   -28,    -8,   -14,   -20,   -20,   -41,   -40,   -15,     5,   -55,   -43,   -49,   -87,   -43,    -1,    18,    11,    -3,    18,   -13,    -2,    -5,   -56,   -68,   -51,   -15,    -5,     3,   -26,   -10,   -15,   -22,   -18,   -19,   -19,    -4,   -73,   -82,   -87,  -140,  -123,     0,    32,     6,    14,    -7,   -10,   -13,     3,    -3,   -14,   -41,   -15,   -30,    -7,     4,   -13,    -5,     0,     0,   -45,   -47,   -66,   -40,   -73,   -71,   -96,  -118,   -58,    -4,    54,     9,   -18,    -7,    -2,    16,    12,    -4,     9,   -20,   -24,   -19,    -9,     4,    12,     6,   -14,     8,   -20,   -54,   -60,   -48,   -62,   -38,   -57,   -43,   -28,    63,    24,    22,    65,   -13,    -2,     6,   -37,   -54,   -34,     5,   -30,     5,    -4,     2,   -28,    15,    -2,    19,     6,   -43,     5,   -71,   -45,   -50,   -17,   -30,    18,    48,     3,    25,     9,    16,   -48,    -3,   -40,    -8,   -28,     4,   -14,     1,    -8,     3,   -22,    -1,     2,   -23,   -12,   -24,   -19,   -40,   -18,   -10,   -33,     8,    47,    31,     8,    30,    21,   -21,  -109,   -47,   -47,   -17,   -21,   -11,    -1,     2,    -5,    -3,    -4,     0,    13,   -15,   -12,     1,    -7,    29,    35,   -14,    -3,    33,    13,    16,    27,   -44,   -60,  -128,  -139,   -17,    19,    -2,   -11,   -24,   -15,    -6,     2,   -10,    25,    47,    -3,   -52,    -3,     8,    70,    27,    23,     4,   -10,     9,     8,    24,     8,   -39,  -115,  -143,   -84,   -13,    14,     2,   -91,   -68,   -43,     0,     7,     0,     9,   -14,    14,   -13,   -30,     2,    28,    26,   -41,    -4,   -14,    -2,   -34,    22,    22,    -9,   -81,   -77,   -11,    22,    26,    54,    75,   -29,   -47,   -13,     0,     0,    -3,   -26,    -1,   -58,   -26,    15,    -1,     2,   -11,    31,    27,    -3,     7,   -38,    10,    -4,    13,    30,    38,    67,    85,    79,    60,    -4,   -85,   -31,     1,    -1,    -6,    -3,   -36,   -95,   -59,     8,     5,    -5,   -12,    27,   -12,    -7,     3,   -11,   -29,    -3,    14,    23,    23,    -5,    49,    38,     0,    15,    -5,    25,    -4,     8,     7,   -35,   -58,   -17,     5,    15,    11,    -7,   -19,    -7,    -6,   -37,   -77,   -57,   -38,   -56,   -45,   -28,   -24,   -15,    29,    39,    37,    41,    -2,    13,    -4,    -4,    -1,   -28,    14,    31,    27,     5,    13,     1,   -21,    24,   -27,   -54,   -56,   -39,    19,   -27,   -59,   -36,   -38,   -13,    32,    30,    56,     0,     8,    15,    22,    24,     3,     1,    -9,     1,    -5,    10,     7,   -15,   -16,    -6,   -20,   -10,   -18,    12,    30,    22,   -31,   -27,   -40,   -18,    10,    57,    47,    22,     6,     8,    30,    23,     3,     3,    12,    53,    16,    -2,    14,    30,   -17,   -27,   -44,    -4,   -37,    33,    41,    -1,   -34,   -43,   -39,   -39,     5,     8,    10,     2,    11,     3,     1,     1,   -14,    26,     4,     3,     4,     2,    43,    24,   -14,   -38,     9,    17,    20,    35,    13,   -22,   -28,   -35,   -16,    -3,    -6,    -9,    26,    51,    61,     5,    -2,     3,     7,    17,   -46,   -34,   -47,   -62,   -12,    38,    -9,   -27,    35,    56,     6,     6,    -4,     2,     0,   -15,    -1,     7,    10,     7,   -31,     7,     1,     6,    -1,    -4,     9,   -21,   -39,   -39,   -13,   -83,   -20,    17,   -16,    13,    43,    12,   -61,   -37,   -31,   -55,   -32,   -19,   -11,   -30,   -23,   -19,   -21,    -6,     0,    -5,    -2,    -9,    -3,    -5,   -37,   -29,   -30,   -44,   -57,   -47,   -32,   -16,   -30,   -30,   -24,   -26,   -37,   -40,   -16,     2,    -5,    -6,    -4,    -5,     4,    -2,    -9,    -7,     6,     0,    -9,     5,    -3,    -5,     2,     3,     5,    -7,   -31,   -14,    -8,    -5,   -19,   -10,     8,     3,    -9,     0,     0,     0,     7,    -6,    -4,    -5,    -8,     8),
		    12 => (   10,    -8,     9,    -6,     1,    -2,    -2,    10,     3,     6,    -7,     7,     6,    -8,    17,    10,   -10,    -6,     4,    -3,     3,     4,    -6,    -7,     3,     2,     6,    -5,    -9,    -8,    -7,    -5,     0,     0,     2,   -14,   -32,   -12,   -14,   -18,   -16,   -27,    -8,     8,    10,    -4,   -10,   -31,   -20,   -17,    -3,     9,    -1,     4,   -10,    -3,     8,    -3,   -13,   -29,   -21,     7,    -3,   -10,     2,     7,    11,    33,    10,   -15,   -13,   -29,   -35,   -20,    11,    11,     5,     6,   -27,   -10,   -16,     7,     7,     7,     0,     9,   -12,   -58,     2,   -29,   -14,   -28,    -3,    30,    57,    41,    32,     7,     2,     5,    -1,    -1,   -15,     1,     6,    10,   -28,   -50,   -26,   -24,    -7,     4,     0,    -3,    -3,   -23,     7,    17,    36,    50,     4,    -2,    14,    45,    41,    50,     1,    -7,    -2,   -23,    -5,   -34,   -18,   -28,   -32,   -31,   -54,   -44,   -43,    -9,    10,     7,   -34,    -5,     3,    20,    37,    68,    33,    17,    15,     4,    12,    11,   -22,   -16,   -24,   -17,   -22,   -10,     4,     9,   -13,   -26,   -46,   -21,   -24,    -9,   -10,    -6,     1,     0,    -6,     2,    48,    39,    26,    25,     9,     2,   -13,    -2,   -16,   -22,   -16,   -15,    -6,   -28,    -4,    12,     7,   -30,     0,    44,   -23,     3,     7,    -8,    -4,    -4,   -12,     9,     2,    13,    -1,   -25,   -19,     0,   -14,   -21,   -12,    10,    11,   -32,   -29,   -36,     5,    20,   -11,   -32,    14,    52,   -68,   -28,   -29,    20,   -13,     2,    -8,     2,   -12,     6,   -34,   -42,   -21,   -24,    -6,     4,    -2,     6,     8,   -10,   -23,   -11,    -8,    -3,   -10,    13,     8,    -5,   -63,   -32,     5,   -27,    33,     1,   -15,   -11,   -22,   -17,   -28,   -37,   -19,   -24,    -4,   -10,    35,     7,   -25,    -9,   -20,   -15,    -5,    12,    11,    -2,   -18,   -36,     0,   -23,     7,    -5,    10,    -9,   -33,   -13,   -24,   -42,   -60,   -52,   -58,   -21,    -7,   -17,   -15,     1,   -36,   -10,   -39,   -10,   -34,    13,    20,   -19,   -39,   -16,    18,   -35,    -4,   -21,   -12,   -34,   -26,   -20,     2,   -56,   -60,   -59,   -55,   -19,    -5,     7,    16,   -14,   -40,   -26,    12,    -5,   -17,   -16,   -11,   -15,   -27,   -14,    -1,   -15,    -5,   -14,   -35,   -39,   -15,    -7,   -26,   -32,   -13,   -16,   -15,     8,    28,    -1,    -5,   -10,   -21,   -13,   -21,     3,   -36,   -39,   -15,   -33,   -42,     2,    17,     9,     7,   -13,   -21,   -25,   -27,   -42,   -15,   -37,   -25,   -11,     1,    -8,    -2,    -6,    -7,   -12,   -26,   -22,    10,     0,   -14,   -15,   -29,   -34,   -10,    12,    33,     1,    -2,   -24,   -17,   -10,   -31,   -46,    -9,   -29,   -21,   -24,   -21,   -36,   -34,   -22,   -19,   -28,   -35,   -38,     3,    -9,    -8,   -43,   -32,   -30,   -10,    25,    43,    26,     2,   -29,   -20,     2,   -24,     4,   -23,   -16,    -2,   -25,   -13,   -19,   -29,    -4,   -10,   -30,   -57,   -41,    -3,    -2,     4,   -17,   -30,   -37,    16,    40,    52,    38,     4,   -15,    -6,    29,    26,    -1,   -15,   -19,   -11,   -10,    10,     3,    10,    10,     6,   -20,   -31,   -29,   -34,   -23,   -15,   -12,   -24,   -30,     4,    31,    62,    41,    -9,    -9,    10,    31,    27,    -8,    -4,   -35,   -16,   -10,   -18,   -17,    27,     6,   -17,   -18,   -38,   -36,   -22,   -36,   -42,   -25,   -26,   -46,     0,    50,    41,    48,     8,     1,   -10,     9,    32,     1,   -33,   -14,     0,     6,    -4,   -27,    -1,    -7,    -1,    -6,   -42,   -17,   -35,   -29,   -14,   -16,     4,    -1,    31,    29,    31,    37,     2,    -3,    -2,    13,     7,   -17,    -5,   -14,    -6,   -17,     7,    11,     2,     3,   -23,   -19,    -4,   -12,    21,   -49,   -20,    13,    24,    36,    37,    39,    68,    74,     3,   -14,     7,    -5,    15,    14,   -11,   -12,   -18,    -2,     3,    25,    -2,   -14,   -20,   -26,   -12,   -19,    19,   -32,    -6,    19,    30,    41,    46,    25,    21,    -8,     5,     4,    16,    21,   -13,     7,    -3,   -22,   -30,   -24,   -22,    -8,   -22,   -15,   -26,   -15,    -5,     7,   -11,   -20,    11,    23,    45,    42,    21,    -6,     7,   -14,    -1,     5,     4,    12,    21,   -14,    -7,   -18,    -8,   -16,   -30,   -16,   -10,   -10,    14,   -19,    15,   -14,   -24,    -1,     5,    17,    40,    38,    11,    29,   -32,   -16,    -2,     4,     4,    11,     9,     0,    -6,    -1,    15,   -20,   -11,    20,     2,     8,    13,    11,     1,   -29,   -38,   -28,     6,    17,    42,    50,     1,    23,   -16,     6,    -4,     9,   -21,   -10,   -20,   -23,   -22,    -4,   -11,    -8,   -27,     1,    20,     1,    25,    -1,   -29,   -20,   -21,    -1,   -25,   -10,   -26,    18,    13,     7,     2,    -2,    -7,     4,   -36,    -9,    -5,    -6,     2,    -7,   -24,   -33,   -35,   -11,   -30,   -55,   -21,   -25,   -39,    -6,   -26,    -1,   -26,   -24,   -29,   -19,   -13,    -6,     2,     8,     0,     9,     1,     5,   -17,   -32,   -21,   -25,   -30,   -44,   -40,   -19,   -15,   -27,   -51,   -39,   -80,   -86,   -74,   -60,   -31,   -23,   -40,   -27,     3,    -3,    10,   -10,     5,     3,     5,    -3,    -1,     6,   -11,   -14,   -22,   -12,   -23,   -28,   -14,   -44,   -27,   -26,   -30,   -26,   -35,   -13,   -22,   -15,   -23,     8,     2,    -4,   -10,     9),
		    13 => (   -4,   -10,     9,    -4,    -7,     3,   -10,    -9,     9,     4,     7,    -7,   -10,   -10,    -3,     0,     7,    10,    -3,     4,     9,     5,    -5,    -9,     5,    -2,    -3,     4,     4,     3,    -7,     7,     2,    -4,    -8,    -3,     8,    -1,    -6,     5,     0,    -5,   -15,    -9,   -19,    -5,     7,    -4,    -7,    -1,    -6,     4,    -4,    -7,     9,     2,     4,     4,     1,    -4,     7,    -5,     5,    -1,   -23,   -43,    34,    22,    39,   -14,   -16,   -21,   -11,     2,    -5,    -4,   -21,   -14,   -31,   -17,     1,     0,     3,     8,     0,     6,    -4,     4,     2,   -15,     8,   -13,   -25,   -39,   -48,   -31,   -39,   -99,  -142,  -110,   -89,   -12,    12,    -2,   -37,   -31,   -25,   -45,    -5,    -6,     0,    -9,    10,    27,     2,    15,   -36,   -45,   -28,   -21,    43,   -27,    24,    45,   -36,   -22,     1,   -12,   -38,    32,    10,   -37,   -16,    27,   -18,   -19,   -36,   -18,   -14,    -1,     7,    -2,    39,     0,    51,    61,    34,    27,   -25,   -39,    -1,    -1,    -6,   -15,     7,    -1,   -22,   -17,   -11,    -8,   -54,   -51,   -25,   -45,   -17,   -43,   -22,    -9,    -3,    -1,    10,    16,    43,    49,    15,     2,   -19,     0,    -4,    33,     0,    29,    16,     9,    -4,    23,     2,   -94,    -5,   -31,   -66,   -35,   -15,   -18,    -4,    -9,    -7,     9,    17,   -24,    60,   -23,    54,    17,     7,    29,     5,    20,     4,    19,    18,   -46,   -25,    -1,     7,   -24,   -16,     0,   -63,   -42,   -27,   -24,   -30,   -10,    -4,    -8,    15,   -25,    55,    11,     8,    17,     0,    67,    36,    20,   -16,    -6,   -24,     0,    -3,    16,    26,   -20,   -41,     3,   -36,   -95,   -58,   -18,   -41,     8,     7,   -27,    35,    16,    42,     4,    63,    72,    33,    33,    -2,   -58,   -43,    -7,     8,    23,    -2,     5,     5,    21,     9,   -15,   -69,   -71,   -77,   -29,   -21,     0,     7,   -34,    40,    61,    52,    30,    35,    19,   -62,   -90,  -123,   -62,   -49,    12,    18,    39,   -10,    59,    -4,     7,     9,   -21,   -52,    -2,   -41,   -28,   -25,     3,     7,   -21,     4,    58,    22,   -31,   -59,   -98,  -155,   -82,   -17,   -20,    26,    53,     5,    -5,   -31,   -25,    11,    -5,    16,    -3,   -70,   -50,   -28,   -24,    -7,    -2,    -6,    -5,    48,    55,   -35,   -78,  -127,   -77,   -77,     7,    44,    28,    41,    32,     8,   -28,   -48,   -38,   -38,   -78,   -49,  -101,   -50,   -78,   -34,    -1,     2,   -14,    -8,     4,   -14,   -17,   -11,   -50,   -78,   -62,   -31,     4,    40,    13,    21,    13,    11,   -37,   -15,   -27,   -44,   -43,   -59,   -65,   -26,   -18,   -16,   -33,   -26,   -15,   -10,    18,     4,    25,     1,   -37,   -45,   -27,    47,    -2,    13,    -5,     7,    -3,    30,   -16,   -15,   -20,   -54,    13,   -37,   -34,   -39,    17,    -5,   -76,   -37,   -19,   -16,    17,    15,    41,   -24,   -34,   -18,   -12,    -7,    23,    39,    73,     1,     9,    12,    21,    -2,   -41,   -45,     1,     3,    36,   -43,    49,    -6,   -38,   -15,   -25,    10,     7,    19,    38,   -44,   -60,   -35,   -25,    16,    50,     1,     2,    39,    35,    29,   -11,     3,    -7,    -2,   -27,     9,    57,    24,    29,    -9,   -55,   -57,   -24,     5,    12,    20,    41,   -47,   -86,   -85,   -73,   -32,   -18,   -52,    -8,     9,    25,     4,     5,    25,     5,    -7,     9,   -19,    45,    48,     5,   -26,   -86,   -39,   -16,   -14,    -2,    35,    69,   -16,   -49,   -70,   -90,  -144,  -191,  -158,  -167,  -159,  -120,   -81,  -106,   -27,    65,     6,    20,    21,    16,    73,    40,   -29,   -68,   -34,   -28,    -1,   -12,   -58,    37,    31,    36,   -30,   -35,   -60,   -85,  -129,  -140,  -127,  -109,   -87,   -98,   -52,   -23,     9,    44,    41,    31,    47,    53,   -10,   -45,   -57,   -30,     4,    10,   -40,   -23,   -10,    37,    14,   -11,    -4,   -44,   -45,   -38,   -31,    -8,   -12,   -52,   -60,   -10,    -2,    31,    27,   -10,     7,   100,    -6,   -44,     3,     3,    -5,     5,    27,    30,    22,    -4,    30,    18,    -5,   -12,     5,    -2,    20,    25,   -18,   -10,   -25,    -4,    18,    11,    46,   -26,   -28,    -9,   -35,   -40,   -12,     5,     8,    -7,    42,    38,    54,    32,    16,    26,    46,    18,    -5,   -21,    -3,    25,   -32,     4,    -6,   -31,    12,     7,    21,    16,    -2,    18,   -67,   -48,     1,    -7,    -2,     4,    42,    56,    51,    -5,     2,    20,    17,    11,    -9,    22,   -20,    18,   -19,   -14,   -20,   -20,   -52,     0,   -39,   -16,   -40,    -2,   -44,    -7,     8,     9,     9,     9,    14,    -7,    61,    39,    16,    57,    40,     0,    42,    32,    18,    -7,    11,   -20,   -25,     8,   -12,   -38,   -64,     3,    26,     6,   -42,     2,    -2,     1,     9,     2,   -10,   -35,    13,    47,    11,    24,    38,    21,    -9,   -23,   -33,   -43,   -55,   -35,   -12,   -61,   -63,   -62,   -44,   -37,   -21,  -110,   -47,    -9,    -7,     2,     7,     0,     9,   -25,     3,     2,   -33,   -14,   -45,   -53,   -60,   -62,   -53,    20,   -19,   -40,    44,    -2,    11,    -9,    -6,     4,   -31,    -5,    -3,    -8,     6,     1,    10,    -9,    -2,    -5,   -11,     7,    -7,     7,    -2,   -49,   -36,   -26,     3,   -33,   -20,   -24,   -12,    -2,   -15,   -36,   -41,    -7,   -18,    -6,    -3,    -7,    -9,     3),
		    14 => (    0,   -10,     7,    -7,     6,     7,     5,   -10,     1,    -6,    -1,     1,   -27,   -18,     0,    -3,     3,    -9,    -4,    -8,     7,    -1,    -6,    10,     9,     6,     6,     6,     3,    -3,     7,     6,     4,     0,    -1,   -18,    -8,   -13,   -30,   -28,   -38,   -25,   -10,   -84,   -69,   -54,   -15,   -12,   -31,   -16,    -9,    -7,    -6,    -3,     0,     7,     7,   -10,    -3,   -30,   -84,     2,    -7,   -27,   -47,   -34,   -68,   -66,   -68,    -2,    16,    17,   -65,   -44,   -22,   -22,   -63,   -32,     6,    -4,    -7,   -42,    -1,    -7,    -2,     1,     2,   -29,   -84,   -65,   -28,   -13,   -15,   -25,   -61,   -65,   -44,     3,    24,     3,   -49,   -61,     1,    31,    44,    35,   -17,   -42,   -66,   -35,     4,     0,     6,    -4,   -12,   -58,   -25,   -31,   -17,    14,    26,    37,    -4,   -64,   -66,     4,     6,   -11,   -18,   -19,    24,    -6,    36,     8,    -5,   -33,   -64,   -39,   -48,    -7,     1,     7,   -23,    -9,   -22,     0,    25,    16,    41,    22,    -6,   -54,   -55,   -36,    -2,   -25,   -43,    10,    12,    28,    -4,    -7,     2,    -2,   -19,    23,   -53,   -14,    -5,     1,   -41,   -16,    26,    29,     7,    12,     1,   -23,     5,   -21,    25,    20,    47,    96,    96,    72,    45,    40,     8,    46,   -24,    -6,   -13,   -29,     3,   -22,    -2,   -72,   -18,    12,    15,    19,    45,    44,     2,    16,    19,    -5,    24,    28,    25,    63,    72,    57,     7,   -11,     2,    -2,     4,     4,   -20,    12,   -10,   -73,   -34,   -84,    -8,     5,     3,     6,    52,    34,    42,    -9,   -38,    -6,   -21,    -3,   -16,     9,     3,   -17,     1,     1,    -9,     6,    -8,    -4,    13,    27,    -5,   -62,    -4,   -37,   -44,     4,    -1,    11,    -3,    -6,    -7,   -63,   -64,   -11,   -35,   -56,   -67,   -31,   -24,   -26,    -3,   -27,     3,    27,     7,    10,   -22,   -12,   -23,   -47,     3,   -31,     7,    -2,   -22,   -15,   -31,   -23,   -35,   -38,   -25,   -24,   -32,   -81,   -91,   -58,   -49,   -32,     7,   -15,   -35,    35,   -14,   -64,   -77,   -48,   -28,   -14,    -2,   -28,   -24,     1,   -35,     1,   -31,   -16,   -38,   -37,   -30,   -38,     2,   -33,   -73,    -7,   -28,    12,    12,    19,   -14,    18,   -31,   -94,   -89,   -59,   -39,   -60,    -6,     4,     6,    16,   -19,    13,    24,    -5,    20,    21,    24,     8,    34,    27,   -43,    20,    16,    -3,    -3,    16,    23,    73,    17,   -20,   -54,   -34,   -70,   -75,    -6,   -13,   -31,    -2,    38,    -8,     1,    -6,    25,    16,     3,    34,    20,   -12,    13,    56,    28,    32,    35,    41,    27,    17,   -14,   -14,   -56,   -25,   -53,    -3,    -6,   -14,   -83,   -17,    38,   -12,    -9,    -4,    -9,     0,   -29,   -11,   -38,   -14,     9,    53,    15,    36,    54,    37,    41,    11,     2,   -23,     5,   -32,    48,     7,     5,     2,    42,    11,    29,   -51,   -23,     1,   -14,   -36,   -78,   -46,   -28,    25,    43,    75,    68,    59,    58,    -7,     2,    13,    17,   -17,   -41,   -45,    50,   -41,     4,    -2,     7,    26,    29,   -36,   -38,   -21,   -27,   -47,   -63,    -7,    12,    58,    85,    69,    81,    20,    52,   -20,     4,    -8,   -16,   -24,   -20,     7,     5,   -17,     9,    -3,    20,   -17,    60,   -47,   -20,   -23,    -5,   -45,   -11,    22,    60,    57,    51,    58,    81,    25,    38,   -32,   -16,    -7,     7,     3,   -32,     6,    34,   -42,   -54,    -9,    -2,    -8,    50,   -33,   -21,   -27,   -88,   -20,    12,    20,    44,     8,    52,    49,    57,    19,    -5,   -40,     8,     5,    -9,    57,   -48,   -59,   -16,    -7,    -2,   -14,   -33,    38,    -3,   -10,     3,     3,    -6,    20,    26,    67,     1,   -33,    28,    29,    -4,   -26,    30,    12,   -15,    10,    -5,    -4,   -36,   -29,   -19,    -7,     7,     5,   -17,   -34,   -56,   -46,   -35,     6,    41,    32,    41,    39,    34,    36,    -9,    15,    58,     6,    42,    21,    33,    13,     7,    -3,   -48,   -72,   -41,     2,    -8,   -14,   -53,   -26,   -65,    -7,   -72,    -4,    20,    13,     3,   -23,   -51,   -48,    52,    36,    20,    15,    -8,    20,    15,   -15,    23,    10,   -16,  -107,   -62,     3,   -10,   -15,   -10,   -44,  -132,   -62,   -13,    -9,     7,   -65,     5,   -21,   -29,   -15,   -12,    28,    -3,   -42,   -18,    17,   -10,    21,     2,    23,   -32,   -55,   -24,   -18,     2,     0,    -2,   -73,  -112,   -99,    30,    -3,   -43,   -46,   -20,   -32,   -34,   -15,    15,   -16,   -20,   -19,    11,    38,     6,   -18,   -37,    -5,   -25,    -8,   -14,    -6,     7,     0,   -12,   -14,   -80,    14,    -3,   -28,   -54,   -43,   -48,   -28,   -23,     6,    -7,   -28,     3,   -25,     2,    54,   -33,   -46,   -13,    12,   -51,    28,   -37,     5,     2,    10,    -3,    -4,    52,    38,   -47,   -55,   -45,    -2,   -49,    14,    -4,    29,    14,    12,    -6,   -38,   -22,   -13,   -47,   -61,   -21,    23,   -14,   -40,   -39,    -7,    -9,     6,     8,   -39,    55,     5,   -32,   -76,   -45,   -41,   -51,   -32,   -89,   -68,   -77,   -80,   -54,   -78,   -60,   -29,   -84,  -127,  -134,     3,    -4,    -4,    -8,    -2,     5,     3,    -5,     3,    -7,   -15,   -19,   -34,   -39,   -38,   -70,   -54,   -40,   -45,   -79,    -9,   -43,   -57,   -34,   -47,   -55,   -44,   -53,    -4,    -6,    -3,     4,     6),
		    15 => (   -3,    -9,    -1,    10,    -7,    -4,     3,    -8,     8,     9,    -3,     0,     3,    -2,    -2,    -4,    10,    10,    -4,    -3,    -9,    -4,     6,    -1,     2,    -8,    -1,    -5,    -6,    -1,    -4,     0,     8,    10,    -9,     6,     9,     1,    -8,   -10,   -21,   -25,   -22,   -15,   -21,   -39,   -21,   -15,   -18,    -9,     4,     3,    -2,   -10,     0,    -8,   -10,   -10,    -7,   -12,    -6,     7,   -12,   -29,   -26,   -55,   -25,    -9,   -24,   -43,   -51,   -68,   -29,   -17,     5,     0,   -13,   -30,    -7,     5,   -16,   -11,   -10,    -5,     2,    -3,   -19,    18,     8,   -21,    -1,   -42,   -43,   -42,   -44,   -22,   -18,   -46,   -47,   -72,   -84,   -46,   -19,    -9,    -9,    15,    14,    -9,   -21,   -25,     5,    -8,    -8,     2,   -12,    13,   -12,   -10,    -5,    17,   -18,    11,   -42,   -35,   -57,   -59,   -11,    15,   -43,   -18,   -24,   -17,   -39,    -9,   -24,    18,    21,   -25,   -44,   -45,     2,    -8,   -13,    -1,    -7,    11,    26,    21,   -40,   -37,     9,    -9,   -29,   -52,     6,    15,   -14,   -32,   -30,   -24,     9,   -10,   -44,   -63,   -48,   -11,   -22,   -31,     6,   -11,    -5,   -26,   -19,    24,    19,    -7,   -28,   -32,   -23,     9,   -19,    -4,    35,   -26,   -42,   -56,   -45,    -5,    -6,   -22,    -4,    -9,   -27,    -3,    -2,    33,     6,   -13,   -12,   -37,    -8,     9,     9,   -25,   -32,   -53,     8,     5,   -19,   -36,    14,   -34,   -51,   -50,   -99,   -92,   -80,   -30,    -5,   -14,    14,    12,    13,    25,    -3,   -44,   -42,   -44,   -32,    37,     1,   -14,   -64,   -18,    25,   -31,   -12,     3,   -41,   -81,   -44,   -35,   -80,   -74,   -40,   -34,   -33,    -9,     4,   -33,   -75,    -1,    -2,    -9,   -15,   -38,   -22,    31,   -32,   -60,   -22,    -4,    16,     0,     3,   -67,   -16,   -59,    17,    17,    21,   -22,   -29,    -3,   -17,     8,    47,    14,   -17,   -12,    -6,   -16,    -4,    -8,   -35,   -15,    -3,   -47,    -8,    -6,    21,     3,   -14,    32,   -10,    13,    46,    47,    52,    53,    42,    23,    30,    89,    57,    74,    17,   -14,     4,    -8,   -11,   -12,   -19,   -23,    26,   -24,    -3,     7,    19,    42,     5,   -13,   -12,   -11,    40,     3,    29,    35,    62,    73,    81,    87,    22,    38,     3,     1,    -7,    -2,    -5,   -30,   -52,   -19,    -5,   -17,    -6,    43,    41,     7,    14,    -1,    26,     4,   -15,    -9,     2,    14,    72,    37,    61,    44,    10,    38,    82,   -10,    -6,    -5,    -6,   -15,   -64,   -13,   -35,   -30,    16,    12,    34,     9,     7,    -9,   -22,   -69,   -15,   -10,   -99,   -62,   -39,   -53,    -8,   -20,    -8,     4,    73,   -22,     0,    -5,   -21,   -49,    31,    24,   -10,    -4,    43,    16,    21,    49,    20,    28,   -64,   -69,   -56,   -50,   -33,   -70,   -24,   -37,   -17,   -34,   -43,   -49,   -25,     3,    11,     8,   -14,   -27,    70,    -4,    14,    -8,   -14,    28,    -7,    10,    49,    -4,   -48,   -37,   -62,   -63,   -19,   -45,   -30,   -21,   -28,   -47,    -6,   -71,   -14,   -20,   -13,   -17,   -18,    -3,   -59,   -38,   -62,   -23,   -46,   -30,   -15,   -15,     3,     0,   -16,    -8,    -5,    -3,    -7,   -40,   -50,   -14,   -50,   -12,   -25,   -63,   -33,   -23,    -8,   -10,   -15,   -24,   -36,   -51,   -56,   -84,   -71,   -14,   -62,    -2,   -14,   -46,     6,    -4,   -22,    -5,    -2,   -19,    -3,   -16,   -66,    31,   -42,   -75,   -40,   -67,    -7,     1,   -14,     9,    -4,    -8,    -1,   -14,   -51,   -28,   -25,    19,    16,   -30,   -46,   -54,    30,    16,     5,   -32,    -7,   -29,   -30,    18,   -28,   -17,   -43,   -35,    -3,    -8,    20,   -42,    -9,   -42,    28,    25,   -32,   -18,    -6,     8,   -16,     0,    19,     7,    38,     7,    23,     4,   -16,   -41,    13,    37,   -16,   -50,   -46,   -39,    -5,   -25,    15,   -42,   -32,   -22,    23,    39,    -6,    17,    35,   -22,    -7,    11,   -30,     3,    30,    26,   -13,   -11,   -32,    12,    33,     8,   -13,    -3,   -59,     9,     1,    -8,    -7,    -3,   -30,    15,    41,    45,     7,    -1,    10,   -27,   -43,    17,   -35,    14,    13,    -4,    31,     5,    27,    22,    -2,    -4,   -47,   -10,   -46,    -7,     1,     7,    -8,    25,    -5,   -12,    16,   -13,    22,     3,    22,    20,    44,    14,    23,    23,     4,    17,     0,    17,    27,     8,   -16,    -7,   -41,    -3,   -17,    -4,     2,     5,    21,   -18,   -35,   -47,   -16,    -9,    36,    15,    17,     8,    27,    53,    34,   -19,    -7,     6,   -31,    17,    23,   -17,   -32,     4,    -3,     2,    -8,    -2,   -10,    -6,   -21,    -4,    -6,   -44,   -44,   -41,    35,    39,    28,    13,     6,   -13,    31,    12,    10,    34,   -16,    13,     6,   -44,   -21,    12,    -4,   -46,   -13,     9,     2,    -9,    -9,     8,   -24,   -61,   -31,   -71,   -45,   -66,   -44,   -31,   -42,   -58,   -40,   -25,   -50,   -67,   -43,   -33,   -17,   -13,   -17,    -9,    -4,    -5,     9,    -7,    -2,     7,    -6,   -12,    -9,   -43,   -54,   -51,     1,   -22,    13,   -14,   -40,   -74,   -67,   -70,   -57,   -31,   -45,    -9,   -13,     7,     1,   -25,    -1,     7,     4,    -8,     8,    -6,    -4,    -9,   -14,    -1,    -9,   -14,     1,     3,     2,    -5,   -11,   -12,   -59,   -28,   -20,    -5,    -5,   -23,   -29,   -39,   -38,   -12,    -7,    -5,     0,    -6),
		    16 => (    5,    -9,     8,     0,     8,    -4,    -5,     1,    10,    -1,    -1,    -4,    15,     3,    -6,     1,    -2,    -5,     8,     7,    -2,    -2,     2,    -7,    -3,    -3,     6,    -9,    -2,     3,     4,    -6,     5,    -7,     2,    28,     9,     7,     9,    11,    35,    16,   -27,     3,    15,    14,     6,     2,    44,     8,    14,     9,     6,     2,    -1,    10,    -4,    -4,    18,     4,    10,    12,    19,    22,    22,   -13,   -16,    -4,   -36,   -28,    16,    13,    60,    68,     7,   -34,   -46,    24,    40,    28,    13,   -12,     1,    -1,    -8,     0,   -11,    -2,    15,    30,    -7,    -4,    -1,   -19,   -15,    -7,   -43,   -13,    30,    34,    62,    26,   -11,    13,    55,    26,   -23,    -8,     4,     1,    -3,    -9,     7,     3,   -29,   -27,    50,    45,    -9,   -11,   -26,   -15,   -14,   -40,   -45,   -19,   -40,     3,   -10,     2,   -26,   -12,     4,   -39,     6,   -35,   -31,   -17,    24,    23,     7,    -2,   -19,    -4,    55,    49,     6,    -5,   -10,    -4,   -52,   -83,   -28,   -51,   -12,   -14,    24,    23,   -15,   -11,   -64,   -53,    -5,   -36,    -7,     0,    21,    10,     5,    -1,     5,   -26,    34,    28,    -6,    -1,   -13,   -25,   -71,   -78,   -48,    -9,    11,    43,     4,   -45,    24,    21,   -10,   -63,   -11,   -13,     3,    -5,    -9,    12,     8,    -4,    -1,   -49,    25,    34,    -3,   -25,   -20,   -32,   -58,   -77,   -44,     3,     8,   -58,   -35,   -61,   -36,     5,     6,    24,    27,     4,    -8,    14,     5,   -15,    -2,     3,    -7,   -49,    27,    31,     7,    -2,   -30,   -37,   -55,   -82,   -20,     9,     9,   -41,   -22,   -37,   -57,   -39,   -17,    44,    17,   -14,   -11,    -4,   -34,   -47,     5,     0,    -3,   -23,    47,    37,     6,    13,   -17,   -39,   -43,   -10,    15,    21,   -10,     8,   -40,   -27,   -46,   -40,   -39,   -37,   -35,     3,    -9,     3,     1,   -14,     9,    -8,   -16,   -30,    45,    49,   -12,   -17,   -27,   -12,    -8,   -31,    22,     0,    -3,   -65,   -40,   -46,   -82,   -60,   -49,   -56,   -30,     4,     9,     3,   -15,    -8,    -5,     6,     2,   -35,    57,    54,   -10,   -14,   -27,   -45,   -34,    10,    -4,   -21,   -33,   -46,   -30,   -55,   -75,   -61,   -41,   -62,   -47,    10,    15,     5,   -11,   -23,     4,    -2,    -9,   -26,    31,    46,   -15,   -33,   -32,   -16,    -5,    43,    14,   -24,   -18,     0,   -45,   -69,   -48,   -27,   -22,   -55,   -46,    30,    25,     0,   -29,   -21,     4,     2,    10,   -24,    34,    33,    -2,   -21,   -17,   -24,    -4,    21,    -5,    -5,    11,    16,    44,    13,   -24,   -23,   -14,   -42,   -37,    15,   -30,   -38,   -28,     0,     7,     7,    -9,    -7,     0,    26,    20,     5,    -7,   -54,     1,    -3,    -2,   -16,   -29,    -8,    35,   -27,   -45,     0,    25,   -32,   -35,    -7,   -17,   -18,   -19,   -11,    10,    -1,   -10,   -29,   -10,     7,    12,     0,   -21,   -38,    -2,     3,    -2,   -69,   -11,   -11,    12,    45,    -1,    46,    37,   -27,    -8,   -15,   -27,   -27,   -14,   -38,    -5,     9,    -6,   -31,   -12,    13,    -3,    21,    18,   -40,    -4,    51,    43,   -39,   -11,   -47,    -8,    12,   -28,    25,    -3,   -42,   -19,   -33,   -16,   -10,   -20,   -16,     4,    10,     4,   -34,   -22,   -10,     7,    12,    15,   -41,    27,    64,    16,   -71,   -64,   -24,     7,   -28,    -5,    20,    -3,   -34,   -29,   -15,   -27,   -51,    -9,   -28,     9,     1,    -1,     8,   -26,     0,     0,    -1,   -46,   -35,     1,     7,    27,     2,   -53,   -39,     1,    18,    14,    18,   -53,   -32,   -46,   -38,   -47,   -53,    -8,   -27,     4,    -4,     2,     2,   -13,   -24,   -29,   -30,   -34,   -47,    -5,    53,    30,    32,    -1,   -18,   -33,    25,    11,    11,   -31,   -21,   -41,   -36,   -38,   -28,   -29,   -12,     6,    -6,    -8,    -8,    -1,   -15,   -24,   -38,   -42,   -64,   -55,    -5,    15,    35,    -7,     2,   -12,    38,    -6,    20,    13,   -22,   -18,   -20,   -14,   -15,    -5,     1,    -4,     2,     5,    -4,     8,    -8,   -13,   -27,   -36,   -57,   -53,   -53,     0,    26,     3,    -9,   -20,    -9,    -1,    -4,   -45,   -25,   -15,   -11,   -22,   -27,    -1,     6,     7,     1,     0,   -13,     3,    -9,     9,     0,   -28,   -64,     7,   -21,    -1,     8,    30,    32,   -21,   -47,   -52,    16,   -10,   -14,     5,   -13,   -39,   -11,     7,     4,     6,    -8,    -5,   -13,     5,    -5,     0,   -10,   -11,   -41,   -49,   -29,     7,   -14,     4,   -14,   -17,   -21,    -5,     5,   -19,   -15,     5,    -4,    -4,   -12,     8,     2,     9,     5,    -1,   -10,   -13,   -15,   -12,    -1,   -23,   -13,   -27,     8,    13,    15,     1,    43,    77,    32,   -51,   -76,   -21,    -2,    -2,    -4,    -6,   -13,     1,     2,     3,   -10,     1,    -9,     6,   -11,    -8,    -8,     2,   -14,    -9,     4,    22,    15,    -9,    -4,   -13,    -5,    -9,   -13,   -26,    -4,   -11,   -16,     2,     8,     6,     1,    -2,     5,     4,     3,    -5,    -3,     7,     4,     4,    -2,    -9,   -12,    -6,     4,     7,   -10,     1,     0,     4,    -9,    -3,   -16,     2,    -2,     9,     8,    -9,     6,    -4,    -5,     8,     8,     1,    -1,    -7,    -4,     5,    -7,    -3,     5,     0,     2,     3,   -12,    -7,    -1,     6,    -3,     2,     3,     4,    -7,     7,     0,     0,     0),
		    17 => (   -2,     2,    -7,     5,     0,    -6,    -8,    -9,     7,     6,    -7,     9,     3,    10,     8,    -7,    -1,    -7,     8,    -4,    -6,     4,    -5,    10,    -3,     1,     3,     6,    -5,     0,    10,    -1,    10,     8,     3,    -3,    -5,     4,    -8,   -40,   -36,   -25,    -6,   -31,   -33,   -25,     3,     4,     7,     5,     1,    -7,     9,     2,     4,    -2,    -2,     6,     3,   -22,   -16,     2,    -9,    -2,   -14,   -11,   -10,   -31,   -18,   -15,     0,   -23,   -25,    -4,    -4,     6,    -6,     3,    -9,     1,     8,     3,    10,    -3,     6,     0,     6,   -35,    -7,   -13,   -14,   -26,   -36,   -28,   -22,   -17,   -19,   -27,   -15,   -27,    -7,    -8,   -15,   -10,   -10,   -16,   -47,   -20,    -3,   -14,     9,    -7,     3,    -3,    -8,    -3,   -46,   -22,    -7,   -63,   -60,   -30,   -63,  -102,   -87,   -80,   -61,   -32,   -18,    -4,     3,    -7,   -39,   -48,   -27,   -50,   -13,   -22,   -12,     2,     7,    10,    -4,   -10,   -49,   -23,   -15,    14,    13,    -8,   -40,   -24,     6,     2,   -55,   -67,   -74,  -136,  -156,  -145,  -139,   -82,    -8,   -50,   -32,   -24,   -10,    -6,    -7,     7,    47,    51,    -4,    -8,    -1,   -26,   -25,   -46,   -65,    22,    37,    19,   -22,   -81,   -61,    -1,    -8,    -6,   -19,    49,    29,    11,   -36,   -40,   -66,   -20,    -7,    93,    85,    56,     7,    -8,    -1,    41,   -10,     0,     8,   -25,    21,    -7,   -29,   -42,   -41,   -13,    -5,   -14,   -31,     5,   -11,    24,    20,    -4,   -49,   -23,   -59,    99,    31,     9,   -20,   -33,   -25,   -10,   -43,    -6,    40,     4,    16,   -34,   -29,   -19,   -29,    19,    23,     3,   -12,   -35,   -15,    39,    63,    17,   -38,   -32,     5,    57,   -43,    -5,    16,     3,    24,    -9,   -23,     7,     8,    20,    10,     2,    44,    -3,   -29,    15,    33,    28,     5,    10,    10,    23,    69,   -10,   -64,    -2,     8,    43,    30,     7,    17,     9,    39,    16,    19,    -3,     3,    37,    37,    51,    -3,   -41,   -31,    14,     1,    27,    41,    35,   -28,   -19,   -30,   -22,   -53,    17,    -3,     9,    36,    46,    17,    55,    11,   -22,   -40,    41,    14,    68,    77,    -3,   -62,   -41,   -23,    -9,    55,    29,    39,   -14,   -35,     0,   -17,   -44,   -23,     7,    10,    13,    21,    30,     5,    29,    11,    42,    27,    20,    44,    23,    47,  -123,  -133,   -22,    20,    18,    30,     0,    16,   -17,   -40,   -40,   -25,   -32,    -5,    28,     1,    17,    46,   -12,   -10,    47,    32,    44,    35,    -6,     6,     4,   -27,  -168,  -113,   -59,    26,    -4,    31,   -27,     0,    19,   -36,   -66,    -3,   -53,   -14,    -8,   -10,    32,    88,    33,   -24,    52,    16,   -14,    -6,    34,    50,    11,   -78,  -220,  -101,   -37,    22,    -6,    44,    24,    -7,    -9,   -10,    -7,     3,   -33,   -24,    -6,    -9,     0,    23,    33,   -80,    20,    29,    26,   -36,   -22,    57,   -28,  -192,  -135,   -71,   -31,    27,    26,    18,    39,     2,   -15,     5,   -32,   -44,   -44,    -5,   -16,   -12,   -13,    14,    13,   -39,   -30,     7,    55,    -9,    -5,    61,   -82,  -186,   -24,     3,   -11,   -14,     8,    35,    31,   -38,    -4,    25,   -23,   -23,   -39,    -2,   -37,   -10,     5,    26,   -14,     7,   -27,     7,    -5,   -31,   -63,   -94,  -128,  -102,    -9,    13,    -7,   -12,   -22,    32,   -27,    10,    -5,    31,   -94,  -123,   -20,    -1,   -45,    23,    -8,    53,   -81,   -34,    -8,    19,     5,   -48,   -95,  -160,   -42,   -13,    26,    45,    -8,    17,    23,    23,   -26,    30,   -22,   -34,  -120,  -113,    13,    -1,   -14,    -7,    30,    20,   -65,   -10,    13,    16,  -101,  -101,  -117,  -124,   -41,    -4,     2,    11,    -2,   -14,   -24,    18,     1,   -19,   -48,   -75,   -88,   -55,    39,    -1,    -9,     1,    35,    -4,   -38,   -23,   -22,   -40,   -95,   -96,  -126,   -27,    46,    33,   -25,     1,   -33,   -21,     7,   -26,    -8,   -31,   -75,   -66,   -93,   -35,     1,    -4,    -3,    -6,     1,   -14,   -46,   -92,   -24,   -84,   -78,   -71,   -28,    64,    21,   -22,   -33,   -20,   -58,   -31,    -5,    26,     6,    -5,   -16,    -2,   -14,   125,     6,    -9,     4,     1,     9,    -9,   -24,   -59,     6,     5,     0,    10,    22,     4,    13,   -25,    -1,     5,     1,   -12,     6,    12,    24,     6,   -21,    -2,   -14,    -8,    -2,   -26,    -4,     5,     4,    -9,   -59,   -32,    34,    44,    28,    31,    -3,    16,   -64,     2,    20,    -1,     0,   -26,   -20,    22,   -40,   -20,    -8,   -85,   -55,   -10,   -18,    -8,    -6,    -6,     1,    14,    15,    -3,    42,   -17,   -48,    30,    -4,     8,    16,    11,    -1,    28,   -17,   -27,   -20,   -62,   -39,   -19,    13,   -69,   -69,   -16,   -58,     8,     3,     7,     0,    -7,    -2,   -70,   -89,   -33,   -24,    -1,    -8,    15,    12,    19,     4,    30,    -1,    18,    27,   -41,   -13,   -18,    18,    -3,   -45,    20,   -10,    -8,     5,     3,     3,     8,    -5,   -78,   -72,   -59,   -64,   -27,   -39,   -37,   -47,     8,    38,    42,     5,    26,   -11,     1,    18,   -17,   -20,   -12,     1,   -19,     6,     0,     3,     8,     9,     5,    -5,    23,    23,     9,    20,    39,    14,    21,    11,   -13,    -9,    10,   -20,   -23,    47,    43,   -37,    21,    70,    17,    37,    -5,     8,     1,     0),
		    18 => (    7,    -7,     2,     0,     7,    -1,     1,    -8,    -1,    -6,    -9,    -6,    -2,     8,    -4,     3,     4,     3,    -3,    -9,     3,     7,    -8,    -8,     1,     3,    -9,     4,     7,    -8,    -2,    -3,    -7,     8,    -6,    -4,     6,    -9,     4,     2,   -10,   -16,   -25,   -44,   -69,   -32,   -12,   -16,   -13,   -22,   -19,    -1,     7,     8,    -5,    -1,     8,    -2,   -13,     0,    -1,    -4,   -26,   -16,   -20,   -59,   -73,   -40,   -10,     3,   -13,   -50,   -32,   -12,    14,   -25,   -77,   -64,   -71,   -21,   -15,   -13,     7,     5,    -6,     4,   -30,   -31,     0,   -26,   -35,   -81,    15,     8,    -9,   -34,   -38,   -58,   -86,    -4,    12,     7,    29,    18,    72,    60,    27,    24,   -26,   -10,   -22,     2,    -1,     9,    -3,   -49,   -45,   -76,    -1,     0,   -32,   -51,     7,   -25,   -67,   -56,    28,     3,    11,   -10,   -10,    23,    53,    58,    33,    22,     1,    71,    31,   -12,    -9,     3,   -38,   -52,   -78,   -26,    -5,     5,    21,    -7,    -3,    -1,   -28,   -27,   -23,     8,     0,   -33,   -41,   -16,    51,    28,    13,    66,    67,    29,   -26,    -3,     3,     2,   -29,   -47,   -13,   -42,    11,    18,    20,    -6,   -15,   -27,    17,    -2,    11,    -2,   -46,   -49,   -16,    27,     2,   -23,   -48,    17,    -6,    81,     6,   -40,    -4,   -55,   -30,    -9,    -2,   -48,    19,    53,    -2,   -28,   -20,   -12,     4,    -1,     6,    19,   -47,   -10,    33,    14,   -26,     3,    23,    24,    18,    -6,    -9,   -45,   -18,   -15,   -30,    17,    53,   -20,    39,    41,   -37,    21,   -11,     7,     9,    43,   -20,   -66,   -28,   -21,   -25,   -54,     5,    47,    29,    -5,     9,    32,    27,    14,    -4,    10,    -8,    33,    16,   -47,   -21,   -14,   -22,   -16,    16,    39,   -14,   -15,   -48,   -67,    -2,   -10,   -38,    19,    19,    16,     7,    41,     9,    11,   -46,  -108,     5,   -11,   -14,   -33,    -4,   -46,   -33,   -54,    10,    29,    39,     9,    -9,   -38,   -42,   -40,     8,    41,   -15,   -20,   -12,   -17,     1,    27,     1,   -75,   -40,   -85,    -3,    -8,   -30,   -41,   -40,   -28,   -14,     6,   -23,    27,    -1,    46,    38,    -8,   -16,   -29,    -1,   -23,   -15,   -67,   -34,   -80,   -37,    37,    70,     7,    64,   -50,     1,     5,   -46,    52,   -27,    48,     5,    14,   -46,   -22,     1,   -34,    21,    37,    -8,   -28,   -31,    -1,    11,    30,   -48,   -12,    43,    85,    80,    24,    18,   -88,     0,    -2,   -44,    42,   -13,   -27,   -82,   -31,   -37,   -42,    -8,    -9,     8,    23,     5,    -8,   -54,    12,    -6,    22,    30,    68,    98,    85,    43,   -24,   -26,    14,   -15,    -1,    -1,   -72,     0,   -68,   -33,   -33,   -55,   -70,    -1,   -30,     0,    44,    13,     6,   -49,    36,   -46,    20,     1,    46,     8,    70,    42,   -24,   -59,    -1,    -1,     5,   -11,    27,    -8,    15,     5,   -20,     1,   -62,   -17,     8,    26,    12,    -2,   -20,    29,   -86,   -29,    13,   -31,   -62,   -15,    50,    52,     0,   -72,   -47,    -3,    -8,   -21,    35,   -50,    48,   -12,    11,   -39,   -46,   -23,    -6,    42,     8,    -5,    10,   -41,   -19,   -16,   -55,   -71,   -53,   -36,    25,    10,    19,   -54,   -41,    -1,    -7,   -23,    22,   -75,   -12,    -6,    31,   -23,   -37,     5,    32,    36,   -26,    40,    36,   -13,   -13,   -71,   -60,   -30,   -54,   -33,     0,    -7,     6,   -10,   -26,   -17,    -6,   -10,   -29,   -51,   -25,   -15,   -31,   -38,    38,    29,    55,   -27,   -88,   -17,    43,     1,   -10,   -20,    22,   -17,   -87,   -22,     3,   -55,     6,    -5,   -28,     3,    -8,   -21,   -20,   -59,   -23,   -22,   -52,    42,    14,    47,    44,   -41,   -83,   -38,    14,    10,    33,   -39,    -9,   -27,   -53,    -4,   -34,   -38,     1,   -35,   -14,     0,     8,   -11,   -26,   -90,    -9,   -44,    29,    22,    21,    40,    52,     8,   -23,    -9,     6,     1,   -22,     0,     5,   -27,   -26,   -29,   -36,     0,    10,   -41,     4,    -9,   -30,   -24,    -4,   -76,   -92,     8,    17,    17,    17,     4,    -6,    16,   -39,   -34,    20,   -44,   -23,    13,   -22,   -86,   -49,    -7,   -31,   -14,    22,   -49,     1,   -11,    -9,   -13,   -35,   -53,  -110,   -52,    14,   -13,     5,    -2,    24,   -11,    24,   -29,    -7,   -81,     0,     7,   -75,  -118,   -53,   -31,   -33,     6,    25,   -70,    -1,     2,     3,   -29,   -50,   -62,   -76,   -27,     3,    45,   -29,   -49,     6,    24,    11,    17,   -38,   -13,    47,   -52,  -115,  -104,   -47,   -50,   -17,    24,    21,   -68,     5,    -4,    -2,    -8,    -6,   -69,   -93,   -50,    -4,    23,     2,    -7,    11,    42,    42,    22,   -10,    20,   -38,   -55,   -68,   -34,   -25,   -31,   -10,   -26,   -56,   -53,     1,     0,    -3,   -34,   -21,   -33,   -49,   -18,   -10,   -38,   -38,    42,   -50,   -57,   -25,   -10,    28,   -19,     1,    16,    31,    30,   -14,   -34,   -17,   -46,   -24,   -26,    -3,    -4,    -1,     8,    -7,   -12,   -36,   -53,    -6,     4,   -29,   -73,   -51,   -42,   -57,   -81,   -76,   -30,   -14,    -4,   -16,   -28,   -30,   -27,    -9,    -3,     4,     7,     4,    -3,     2,    -9,     6,   -18,    -6,    -3,   -26,   -30,   -14,   -15,   -15,    -5,   -19,   -16,     2,    -6,    -8,     1,    -4,    -6,    -6,   -10,     3,    -1,    -6,     7,    -1),
		    19 => (   -4,     4,    -2,    -3,    -1,     2,     0,    -7,     6,     9,    -3,    -5,    -5,    -5,     7,    -1,     9,     6,    -2,    -2,     4,     4,     1,    -5,    -8,     2,   -10,     9,     3,     9,    -7,    -3,     6,    -1,     9,    -6,   -10,    -8,     0,    11,   -12,   -13,    -1,   -24,   -21,   -33,   -12,   -10,     3,   -12,    -1,     1,     9,     7,    -8,    -2,    -8,     8,    10,    -3,     0,    -2,    -5,    -2,    -2,   -11,    -6,    -9,     5,    -3,   -23,   -11,    -1,    -8,   -22,    -5,   -18,     6,    -5,   -10,   -10,    -9,    -5,     7,     1,     5,    -7,    -2,   -10,   -44,    -2,    -6,   -31,    -2,    -6,    -2,    -5,    -1,   -28,   -65,   -32,    14,    66,    24,   -39,   -18,   -22,    -2,    -5,   -14,    -8,     7,    -8,    -3,   -10,   -12,    -1,   -25,   -26,     1,   -12,     3,     9,    -7,   -33,   -45,   -58,   -93,  -102,  -104,   -63,   -76,   -92,   -48,   -46,   -56,   -36,   -51,   -27,    -6,     5,     4,   -18,    -6,    -9,    -6,   -11,    -4,   -42,    -5,   -17,   -38,   -88,  -100,  -129,  -128,  -102,   -86,   -27,   -26,     4,   -11,   -39,   -73,   -54,   -40,   -48,     6,    -5,   -16,   -30,   -31,    20,    -4,   -26,   -29,   -33,   -68,   -53,  -120,  -134,   -72,    -5,   -15,    -6,    41,    34,   -32,   -10,   -20,   -43,   -66,   -36,   -32,   -41,   -46,     4,   -26,   -36,   -16,   -21,   -15,   -30,   -42,   -16,   -94,  -134,   -78,   -26,    20,    21,    57,    50,   -25,    28,    -5,    38,   -30,   -18,    18,   -55,   -40,   -34,   -25,   -41,   -28,   -32,     6,    -9,     0,    62,   -26,    -4,   -43,   -54,   -28,    17,    23,   -21,   -38,    -3,    10,    16,    32,   -57,     3,    47,    34,   -64,   -65,   -34,   -12,    -2,   -31,    33,    30,    36,     8,   -12,   -29,   -75,   -23,    12,    22,    28,     0,   -52,    -2,   -56,   -95,   -31,     1,   -32,   -29,    77,   -30,   -34,   -69,   -12,   -28,     3,   -43,   -75,    34,    39,    11,   -35,   -64,   -28,    18,    22,    41,    13,     9,     5,    -5,   -45,   -53,    -2,    -1,   -17,     6,     1,   -34,   -14,   -56,   -44,   -25,     2,   -18,   -31,     6,    -8,    -6,   -20,    -4,   -25,   -22,    -6,    35,     5,    23,     0,    -5,    13,   -23,    34,     3,   -17,     6,    11,   -24,   -16,   -23,   -46,   -24,     0,     0,    17,     5,    13,   -33,   -41,    -3,    -6,   -24,    17,     8,    12,     2,    84,    55,    37,    -8,     8,   -54,  -100,   -18,   -55,   -16,   -39,   -63,   -53,   -57,     7,   -20,   -18,   -16,   -11,   -25,     5,   -39,     6,   -19,    43,    61,    31,    26,    24,    29,   -16,     2,   -13,  -125,  -116,   -41,   -56,   -15,     5,   -29,   -27,     2,   -13,   -10,   -30,   -17,   -14,   -10,   -14,     8,   -30,   -30,     4,     7,     0,     8,    37,    13,    -5,    -7,     1,  -103,   -71,   -51,   -31,   -20,     6,     0,    -2,    -7,    -6,    -4,   -40,   -10,   -18,   -39,    -5,    -3,     9,   -25,    20,     7,    15,    16,    30,    19,    50,    18,    29,  -139,   -92,   -29,   -42,    19,    20,   -14,    56,     7,     3,    -7,   -29,    -2,    -9,   -84,   -61,   -23,     3,     3,    78,    34,    31,   -35,   -25,    -5,     5,     7,  -117,  -161,   -48,    42,    13,     4,    65,   -39,   -13,     3,     7,   -13,   -21,   -11,   -14,   -73,   -71,   -38,   -48,   -23,    34,    15,   -48,    -1,    37,    -4,   -24,   -31,   -73,   -75,    27,    55,   -45,   -28,    50,   -19,   -43,    -2,    28,    -4,   -25,   -17,   -28,   -30,   -21,   -97,  -104,   -40,    -6,   -22,   -59,    12,    21,    20,   -51,   -37,   -61,   -64,    48,    47,     5,   -13,    -2,     3,   -51,   -29,     0,   -27,   -31,   -15,   -44,   -60,   -49,   -73,  -127,  -102,   -77,   -73,    -9,     6,   -14,    -7,   -53,   -25,   -70,   -14,    24,    64,     8,   -21,   -12,     0,   -19,   -27,    -4,     1,   -23,   -24,   -44,    -7,   -29,   -84,   -62,   -32,   -46,     0,    -1,   -28,    -3,   -59,   -42,   -40,   -52,    37,    12,   -12,   -10,   -14,    38,    22,    -7,    -6,   -10,     0,   -30,   -31,   -39,   -18,    14,   -16,     5,    -6,    -7,   -26,     5,   -11,   -17,     1,   -20,   -60,   -33,    42,    43,    -5,     0,    45,   -67,    41,   -29,    -9,     0,     6,   -23,   -46,    -4,    14,   -30,     5,    18,     4,   -22,     9,   -37,   -52,   -27,   -24,   -26,   -79,   -32,    30,    60,    -2,   -18,    39,    61,    -2,     5,    -5,    -6,    -6,   -16,   -14,   -45,     8,   -15,    43,     8,    12,     7,   -43,   -15,   -30,   -40,   -55,   -31,   -50,   -41,    22,    73,    10,    -2,   -15,    43,   -30,     5,     4,     0,    -1,    -9,   -31,   -21,    17,     4,    31,    -5,     7,   -11,   -37,    -4,   -25,   -31,   -42,   -25,   -18,   -64,   -37,    24,    -6,    -1,     5,   -41,   -26,   -34,    -8,    -9,    -1,    27,   -11,    48,   -14,     2,    36,     3,   -49,   -29,    29,   -18,    17,   -37,   -26,    85,    28,   -37,   -22,    15,    17,   -12,    13,   -52,   -43,   -32,     2,   -10,    -4,     4,    55,    61,     6,    -8,    39,   -10,    25,   -22,    33,    60,    26,    56,    13,   107,    97,     3,   -66,     4,    24,   -18,   -15,     3,   -10,    -1,    -7,   -10,    10,    -2,    -4,    -2,    -6,     6,     4,     2,     4,    34,    68,    58,    58,    74,    44,    26,   -12,   -20,   -13,   -21,   -17,     3,   -10,     5,     1,     3,     7),
		    20 => (    2,    -8,    -4,     0,    -8,    -9,     6,     8,    -2,     7,     2,    -9,    -8,   -13,    -8,   -11,    -4,     6,     5,     9,    -7,    -2,    -8,    -5,    -3,    -1,     9,    -7,   -10,   -10,    -4,     2,     8,    10,    -1,   -17,   -31,   -39,   -43,    11,    10,     3,    -4,    37,    22,    21,   -10,    -3,    -4,    -2,    -9,    -4,    -8,     4,    -8,    -3,     1,     7,    -3,    14,    27,   -10,   -14,    -3,   -21,   -40,   -26,    -5,     5,   -17,   -44,   -34,     4,    -3,     6,    -7,    -3,   -11,   -43,   -36,   -13,   -15,     1,     9,     0,     5,    -7,    17,     3,   -37,   -21,    -8,   -41,   -78,   -26,   -28,   -26,   -62,   -44,   -19,   -18,     6,   -19,   -12,   -52,   -50,   -39,   -62,   -26,   -30,   -44,     2,     5,     0,   -17,   -29,   -26,   -68,   -23,   -16,   -23,   -14,     0,     2,   -40,   -33,   -26,   -13,    23,    33,    24,    23,   -14,   -37,   -32,   -38,     4,   -76,   -32,    10,     2,    -2,   -21,    -9,    13,   -33,   -14,   -40,   -38,    -1,     9,     7,   -13,   -24,     6,    16,    49,    38,    49,    24,   -14,    -9,   -60,   -46,    -5,   -69,   -33,    -1,    -2,    -6,   -25,     0,    -5,     0,    -5,   -17,   -41,   -34,   -11,   -12,   -28,     5,   -10,    26,    34,    33,    40,    21,    41,    19,     0,    -7,   -21,   -43,   -12,    24,    -9,   -31,   -46,   -31,   -23,   -14,     1,     6,   -48,   -23,   -13,    -7,   -12,     3,    18,     2,     8,    24,     6,    17,    23,   -13,    17,     3,     0,    17,   -38,     6,    19,   -60,     8,   -27,   -36,   -18,   -39,   -23,   -42,   -30,   -25,    -3,     1,    -5,   -15,   -29,   -17,     3,    20,    -8,     5,    24,     6,     5,    -7,   -26,   -36,    -8,   -12,   -13,    11,    -5,   -35,   -33,   -59,   -14,   -39,   -29,   -38,    -2,   -13,   -19,   -51,   -41,   -22,   -36,   -49,   -47,   -29,   -29,   -22,   -22,    -9,   -52,   -56,     0,    -8,     7,    29,    -3,   -41,   -53,   -24,    -1,   -36,   -38,   -47,   -56,   -64,   -62,   -30,   -42,   -28,   -19,   -44,   -41,   -74,   -81,   -23,   -17,   -30,   -23,   -42,    -7,    -6,    46,   -47,     6,   -34,   -13,    19,   -22,   -63,   -49,   -48,   -51,   -49,   -31,   -33,   -17,   -30,   -21,   -19,   -11,   -29,   -39,    -7,   -18,   -13,   -21,   -16,    -9,    -4,     8,   -60,    16,   -21,    -3,    -5,   -25,   -22,    -6,   -17,    -3,     5,     7,     7,    -7,    -2,   -10,    12,     4,     4,    -5,     8,   -11,   -15,   -30,   -25,   -13,     1,    15,    -3,    11,    -4,    -9,     5,   -12,   -30,    -2,   -25,   -12,    -8,     5,    -2,   -34,   -18,     0,    33,     4,   -31,     3,     8,    12,    -5,    -5,   -42,   -30,     4,    -3,   -14,   -38,     6,    -1,    -7,     9,    10,    -6,   -54,   -35,   -25,   -19,   -59,   -48,   -36,    -5,    -4,   -37,   -14,    -9,    -3,   -30,   -12,    27,   -46,    -6,     6,     6,   -11,   -54,    18,    15,   -35,    10,    12,   -38,   -54,   -63,   -39,   -92,   -93,   -43,   -31,     0,    -8,    -8,    18,     3,   -25,   -38,    -7,     6,   -57,   -20,     7,    -2,   -30,   -10,    43,    -1,   -33,   -37,    -6,   -57,   -72,   -51,   -74,   -86,   -57,    -2,     1,    23,     8,     1,    25,   -16,   -26,    -5,    18,    17,   -76,    12,    -2,    -5,   -33,    -8,    10,     1,    12,     6,    -6,    -3,   -45,   -42,   -23,   -27,   -16,    25,    12,    28,    -6,    16,    -9,   -21,   -14,    22,    16,     6,   -70,    14,   -14,    -6,   -24,    -7,    18,   -13,     9,    11,    11,    11,   -12,   -34,   -45,   -32,    -2,    38,    28,    21,    -4,   -19,   -21,   -17,     5,    18,     4,    -3,   -41,   -29,     4,     5,     1,    -1,     7,     6,   -10,    30,    18,    17,   -11,   -12,    -2,   -38,     1,    24,     2,   -39,   -60,   -38,    -4,    36,    18,     6,    35,   -66,   -27,   -23,    -6,    16,    17,     9,     4,     8,   -14,   -11,    -7,   -16,    -2,   -16,   -19,   -34,    -6,    -2,   -24,   -50,   -22,    -6,    -4,    -9,    -5,    20,    17,   -19,   -10,    -9,     8,     6,   -14,    -1,    -7,    -4,   -12,    -7,     3,    -1,   -15,   -48,   -31,   -57,   -26,     5,   -21,   -26,     2,     6,     6,   -34,    -7,    21,    20,     1,    15,     5,     0,   -10,   -38,     0,    20,     2,    -4,    -6,    -8,    -4,   -42,   -14,   -22,   -12,    -3,   -40,    -7,   -34,    -1,     0,   -21,    -2,    18,    10,     6,   -10,     1,     4,    -8,    -1,   -35,   -31,   -28,   -17,   -10,   -10,   -44,   -33,   -11,     7,     6,     4,   -23,   -16,   -12,     6,    18,    11,   -12,    18,    22,     8,   -54,   -37,   -23,     3,    -6,     4,    -3,   -24,   -28,    13,   -42,   -16,   -18,   -35,   -75,   -54,   -41,   -38,   -45,   -32,   -22,    13,    -7,    -3,   -15,   -15,   -13,   -22,   -20,    -6,    -5,     6,    -6,     3,     2,   -30,   -52,   -29,   -30,   -26,   -27,   -21,   -33,   -55,   -60,   -72,   -64,   -46,   -51,   -19,   -13,   -61,   -39,   -37,   -41,   -24,     2,    -2,     7,    -4,     2,    -5,    -7,     6,   -38,   -50,   -60,   -29,   -20,   -35,   -38,    -8,   -17,   -36,   -34,   -48,   -42,   -61,   -61,   -68,   -51,   -49,   -39,   -15,     7,     1,     1,     2,     0,    -2,     2,     1,    -2,     4,   -18,   -32,   -29,   -23,    -4,     3,    -4,   -23,     7,   -11,   -15,   -25,   -15,   -23,    -8,   -17,   -25,   -15,    -6,    -3,    10,    -8),
		    21 => (    8,    -3,    -9,     4,    -6,    -8,     3,    -8,    -8,    -9,    -8,    10,     8,     8,     0,     6,    -1,    -8,     6,    -3,     7,    -3,    -4,     1,     9,     1,    -4,    -9,     6,     6,     4,     7,    -7,     2,     7,    -2,     9,    -5,    -8,     8,     1,   -25,    43,    46,    -7,   -36,   -13,   -20,     2,    -6,    -4,     9,     6,     5,    -5,   -10,     4,     2,     2,    -8,   -10,     3,    -6,    -3,    -8,   -49,   -45,   -31,   -79,   -22,   -44,   -42,    -8,   -43,   -22,   -12,   -14,   -56,   -71,   -41,   -31,   -15,     4,    -4,    -2,   -10,    70,    45,    -5,   -38,    -9,    43,    37,    45,    12,   -62,   -42,    58,   -10,   -57,   -44,   -16,   -19,   -35,   -12,   -95,   -63,   -40,   -37,   -13,     8,     7,    -8,    -9,    61,    61,     7,   -20,    -2,    58,    58,    53,    35,   -16,    -5,    20,    -6,     0,   -46,   -48,   -14,     5,   -25,   -64,   -33,   -35,   -34,   -71,   -76,   -57,    -6,     2,    56,     8,    17,    30,    30,    58,    19,    47,    76,    79,    39,    41,     5,   -23,   -26,   -18,   -28,    11,   -22,   -47,   -37,    27,     6,  -120,   -55,   -50,     1,     2,   -26,     4,    25,    11,    38,    71,    18,    23,    87,    38,    14,    31,     7,     1,   -13,     0,    -4,     1,    -7,   -43,   -26,    33,     2,   -53,   -66,   -33,    -4,   -49,   -68,   -58,   -85,    34,    53,    84,   -27,   -31,    38,    12,    37,   -18,    37,    -1,    17,    14,   -39,   -31,    28,   -23,    31,    27,   -16,   -43,  -109,   -69,   -13,   -48,   -63,   -91,   -88,    -8,    55,    60,   -32,   -71,    35,   -36,    13,    46,    31,    24,     9,    33,    44,    15,   -16,    -7,    22,    -8,   -53,   -46,  -116,   -45,     8,   -19,   -64,   -87,   -62,   -29,     0,    42,   -16,   -21,   -40,   -54,   -22,    55,    10,    13,    -6,    42,    57,   -12,     9,    19,     4,   -33,   -45,   -47,   -45,   -66,     3,   -31,   -56,   -82,   -67,   -40,   -38,     1,    28,   -33,   -47,   -55,   -11,    35,     1,    -3,    55,    63,    19,   -13,    -4,   -29,   -38,   -57,   -63,   -40,   -72,     7,    -1,    -4,   -21,   -51,     3,   -14,   -22,    54,    20,     4,   -28,   -40,   -10,    13,     1,     8,    72,   106,    30,    -2,    44,   -51,   -68,   -53,   -67,   -58,   -72,    60,     3,     9,   -86,   -36,    -6,     8,    45,    49,    10,   -26,   -23,    -1,    19,    -2,    22,    46,    45,    63,    40,   -12,     7,   -60,   -63,   -17,   -66,   -22,     6,    55,     3,   -10,   -43,     2,   -26,    24,    44,    21,   -27,   -44,   -19,   -27,    -9,   -19,     2,   -17,     4,    75,   -38,     6,    -1,   -46,   -48,   -95,   -75,    18,    45,     5,     2,    -8,     6,    16,   -34,     9,   -30,   -40,     1,   -29,   -42,    12,    -9,    -9,    38,    -5,   -20,    -6,   -84,   -28,    14,   -17,   -18,   -38,   -68,    26,    80,    -1,     3,    -8,     6,   -23,   -63,   -44,   -21,    -1,   -18,    -6,    13,   -30,    -2,     6,    23,     5,   -23,   -49,   -81,   -58,   -17,    12,   -62,   -64,   -90,   -34,    -3,   -19,    -2,    -3,    11,   -59,   -55,    11,     4,   -40,   -41,    25,     2,   -22,    -2,    31,    27,   -49,   -80,   -79,   -24,   -32,     2,    -3,   -14,    -4,    33,     3,   -26,   -19,     1,    -7,   -13,   -90,   -46,    22,   -10,   -31,   -29,   -49,   -39,    30,    34,    23,    35,   -76,   -63,   -84,   -56,    -5,    12,    30,    52,    56,    45,     0,   -41,   -52,    -9,    -6,   -23,   -88,   -59,   -57,   -96,   -62,   -51,   -34,   -21,     0,   -10,    11,     4,   -23,   -47,   -46,    49,    53,    58,    51,    10,    -6,    22,    35,   -28,    19,     8,    -1,    13,  -104,   -77,   -27,   -15,   -11,    -5,     9,    29,    30,   -24,   -34,    23,   -14,   -18,     2,     6,    35,    97,    49,     6,    41,    57,    46,   -18,     7,    -8,    -2,   -47,   -85,   -16,    -6,    26,   -11,    20,    44,    63,    20,    -4,   -23,   -17,     6,    -2,    26,    63,    57,    90,    33,     4,    -5,    25,    15,    -4,     0,    20,    16,   -70,    -3,   -16,    17,    -6,     7,    -9,    21,    42,   -21,   -50,   -33,   -20,    33,    22,   -12,    75,    69,    85,    70,    -9,   -18,    30,    22,   -28,     2,     7,     7,   -61,   -48,   -21,    18,    -8,   -13,    40,    12,    19,   -18,   -37,     0,   -36,    43,   -11,    20,   122,    81,    50,    71,    16,     1,    27,    42,    -7,     1,    -7,     8,   -21,    -5,   -46,   -13,     6,     5,   -51,   -12,   -24,    -4,    51,    14,    27,    80,    31,    48,    57,    37,    53,    17,    -5,   -44,   -60,   -36,    35,   -10,    -3,    -8,     1,   -11,   -52,   -46,   -50,    -6,   -64,   -71,    15,   -36,     6,     9,     8,    37,    24,    63,    19,    22,     7,    41,    18,   -46,   -40,    19,    10,     3,     3,    -1,    -5,   -26,   -48,   -89,   -99,  -103,   -61,  -150,  -143,  -117,   -13,    -4,   -28,     5,   -54,  -109,  -101,  -125,  -105,   -81,   -33,   -32,   -34,   -29,   -23,     8,     5,     1,    -4,   -23,   -66,  -124,  -115,   -81,  -154,  -151,   -82,   -57,   -76,   -96,    -8,    -9,    18,   -59,   -46,   -16,   -26,   -56,    -5,    -7,     7,     7,    -4,    -4,     7,     6,    -1,    -8,   -14,   -17,   -16,     2,    -5,   -13,   -68,   -39,   -14,   -21,   -32,   -18,    -9,    -5,    12,   -10,   -11,     5,    -5,     0,     0,     6,     9,   -10),
		    22 => (   -1,    -3,    -4,    -2,     1,    -2,     1,    -8,     6,     5,     2,     4,   -18,   -25,    17,    17,    -2,    -6,     0,    -9,    -8,    -1,     2,    -2,     6,     0,     0,    -9,    -9,     1,     5,     6,     6,    -4,   -24,   -25,   -57,   -43,   -25,   -35,   -25,   -53,   -18,     0,     1,   -11,   -25,   -97,   -56,   -30,   -33,   -21,     9,     2,     0,    10,     0,    -5,    -9,   -17,   -32,   -13,    -7,   -32,    22,    43,    51,    47,    39,    27,   -26,   -19,   -11,   -29,   -50,   -60,   -57,   -34,   -23,    -8,     7,    43,     7,    -1,     6,     4,   -20,   -54,   -53,    45,    36,   -29,    -5,    82,    31,    55,    56,    18,    10,   -18,     0,    -7,   -54,   -41,   -20,    35,    -1,   -53,     6,    14,    -7,     3,    -5,    -4,    -2,   -21,    44,   -16,    19,    40,    24,    65,    41,    36,    38,    32,    -3,    11,    20,    31,    14,    -9,    -5,   -38,   -19,   -30,   -22,   -28,   -21,   -23,    -4,     6,    17,    11,    34,    27,    -9,    19,    25,    11,    -4,    -3,     2,     9,    14,    17,    57,    19,    42,   -22,   -16,    -9,    14,   -27,   -28,   -26,   -20,   -21,    -1,     1,    11,     4,    -1,    18,   -16,     6,    39,    13,     8,    -8,    21,     2,    43,    77,    47,     4,    10,     8,   -48,   -32,   -24,   -54,   -93,    -4,   -13,   -16,    -6,     0,    11,   -29,     5,   -11,    34,    33,    27,    32,     0,    10,     2,    19,     6,   -38,     1,    -7,   -13,   -16,   -37,   -49,   -30,   -92,   -35,     7,   -26,    -5,   -31,    25,   -38,   -42,    -7,   -25,   -11,     2,   -16,    -1,    44,    12,   -36,   -18,   -12,   -13,   -13,     6,    25,    24,     6,    -2,   -60,   -58,   -34,   -34,   -11,   -25,     5,     2,    -7,   -50,   -49,   -65,   -56,   -45,   -68,   -69,    -6,    -7,    -5,   -32,   -44,   -45,    -1,   -18,    -7,   -26,     2,   -18,   -21,   -65,   -74,   -53,     9,   -11,     2,    -1,    -5,   -67,   -42,   -15,    10,   -30,   -60,   -73,   -47,   -66,   -43,   -89,   -64,   -63,   -24,    18,    21,    26,    13,   -32,   -92,   -32,   -10,   -16,    -7,   -24,    -7,   -30,   -28,   -54,   -40,   -66,   -68,  -123,  -106,  -110,  -107,  -105,   -91,   -64,   -65,   -87,   -45,    -5,   -32,    27,    -8,   -26,   -20,    24,    25,    -1,   -65,   -19,    -1,   -44,   -48,   -43,   -88,   -80,   -79,  -122,   -96,   -62,   -53,   -81,   -23,    -1,   -17,   -31,   -16,   -21,   -14,    26,   -15,    -9,   -19,   -31,   -80,    16,   -47,   -12,    -5,   -41,   -15,   -33,   -61,   -69,   -37,    -4,   -19,   -39,   -36,    29,    75,    55,    34,   -24,   -14,     3,    37,   -12,    -8,   -46,   -24,     1,    35,    34,    34,    13,    -9,   -45,   -40,    46,    -9,   -19,    16,    23,    28,    49,    67,    76,    84,    15,    44,    19,    23,     4,    23,   -10,     1,   -30,     1,     7,    45,     7,    42,    48,     3,   -20,    -1,    39,    36,    65,    39,     4,    23,    57,    53,    41,    -9,    -6,    20,    29,     3,   -11,    12,   -11,   -34,    14,   -10,   -17,   -10,    44,    42,    71,    -7,     7,    36,     6,    55,    19,    36,    23,     5,    15,    -9,    25,    -1,   -13,    14,    12,    22,    41,    29,    27,    43,    53,    25,     9,   -17,    76,    64,    17,     8,    -2,    29,   -18,    18,    25,    46,    -1,    45,    -1,    34,   -18,     1,   -48,    12,    30,   -15,    35,    27,    11,    -2,   -32,    16,   -18,   -77,    48,   -10,    37,    -5,    -1,   -21,   -62,   -28,    48,    33,    42,    66,    28,     5,   -39,   -49,     0,    11,    15,    28,   -12,   -28,    10,    30,   -31,    41,     5,    22,     2,   -15,    86,    -4,   -27,    -7,   -82,   -19,   -66,     9,    13,    20,     0,    -6,   -58,   -49,   -48,     6,    59,    16,    18,    13,   -31,     0,   -10,    16,   -27,    -3,   -22,    52,    75,    -3,   -39,    35,    -4,    14,     7,   -58,     3,    58,    -7,   -39,   -13,   -26,   -10,   -26,   -28,   -26,   -31,    27,   -18,     4,   -29,   -16,   -38,    45,   -44,    44,    -1,     9,    11,    25,    39,    25,    -9,    -3,    -2,    14,    -3,    33,     1,   -26,   -18,   -21,   -73,   -77,   -40,   -32,     5,   -32,    25,     0,    12,   -48,   -42,   -98,    -5,     8,    10,    23,    70,    34,     8,     9,   -39,   -27,     3,   -18,    -5,   -58,   -33,   -88,  -133,   -25,   -55,     8,     2,   -46,   -38,    21,     9,   -12,   -65,  -105,    -2,     8,    -2,    10,    18,   -16,   -14,   -52,   -42,   -26,   -16,     2,   -24,   -33,   -94,   -58,   -81,   -62,   -65,   -37,  -108,   -67,   -48,     8,   -43,   -37,   -56,  -100,     2,    -5,    -4,   -54,   -24,   -62,   -40,  -118,   -57,   -67,   -86,   -94,   -64,  -108,  -126,  -113,  -109,   -78,   -41,  -127,  -128,   -81,   -34,   -15,   -72,    10,    15,     0,    -9,     7,     8,    -2,    -6,    -2,   -21,   -25,   -48,   -79,   -96,   -56,   -40,   -60,   -69,   -64,   -69,   -92,  -102,   -70,   -88,   -69,   -33,   -25,    -1,    22,    40,    44,    -5,     5,     0,     3,    -4,    -9,   -18,   -16,    -9,   -14,   -20,    -1,    -7,     2,   -14,   -10,   -25,   -35,   -42,   -30,   -13,   -17,     7,   -31,    -5,   -17,    10,    -7,    -8,    -9,    -5,     7,    -2,    -7,     7,    -5,    -9,     0,     4,    -8,   -10,    -4,     0,   -14,     2,     0,    -5,    -6,     4,   -11,   -19,   -10,    -2,    10,     0,     9,     4),
		    23 => (    2,    -3,    -4,    -3,     8,    -7,    -2,     1,    -4,     3,     2,     4,    -4,   -14,     3,    -3,     2,     1,    -7,    -8,     1,    -4,    -4,    10,    -9,     9,     2,     4,     4,    -7,    -1,     5,    -3,     0,    -3,     5,    -4,    -6,   -25,   -24,   -29,   -15,   -26,   -26,   -25,   -38,   -34,   -14,   -12,   -12,   -10,    -9,     9,     8,     1,    -1,     4,    -5,     6,     9,    -8,   -10,     0,   -10,   -51,   -40,     6,     0,   -31,   -25,   -34,   -51,   -80,   -55,   -39,   -45,   -27,   -14,   -19,   -42,    -2,     5,    -5,    -3,     7,     3,   -14,    15,   -15,    35,    54,    80,    38,    20,   -31,    -8,    -3,     7,   -27,    11,    29,   -16,   -97,   -58,   -20,   -64,   -40,   -68,   -20,   -19,     9,     1,    -6,    16,     4,    12,    42,    43,     9,    28,    62,    45,     4,   -13,    10,    14,    13,    -4,     1,     4,   -56,   -79,  -110,   -43,   -52,   -95,   -55,   -13,   -12,    -2,     9,     4,    31,     6,    12,    39,    29,     4,     7,     0,    24,    28,     9,    40,     6,    13,    16,   -31,   -38,   -23,   -93,   -84,  -106,   -89,   -43,   -38,   -21,    -9,     9,    11,    14,    28,    10,    52,    50,    12,    35,    49,    52,   -14,    -3,    23,     3,    17,    13,     9,    23,   -13,   -28,   -90,   -93,   -85,   -24,   -25,   -48,    -8,    -1,     5,     1,    40,    64,    65,    22,    12,   -11,    -7,     1,   -12,   -26,    26,     9,    -2,    36,    20,   -14,   -13,   -73,   -92,   -96,  -104,   -52,    -6,   -45,   -22,   -17,    -6,    12,    22,     4,    51,    46,    35,    -5,   -73,   -29,  -124,   -80,   -23,   -19,    18,    29,     4,     5,    44,   -60,   -68,   -97,  -106,   -74,   -23,   -51,    -2,     9,   -14,   -10,   -19,   -18,   -14,   -21,   -94,  -152,  -135,   -84,   -86,   -23,   -14,    31,    37,    22,    13,     0,   -63,  -132,   -94,   -86,   -50,   -38,   -25,   -47,     5,    -3,   -26,    13,     3,   -57,   -99,  -169,  -180,  -109,   -39,    38,     4,     7,    32,    47,    -5,    -4,    20,   -58,  -105,  -133,  -105,   -23,     4,   -40,   -19,   -29,   -15,     8,   -14,    -8,   -15,  -103,  -111,  -101,   -77,    49,    32,    43,    71,    39,    49,    24,     1,   -62,   -62,   -46,   -77,   -67,   -64,   -43,     4,   -52,   -11,   -27,    -7,     7,   -15,   -23,   -37,   -33,    -6,   -16,    50,    45,    70,    31,    10,     1,    10,    -9,    18,   -47,   -63,   -30,   -45,   -38,   -41,   -22,   -28,   -47,    -6,   -22,   -10,     7,    -7,   -16,   -32,     1,    16,    45,   109,    72,    27,     0,   -30,     1,    -8,    50,     7,    -2,   -56,   -24,   -14,    -2,    -5,   -30,    -8,   -52,   -48,   -35,   -22,     1,     5,     3,   -39,     9,   -21,   -18,    -1,    21,    -9,   -10,   -29,   -31,     3,     1,   -31,   -13,   -21,   -20,    22,     2,    46,     7,    22,    -3,  -102,    -8,   -28,   -12,    24,     1,   -26,    -5,    -5,   -19,   -78,   -31,   -56,   -31,   -55,   -24,    -4,    -1,   -64,     1,    26,    -7,   -11,    -6,    50,    12,    23,    39,   -56,    -8,   -11,    -1,     2,     4,   -32,   -29,   -26,   -58,  -100,   -24,   -60,   -63,  -101,  -145,   -85,   -28,   -43,    -7,    23,     2,    22,    10,    49,    55,    36,    26,  -106,   -87,   -20,    -6,    16,    27,    21,   -32,   -26,   -17,     9,    49,     9,   -19,   -99,  -124,   -91,   -94,   -46,    -3,    17,   -41,   -47,   -10,    14,    23,   -40,   -20,  -108,   -18,   -27,   -11,    18,   -11,    48,    27,    32,    74,   -32,    76,    14,   -17,    -9,   -20,   -43,   -31,   -22,    33,   -26,   -26,    -3,     6,     5,    -5,   -50,   -41,   -54,   -34,   -24,    -9,    -3,   -54,    12,    23,    21,   -19,   -20,    26,   -14,   -19,    27,    50,    42,   -16,   -10,   -46,   -17,   -12,     3,   -21,   -38,     3,   -16,    11,   -33,   -51,   -26,     4,    -5,   -46,    16,   -29,    12,    22,   -11,    16,    23,     1,   -32,   -27,   -28,     4,   -23,     4,    -4,     8,   -35,     6,   -55,   -43,   -16,    19,   -15,   -43,   -10,   -11,    -1,    15,     3,     2,     3,    10,    16,    14,    27,     3,    19,    36,     5,   -35,   -35,     7,   -28,    -8,     5,   -15,   -41,   -13,   -13,   -30,   -11,   -28,     0,    -2,    -1,    -1,    31,    61,    17,    44,    11,    -1,    17,    14,     9,    -4,     1,    -3,    -1,   -39,   -15,   -14,     2,   -17,    -7,    14,    20,    16,   -40,    -2,    -7,    -3,     5,    20,    81,    82,    17,    11,    38,    12,     9,    10,     2,   -26,    29,   -14,     4,   -11,   -21,    19,     2,    11,     5,   -30,     7,    34,     4,    -9,     3,    -1,    -3,   -21,    15,   -10,    -6,   -58,    29,   -22,   -26,   -21,    19,     0,    -5,    -5,   -23,   -25,   -22,    -8,   -29,   -27,   -48,   -53,   -44,   -28,   -12,     2,    -6,    -6,    -2,     8,   -15,   -12,   -20,    34,    49,    45,   -11,   -19,   -42,   -93,   -38,   -48,   -29,    21,     5,    -3,    41,   -11,   -52,   -74,   -50,     4,   -14,    -7,    -9,    -1,    -7,     8,   -19,   -24,   -29,   -22,    -4,   -27,   -41,   -26,   -33,   -54,   -59,   -72,    -1,    14,   -15,   -10,     6,   -24,   -35,   -52,    -1,     0,    -4,     3,    -2,     2,     4,    -6,     6,    -4,    -7,    -8,    -2,     1,   -11,   -18,   -56,   -35,   -67,    -2,   -15,    -6,     6,    -4,     7,   -14,    -9,   -20,    -9,     9,   -10,     8,     1),
		    24 => (    1,    -3,   -10,     5,     7,    -5,     9,    -4,    -6,     0,    -7,    -4,   -29,   -27,   -14,   -17,    -5,     8,     3,     3,     5,   -10,     2,     7,     6,   -10,    -1,    -2,     3,    -2,     2,     9,     3,    -6,   -28,   -32,   -17,   -43,   -56,   -25,   -84,   -13,    28,   -29,   -55,   -34,   -43,   -16,   -31,   -10,   -15,   -34,    -5,     0,    -3,    -5,    -9,     0,   -11,   -90,   -99,   -22,   -33,   -68,   -72,   -48,   -65,   -89,   -87,   -30,   -10,   -64,   -54,   -51,   -31,   -68,   -30,   -13,    -9,     0,     1,   -11,     6,    -1,     9,    -3,    -9,   -76,   -74,     1,   -35,   -72,   -61,   -88,    -9,   -48,  -100,   -60,     1,     1,    36,    25,    26,     1,   -25,    -3,    29,    23,    40,   -25,     3,    -6,    -8,     8,    -3,   -20,    17,   -59,    -8,   -25,   -21,    -4,   -12,    10,   -23,    23,   -39,    -6,    18,    -6,   -34,   -48,    36,    31,    75,    86,    47,     8,   -39,   -11,    -8,     0,   -18,    23,   -33,    -9,   -27,   -43,   -36,   -25,     3,    26,    12,   -21,   -31,   -31,   -66,   -75,   -38,   -16,    23,    -3,    -4,    13,     6,    -2,     5,     7,    -8,    -7,     6,   -15,   -20,    19,   -34,   -53,   -17,    23,    17,   -31,   -40,   -11,   -28,   -23,  -146,  -181,   -78,    -5,    47,    12,    31,    12,   -44,   -17,     5,   -39,    -3,    -8,    -7,   -28,   -12,   -20,   -29,   -24,    12,     6,     3,    -5,     8,    12,   -12,   -93,  -168,  -149,   -43,    28,    22,    42,    80,    57,   -31,   -58,    45,   -34,   -17,   -28,    26,   -20,   -46,   -41,   -28,   -14,   -16,   -48,    -8,   -27,   -15,    27,   -30,   -83,  -147,  -114,   -21,    20,     4,     8,    45,    40,   -24,    -9,    25,   -44,    -2,   -17,    29,   -29,   -29,   -20,   -16,   -28,     5,     8,   -12,   -27,    15,    13,   -57,  -128,  -154,   -91,   -17,    63,    31,    -4,    42,    23,     5,    -5,   -36,   -13,     5,    -2,    23,    38,   -22,   -25,   -39,   -21,    11,     1,    -9,    18,    21,    -6,  -108,  -142,   -97,   -50,    52,    50,    10,   -10,     1,    12,     9,   -13,   -14,   -27,    -4,   -20,   -14,    11,   -23,   -25,   -12,   -24,    -2,   -20,    18,    14,    -7,   -18,   -45,   -90,   -61,   -11,    13,    56,   -20,    -2,     0,    14,   -12,   -28,   -28,   -48,     0,     3,    24,   -30,   -23,   -41,   -22,     8,     7,   -10,    -2,    -4,    19,   -28,   -98,   -53,   -61,   -12,    52,    26,     4,   -26,    -5,    10,   -37,   -44,   -30,   -52,    -8,   -18,   -15,   -31,   -14,    -2,    -8,    -8,    22,    -8,    -5,   -24,     1,   -41,   -46,   -44,   -42,     0,   -22,   -18,    -9,    21,    21,    -7,   -75,   -10,   -31,     1,     0,    -2,   -42,    61,    12,    79,   -12,    16,   -44,    21,     5,     2,   -30,   -47,   -27,   -36,   -26,     1,   -41,    13,    -4,   -16,    -7,   -23,   -28,   -57,    -3,    -4,    -1,    10,   102,    54,    16,    27,   -27,    -7,    -6,    52,    42,     5,   -31,   -15,   -43,   -42,   -41,    22,    -7,    -3,    -7,   -43,    26,   -18,   -98,   -57,   -40,   -13,     7,    10,    33,     2,   -79,   -14,    35,    45,    78,    47,    90,    -5,   -25,    -1,   -32,    -9,     6,    -6,     2,     0,    11,     0,    31,   -59,   -56,   -58,   -26,   -28,   -10,    -5,    -6,   -50,   -51,   -24,    17,    52,    71,    38,    58,    28,   -33,    -5,     9,     1,    -9,    10,    63,    42,    21,    38,    24,    -3,   -66,   -43,    23,   -29,   -10,     4,    -3,  -101,    13,     8,    -8,    12,    12,     6,     5,     7,    36,    -6,    17,    31,    19,    33,    42,    30,    16,    24,    16,   -36,   -73,   -42,     1,    -4,     1,     1,   -10,   -65,   -15,    33,    41,     8,    -7,     7,   -16,   -24,   -38,   -13,     2,    30,     3,     0,    17,    43,    -5,   -45,   -25,   -38,    -7,   -73,   -23,    -5,    -5,    -7,     5,   -74,   -61,   -16,   -38,   -29,   -41,   -67,   -73,   -65,   -15,   -29,    15,    -8,   -30,   -14,   -39,    45,    17,   -23,     9,     9,    13,   -56,   -26,    -1,     1,     0,   -16,   -60,   -18,   -26,   -30,   -17,   -60,  -113,  -109,   -41,   -31,   -18,     0,   -24,    -5,    -7,    -5,    26,    -8,   -23,    33,    29,    -6,   -64,   -31,    -6,    -9,     2,    -9,   -51,   -58,   -35,   -47,   -69,   -88,   -79,   -86,    39,    -6,   -28,   -36,   -12,    -3,   -28,   -20,     6,   -35,    28,    35,    46,   -27,     6,   -15,    -7,    -6,    -9,    -5,   -15,   -43,   -24,   -48,   -61,   -24,   -23,     0,    31,    14,   -13,    -6,   -35,    14,   -11,    -9,   -13,   -56,    32,     5,    12,   -41,   -24,   -14,    -5,     3,     4,    -2,   -11,   -23,     8,    -6,   -44,   -12,    -1,    -5,   -12,    -9,     2,   -31,    -5,    27,    21,   -49,   -26,   -64,    -3,    41,    27,   -48,   -31,   -12,     3,    -9,     5,   -24,     9,   -11,    -9,   -16,    -1,     5,   -13,     3,   -26,     2,     7,   -67,    -4,   -24,   -45,    10,   -11,   -53,   -61,   -14,    10,   -29,    -5,    -8,    -6,     6,    -3,     2,    -9,    -3,   -11,   -11,    -1,    -7,    21,    25,    17,    28,    12,  -105,   -70,   -28,   -36,   -51,   -12,   -64,   -76,   -66,   -26,   -17,    -2,     3,     7,     8,     7,    -8,    -9,    -3,     2,   -20,   -27,   -34,   -12,   -28,   -24,   -12,     4,    -2,    -7,   -40,   -52,   -12,   -27,   -20,   -43,   -37,     0,     0,    -9,    -9,     1),
		    25 => (   -8,     6,     5,    -8,     3,    -1,     4,     8,     0,    -8,    -4,     3,     2,   -10,    -7,     2,    -1,    10,    -3,     3,     9,    -8,    -6,    -4,     8,    -9,    -4,     3,     3,    -7,    10,     9,    -5,     9,    -3,    -2,     1,     7,   -11,   -20,    -9,   -16,    -7,   -21,   -25,   -34,   -29,   -15,     0,    -1,     0,    -3,     6,     2,    10,     3,    -8,     4,     2,    -9,     3,    -1,     3,     0,   -16,     2,   -23,   -25,   -19,   -11,   -30,    -5,   -25,    43,    33,   -35,    13,    -5,   -12,   -10,   -13,   -28,    -5,     5,     1,    -7,    -8,    12,    22,   -30,   -16,   -22,   -11,   -11,   -14,   -30,   -40,   -65,   -19,    14,     9,    29,    35,   -25,    17,    36,    14,   -36,   -30,   -14,    32,     4,     6,    -4,   -14,    18,   -12,     4,    -7,    -7,   -11,    -7,   -30,   -91,   -66,   -71,    -3,    31,   -27,    19,    32,    -1,   -21,    -4,   -23,    19,    20,    17,     5,   -56,     0,     2,   -22,     5,   -10,    -5,   -14,   -12,   -14,   -33,   -71,   -84,   -40,   -32,   -27,   -14,     5,   -12,   -20,    -2,     2,   -38,   -15,    38,    17,    58,   -14,   -30,     2,     6,     7,   -10,   -15,   -30,     4,   -24,   -16,   -31,   -41,  -116,   -15,   -18,    40,     4,    -6,   -30,     1,    35,    15,   -10,    45,    40,    49,    47,    -4,    -2,    -2,    -2,     3,   -20,   -17,   -13,    11,     0,   -25,   -89,   -16,   -85,   -36,   -10,    -7,    12,    19,     7,   -22,     0,   -11,    19,    41,    44,    31,    71,    13,     7,   -10,   -30,   -36,   -15,    -6,   -10,    22,   -26,   -34,   -25,    -8,     3,    45,    -7,   -12,    -6,   -26,   -23,    11,     8,   -23,    22,    43,    66,    59,    65,     2,    33,    -7,    -1,   -39,   -24,    -6,    16,   -26,   -25,    -1,    -8,    24,   -14,    21,   -34,     1,    -8,   -25,     7,   -11,   -18,    -8,    -6,    42,    64,   107,    64,     0,    47,     0,   -15,    -6,    -2,   -17,    -3,     2,    -1,   -17,   -56,    28,   -20,    17,    22,    50,    -1,   -18,   -29,    23,    25,    30,   -34,    12,    17,    63,    43,    37,    40,    -8,     3,   -13,    -7,    -4,    -2,    13,    -6,    -3,   -13,    28,    -6,    -3,    -9,   -27,   -27,   -71,   -60,   -53,    12,   -70,   -33,    -8,     9,   -11,    15,    54,    15,     7,     5,     4,    -8,   -22,    -6,    13,     9,    29,     1,    12,   -13,     9,    33,   -22,   -70,  -129,  -141,  -129,  -139,  -128,  -129,   -84,   -39,   -43,    -2,    32,   -52,    -6,   -13,     5,     0,   -26,    -6,    30,    23,   -12,     8,    18,   -27,    14,     6,     7,   -54,   -81,  -102,  -135,  -107,  -117,  -115,  -115,   -68,     4,     0,    47,   -27,    14,     2,   -18,     2,   -14,   -21,    -8,     4,    -7,   -20,    26,   -29,    -6,    -2,   -18,   -21,   -49,  -105,  -128,  -103,   -89,   -76,   -59,   -50,     9,     9,     0,   -27,     4,   -15,   -23,     0,   -19,   -55,   -47,   -51,    -5,   -11,   -11,   -10,    35,   -21,    10,    14,    -7,    -2,   -57,   -83,   -99,   -73,   -58,   -31,   -17,     0,    -7,   -13,    10,   -14,   -22,    29,   -19,   -43,   -74,   -83,   -34,   -37,   -22,   -12,    -3,     5,    19,     0,    16,     7,   -46,   -72,  -103,   -70,   -51,   -46,   -14,   -17,   -28,   -11,     7,    -6,   -53,    62,    18,   -44,   -76,   -79,   -35,   -56,   -66,   -12,    25,    -6,     8,    -6,    26,    45,   -47,   -59,   -82,   -52,   -37,   -54,   -45,   -18,   -34,   -32,    -1,   -10,     3,    71,    52,    30,    -1,    -9,   -54,   -63,   -50,   -48,   -27,    10,   -12,   -17,   -24,   -23,   -44,   -28,   -84,   -41,   -28,   -35,   -13,   -14,   -36,   -12,     2,    -5,    13,     7,    49,    37,    49,    61,    -9,   -44,     3,   -35,   -39,    24,   -34,     1,    -3,    39,   -44,   -30,   -38,   -21,   -23,   -32,   -11,   -52,   -26,   -22,    -9,    -6,     3,     8,   -15,    35,    37,    68,    32,     6,    -6,     7,    12,    27,     5,    12,    42,    -3,   -17,   -51,   -34,   -20,   -12,    -2,    -6,     0,   -15,    -4,     3,    -6,    -2,   -13,   -33,   -29,   -38,    32,    38,    17,    -6,    21,    21,     9,    38,    21,    12,   -18,    -8,   -28,   -31,    -9,   -11,   -14,     0,     2,   -11,     1,     0,     8,   -23,    31,    -6,   -35,     4,    18,     3,    -2,     3,    47,    29,    -6,     3,    10,   -33,     3,    -6,   -29,   -35,     1,     3,    -6,     4,   -18,    -5,    -8,    -4,    -5,    28,    22,    26,   -14,    -2,    58,    52,    49,    21,    53,    31,    11,    21,     0,    -3,    34,     3,    -5,   -16,    -1,    -3,    -6,     9,   -12,   -38,     0,    -3,     1,   -18,   -10,    -1,   -34,    11,    38,     6,    65,    44,    40,    37,    18,     4,   -22,   -30,    18,   -20,     9,    -3,    -6,     2,    -5,    -5,   -55,   -19,     9,    -6,     4,     5,    -2,   -45,   -41,    -7,   -35,   -23,    30,    -8,   -20,   -21,    -3,   -54,   -46,   -31,   -22,    36,    17,    -1,   -17,   -10,    -6,     6,     1,    -1,    -1,    -7,    -5,     0,    -6,   -22,   -21,   -71,   -70,   -29,   -12,    20,    35,    45,    20,   -58,   -71,   -18,    -1,   -20,     1,     5,     7,    10,   -26,     6,    -3,     0,     0,     5,     8,     4,    -1,   -14,     2,   -15,    -1,    -9,    -5,    -2,    10,     8,    -5,   -13,    -1,     2,     6,    -3,   -10,     3,    -8,   -35,    -1,     1,    -9,    -9,     0),
		    26 => (    3,    -2,     9,    -3,    -7,    -7,     3,     9,    -4,    -3,     3,    -8,    38,    29,    -4,     3,    -3,    -6,     3,     3,     2,    -3,     5,     1,     6,    -3,     8,    -4,    -9,    10,    -3,     2,    -7,    -4,    27,    40,    44,    28,    86,    77,    14,    36,   -37,     7,   -16,     4,    29,    35,   104,    37,    20,    41,     9,    -1,     4,    -9,    -8,    -1,    15,    26,    54,    73,    32,    49,    94,    76,    40,    44,   -73,   -46,    -2,    -5,    -4,    46,    26,    -3,    31,    31,    59,    34,     7,   -41,    -7,     4,     8,     3,   -84,   -16,    -4,    71,    62,    20,     9,     7,   -11,   -53,   -73,   -13,    33,    20,   -12,    31,    30,    23,    -4,   -24,     7,    73,    36,   -57,   -44,     5,    -2,     5,   -76,    -2,    -1,    57,    -6,   -16,    41,    54,   -19,   -42,  -119,   -31,     3,   -35,    17,   -11,   -41,     3,   -18,    31,    36,    68,    -7,   -79,    44,    69,    10,    -6,   -63,   -50,    22,   -27,   -73,    40,    26,    10,   -48,  -104,   -40,   -25,     2,     0,   -60,   -10,   -58,   -34,    -4,     2,    12,    46,     9,   -39,    94,    62,     0,    -8,    26,   -16,    13,   -25,   -48,    26,   -19,   -71,   -44,   -51,     7,   -55,   -52,    -5,   -22,   -16,    -8,    10,   -16,   -34,    39,     2,    21,   -31,    26,    37,     0,     3,     2,   -31,    17,   -10,   -26,   -12,   -33,   -53,   -53,    -9,   -12,   -25,   -18,   -29,    -9,   -16,   -43,   -13,   -18,    -7,    -1,     8,     9,    -4,    17,    30,    -7,    10,   -39,   -33,    22,   -33,   -49,   -46,   -34,   -63,    -7,   -18,   -33,   -23,   -44,   -45,   -30,   -41,   -84,    -2,   -73,    -3,   -18,   -16,    25,  -100,   -19,   -69,     8,     1,   -47,    16,    11,   -76,   -21,   -55,   -50,     2,    -7,    10,   -34,   -27,   -12,   -68,  -105,   -94,  -100,   -56,   -59,   -56,  -148,   -50,    12,    -5,   -23,   -72,    -6,    -6,   -60,   -50,   -30,   -58,   -80,   -82,   -50,    20,   -32,   -13,     8,    -4,   -36,   -44,   -75,   -58,   -36,   -27,   -29,   -28,   -46,    36,    44,    69,   -40,   -88,     6,    -5,     4,   -36,   -23,   -26,   -44,    -5,   -10,    11,    30,    21,    11,    49,    15,   -16,    -9,   -25,   -55,   -70,    15,   -39,   -34,    11,    11,   -18,   -49,   -23,     5,    -1,    -9,   -38,   -30,   -59,    -1,    24,    47,    65,    61,    21,     6,    12,    -6,   -13,    17,   -11,   -44,   -98,   -74,   -18,    34,    70,    48,    -6,   -82,   -16,     8,     2,   -18,   -31,   -33,    -5,    61,    30,    11,    44,    62,    16,     6,   -23,   -14,    -1,    -3,     5,   -37,   -30,   -50,   -28,    19,    70,    45,    23,   -25,     9,     0,     8,   -10,   -64,   -51,    42,    20,    23,    48,    67,    19,    41,    -4,   -38,    -6,    -6,    17,   -14,   -17,   -12,   -14,    28,    54,    43,    15,    21,   -62,   -43,     4,     3,   -25,   -72,   -63,    51,    54,    61,    88,    82,    50,    38,    39,    10,   -19,   -35,   -10,     0,    -7,    17,     9,   -16,    53,    46,   -53,   -26,   -83,   -42,     3,    -3,    -1,   -60,   -10,    38,    32,    67,   106,    95,    69,    63,    63,     5,    11,    -6,    23,   -13,   -19,    49,    28,    12,    40,    54,   -31,   -54,   -76,   -45,    -7,   -10,    -4,   -57,   -59,    24,    25,    45,    36,    35,    77,    26,    64,    81,     7,    -4,   -11,   -23,   -12,    21,    18,    39,    -5,   -10,   -19,   -59,   -90,   -71,     9,    -3,    -9,    -6,   -34,   -24,    -8,    35,   -21,    23,    21,     2,    56,    80,    25,   -47,     3,    -1,   -28,   -46,    -4,   -12,   -21,   -34,   -95,   -67,   -47,   -48,     5,    -3,   -50,     4,     0,   -69,   -47,   -14,   -41,     1,   -13,    30,    26,    11,    -2,   -14,   -20,    26,   -27,   -21,   -18,    -5,    -9,    -7,   -44,    13,   -36,   -59,     8,   -14,    -4,   -68,    15,   -52,   -45,   -38,   -31,     9,   -12,    -5,   -13,   -39,    32,    -7,   -44,   -29,    -4,   -21,   -10,   -20,    44,     1,    35,    67,   -14,     2,    -8,     1,   -23,   -32,   -31,   -25,   -44,   -14,    -9,    14,     8,   -42,    53,    54,     5,   -33,    -8,     1,     8,    32,    -9,    -3,    41,    47,    44,    19,    -9,   -19,     5,    -6,     0,   -24,   -33,   -88,   -89,   -56,    25,   -32,     4,   -26,    42,    52,    16,    24,    39,     7,     9,    19,   -15,    33,   -15,    -1,   -30,   -72,    -9,   -13,    10,     1,     8,   -10,   -41,   -70,   -83,   -62,   -36,   -20,   -23,     3,   -27,     6,    -8,    17,   -28,     1,    40,    55,     2,   -47,   -75,   -60,   -55,   -55,   -83,     4,    10,     4,    -2,    -2,   -24,   -21,   -11,   -55,   -57,   -82,   -91,   -64,   -23,   -41,     6,    26,    36,    40,    11,   -98,   -41,   -97,   -59,   -46,   -29,   -36,     4,     0,     7,    -3,     0,    -8,     1,   -16,   -14,   -50,   -25,   -31,   -46,    -2,    47,    -2,   -38,   -16,   -44,   -38,   -14,   -37,   -71,   -23,   -28,   -25,   -20,    -3,    -2,    -6,     7,     0,     5,    -7,    -1,   -17,   -24,   -11,    -3,   -12,   -31,   -25,    -5,    -9,     1,   -12,    -6,     3,    -4,    -9,   -13,   -17,   -11,    -6,   -11,     5,    -2,     8,    -9,    -1,    -7,     9,    -8,    -8,     9,     3,    -5,    -3,     1,     2,     8,    -2,    -8,    -3,    -1,   -11,     1,   -10,    -2,   -14,    -3,    -5,    -2,   -10,     1,    -1),
		    27 => (   10,     2,     9,     2,     7,     6,    -4,     9,     4,    -4,    -6,     7,    -5,    -7,    -3,    -3,     2,    -9,    -8,     0,    -8,     7,     2,     0,     1,     2,    -6,    -1,    -9,     5,    -1,    -9,    -8,    -9,    -4,     9,     9,    -4,    -2,   -44,   -31,   -39,    -3,    -8,   -14,   -10,     5,    -5,    -3,    -9,   -10,    -9,    -2,    -5,    -6,    -8,    -8,     5,    10,   -13,   -15,     1,     0,   -14,   -10,    -6,   -12,   -26,   -45,   -28,    -9,    -9,    -3,     7,    -4,   -11,     0,    -4,   -14,    -1,     5,    -7,    -1,     6,     9,   -10,    -1,   -20,   -21,   -16,   -15,   -25,   -39,   -37,   -27,   -51,   -37,   -18,    -8,   -14,   -27,   -23,    -3,   -26,     0,   -34,   -26,   -16,    -8,     2,     9,     5,    -8,     7,     1,    -3,   -53,     1,   -13,   -50,   -45,   -64,   -87,   -81,   -73,   -86,   -63,   -69,   -52,   -24,   -20,   -12,    -2,   -37,   -56,   -42,   -34,   -26,   -15,     5,    -3,     8,     4,   -31,    10,    14,   -13,   -50,    39,    32,   -43,   -34,   -58,   -51,   -44,   -59,   -78,  -161,  -194,  -128,   -89,   -33,    -3,   -88,   -67,   -65,   -32,    -1,    -5,     4,    10,    86,    67,    54,   -24,   -51,    54,    -6,   -32,    -5,    27,    34,     3,   -60,   -11,     8,    34,    -7,    22,    78,    -2,  -111,   -83,   -78,   -55,    -3,    -6,    63,     0,    66,    64,   -20,     1,     4,     7,    28,    49,    42,    29,     1,    -9,   -11,    15,    17,     6,    46,    32,    42,    63,    71,    -4,   -32,   -63,   -31,   -47,    77,    18,    50,    26,   -42,   -36,    13,    28,     7,     5,    19,    13,    15,    -4,    15,    21,    -9,    15,    19,    14,    32,    24,    13,    24,   -44,   -85,   -20,    -5,    48,   -24,     9,    28,    22,    -2,    36,    38,    50,    47,    31,    50,     1,   -13,    -6,   -15,     9,    -3,    40,    15,    70,    15,    -2,    -8,   -17,   -79,     0,     2,    28,    -3,   -32,    52,    41,     7,    19,    24,    23,     9,    55,     9,   -18,   -68,   -36,     5,    55,    -9,    29,    38,    20,    15,   -20,   -40,   -49,   -50,    11,     3,   -23,    61,   -10,    50,    16,    18,    39,     3,     8,    66,    83,   -11,  -101,  -152,   -26,    17,    28,    -9,    -6,    37,   -17,   -10,   -18,    12,   -72,   -18,     6,     0,    33,     8,     6,     5,    41,   -32,    25,     6,     0,    40,   -11,   -91,  -229,  -150,   -15,    20,    -5,    15,   -67,    -4,    11,    -8,   -83,    -4,   -27,   -21,    10,    -6,    39,     3,    -8,   -34,   -11,    14,    30,    38,    31,    24,    -2,  -141,  -243,   -90,   -29,     9,     0,   -47,   -66,     3,     9,   -65,   -81,   -29,   -20,   -26,   -14,     0,     8,    35,     7,    -9,   -23,    42,    23,    18,    19,    51,   -74,  -204,  -207,    -3,    -7,    11,   -12,   -55,    -9,     0,   -32,   -32,     5,    32,   -21,   -13,    -4,     0,    -8,    33,    -9,   -31,    10,    -2,    39,    -2,   -12,     1,  -133,  -226,   -52,   -27,   -45,    -8,   -20,   -13,    -7,    16,   -15,    -7,    13,    34,    -6,     1,    -8,    10,     3,    30,   -30,   -38,     1,   -22,    -2,   -10,   -53,   -62,  -131,   -76,   -26,   -36,   -24,   -37,   -17,   -28,   -17,     8,    -6,   -21,   -62,   -70,   -32,    -3,   -21,     6,     1,    -1,   -25,   -34,   -24,   -88,   -47,   -36,   -36,   -26,   -19,   -70,   -57,   -33,   -21,     6,     3,    34,    14,    -5,    11,    -1,   -65,   -84,   -38,     0,   -42,    10,    -7,    51,   -56,   -65,   -12,   -37,   -41,   -44,    -8,   -12,   -50,   -61,   -37,    -8,   -40,     6,    20,    22,    15,    -3,   -55,   -27,   -44,   -97,   -75,     0,   -26,    10,    24,     4,   -64,    10,    32,   -12,   -75,    38,    38,   -23,    -2,   -26,   -16,    14,   -17,   -13,   -34,   -34,   -10,    -5,   -43,    13,   -44,   -47,   -26,    -7,    -9,     2,    49,   -12,   -17,   -26,   -71,   -57,   -16,    -4,    10,     6,   -17,    46,   -22,    -7,    -9,   -48,   -33,   -40,    -3,   -41,  -102,   -76,   -75,   -61,    -6,   -22,     9,    -2,     9,    -5,   -37,   -67,   -56,   -52,   -79,   -18,   -33,     9,    43,    16,    -4,     5,   -17,   -16,   -42,   -16,     6,    -9,    21,    17,   -36,     4,    -5,   -27,    -2,     3,     3,   -12,   -32,   -46,    15,   -52,   -36,   -12,     6,    -4,   -21,   -20,    10,   -12,     9,   -26,   -22,    15,    15,   -38,   -16,   -25,   -36,   -17,     4,   -81,     4,     1,     5,   -15,   -39,    12,    48,    20,     8,   -32,    20,    35,   -25,   -55,     8,   -26,     2,     5,     5,   -25,    -6,   -42,     4,   -51,   -31,   -15,    -6,   -44,    -5,     1,    -6,    26,    53,   111,    66,    -7,   -20,     3,   -30,    41,   -22,   -16,   -61,   -77,    12,   -17,   -11,   -24,    -7,   -36,     8,   -27,   -16,    -3,   -20,    -2,     4,     7,     8,   -51,    38,     9,   -61,   -45,    -7,    15,    -1,   -52,   -23,    42,    -7,    35,    15,    -2,    10,     4,   -16,    11,    68,    34,   -36,   -10,     2,     6,     0,    -1,     1,   -10,   -31,   -51,   -70,   -29,    42,    56,   -11,   -54,   -45,   -35,    16,    -1,    33,    17,   -22,     0,    47,    33,    -9,    -4,   -12,   -18,   -11,    -3,   -10,     0,    -8,     4,    -1,    43,    49,    17,     3,    27,    27,    18,     4,     7,    50,    49,   -10,     0,    49,    14,    39,    30,    11,     9,    60,   -10,    -5,    -8,     3),
		    28 => (   -1,    -8,    -6,    -2,     1,    10,    -9,    -3,     1,    -5,     9,    -7,    -9,    -9,     0,    -6,     8,     5,    -7,    -1,    -4,     9,     0,     1,     0,     1,    -2,     5,     3,    -9,     3,     8,     1,    10,     3,     0,     7,    -9,    -9,   -35,   -36,   -42,   -41,   -77,   -61,   -78,   -11,   -17,    -5,    14,     4,     4,     6,    -1,     3,   -10,     8,     0,    -1,    -8,   -12,    -5,   -19,    -2,   -29,   -68,  -110,  -101,   -50,   -38,   -16,   -91,   -91,   -81,   -35,   -64,   -37,   -44,   -54,   -43,   -15,   -17,     7,     1,     6,    -9,   -35,   -26,   -17,   -67,  -111,  -138,  -162,  -177,  -111,   -99,   -24,    50,   -28,    -4,   -27,   -55,  -112,  -108,   -27,    18,    39,    48,    32,    -2,   -22,    -3,    -3,   -38,   -22,   -67,   -83,  -133,   -62,   -59,   -19,   -26,    -4,   -46,   -44,    24,    22,    -1,   -12,   -29,   -41,    19,    35,   -41,   -31,   -33,    26,   -41,    48,    -7,     5,    -4,   -58,   -51,   -43,  -111,     1,    -7,    12,    -3,   -38,    -6,   -18,    -1,    26,   -29,   -13,    -7,   -60,   -11,   -10,    43,    30,   -16,    73,    61,   -51,    12,    -2,    -2,   -19,   -91,   -34,   -45,    30,     3,    -1,    -6,   -10,    17,    15,   -29,   -28,   -12,    12,    -8,    29,   -26,    20,    34,    38,    54,    18,   -40,   -44,     4,    -8,   -33,   -21,   -80,     5,    19,    -7,    31,     7,    -9,    25,    -5,   -17,   -28,   -49,     5,     5,     0,     9,     1,   -42,    36,    66,    22,   -20,   -34,   -63,    10,   -32,   -42,   -70,    -5,    -9,   -21,    18,    22,    -7,    35,    -9,   -37,   -23,    13,   -26,   -70,   -46,    13,    31,     3,     1,    -7,    44,    27,    49,   -40,    33,    30,    -7,   -31,   -76,    -7,   -60,   -12,   -12,   -23,    34,    -9,   -22,   -19,   -30,   -14,   -44,   -59,   -24,    21,   -51,    39,   -19,   -23,   -12,    41,    55,    -3,    25,   -31,    -9,   -11,  -103,   -92,    18,   -11,   -17,    27,    -4,    32,   -23,    -8,   -12,   -32,    68,    13,   -19,   -28,   -15,    14,     9,     1,     8,    82,    45,   -48,    17,   -13,     1,    -8,   -63,    66,    21,    18,   -13,    -6,    22,    -5,     8,    -3,    17,    34,    65,    72,     7,    -5,   -14,   -12,    21,    21,    -7,    26,   101,    99,    52,   -42,     2,    -3,   -43,    75,    44,    33,   -24,     5,    -3,   -44,   -45,    43,    70,    72,    39,    45,    23,    57,   -19,    60,    17,     0,   -62,   -12,    26,    69,    32,   -45,    -2,     2,   -27,    88,     5,    10,   -15,    21,   -30,     5,    13,    66,    43,    67,    58,    54,    35,    30,    36,    50,   -18,   -67,     9,   -31,   -61,    -7,   -23,     4,    -6,    -7,   -12,    65,    20,    11,    19,   -30,   -49,    -8,    81,    49,    36,    67,    33,     4,    33,    27,    30,    21,   -62,   -81,   -46,   -33,   -54,    64,   -63,     1,    -5,    -3,   -24,     0,   -87,   -60,   -22,    20,    10,    51,    57,    42,    36,    64,    43,    21,    40,    29,    -7,   -33,   -44,   -65,    11,    18,   -72,    72,  -143,   -48,   -10,    -9,   -13,   -11,   -19,   -15,    15,     9,    20,    26,    80,    22,    71,    -6,    17,    12,    66,   -42,   -28,     5,   -54,   -28,   -12,    64,   -79,    32,  -118,   -54,    -6,    -7,   -14,   -52,    52,    22,    82,   -14,   -31,    34,    58,    77,    69,    76,    56,     0,    71,     2,   -49,   -22,   -36,   -22,    14,    99,    32,   -59,   -29,   -72,    -9,   -12,   -22,   -63,    59,    -6,   -18,    11,   -14,     9,    35,    50,    99,   118,    54,    43,   -13,   -31,   -24,   -57,   -18,   -32,   -20,    22,   -14,   -69,   -38,   -28,    -9,    -8,   -74,   -31,   -32,    -4,    25,   -15,    27,    13,    14,   -38,     9,    57,    15,   -33,   -73,   -42,    -2,   -18,    10,   -17,    25,   -31,   -13,   -84,  -112,   -26,    -2,    -1,   -29,    -3,    -9,     6,    28,    11,   -56,   -15,   -25,   -43,   -32,   -32,   -14,   -28,   -19,   -43,     1,   -17,    24,   -28,    37,   -43,   -34,   -65,   -66,     3,   -34,    -6,   -46,    10,   -19,     8,    -5,   -29,   -50,     0,   -57,   -79,   -64,   -44,   -37,   -50,   -50,    40,    44,   -23,     4,   -13,    -8,   -43,  -103,   -63,  -112,   -19,   -21,   -17,   -26,    -5,    16,   -47,   -18,     4,     8,   -10,   -24,   -50,   -34,   -58,   -44,   -12,   -38,   -56,   -15,   -23,   -10,    43,   -40,   -56,   -81,    15,   -50,    -5,    -4,    -3,   -34,    17,     4,     0,   -60,    -4,    13,    28,   -40,   -34,   -37,    -8,   -47,    -6,    -6,     3,     2,    35,    59,   -36,    16,    36,   -37,    15,   -67,    -4,     8,     9,   -30,   -23,  -110,   -85,   -72,  -100,   -59,    -5,    -1,   -16,    -3,   -11,   -43,   -26,   -53,   -70,   -37,    48,   -19,   -64,   -24,    12,   -26,   -37,   -17,    -9,     3,    -4,   -34,   -25,   -24,    -7,    46,    36,   -18,    -7,    67,     9,   -62,   -31,    -4,    24,    38,    -1,    20,   -46,   -25,   -43,   -65,   -45,   -68,   -46,   -28,    -4,    -1,     3,     5,   -28,   -30,   -62,   -80,   -78,   -96,  -140,  -110,   -55,   -48,   -48,   -53,  -138,   -73,   -45,   -58,  -110,   -83,   -50,   -31,   -30,    -2,    -9,    -1,    -9,    -2,     5,     5,    -5,     0,   -10,    -7,   -34,   -60,   -67,   -41,    -9,   -21,   -50,   -59,   -73,   -45,   -48,   -30,   -37,     4,    -8,    -5,     1,     0,    -1,     7,    -6),
		    29 => (    8,     0,     4,   -10,    -1,     1,    -8,     8,     0,     7,   -10,     1,     9,     7,    -9,     7,    -2,    -4,    -4,    -6,    -4,    -8,    -3,     6,    -2,     0,    -3,    -9,     1,     2,     9,     0,    -6,     5,     1,     3,     6,    -9,    -1,   -16,   -25,   -16,     2,   -11,   -31,   -42,   -35,   -20,     8,   -16,    -3,    -3,     6,    -6,     4,   -10,     1,     6,    -6,   -13,   -16,     1,    -2,   -19,    -7,   -17,   -18,   -33,    -2,    -3,   -60,   -44,   -36,   -11,   -10,    -8,   -74,   -26,   -48,   -29,   -13,    -6,     0,     6,    -3,     3,     5,   -13,   -26,   -62,   -59,   -53,   -68,   -67,  -119,  -120,   -80,   -92,  -174,   -69,   -86,  -127,   -94,   -64,  -101,  -109,   -73,   -40,   -27,   -13,    -5,     4,     6,    -6,   -28,   -28,   -33,  -104,  -145,   -53,   -65,   -79,   -38,   -24,   -17,   -12,   -29,    13,   -16,   -59,   -19,  -147,  -127,   -38,   -54,   -29,   -21,   -72,   -47,    -7,     3,    -8,    -5,   -13,   -10,   -39,   -50,   -48,   -26,     7,    11,    41,     9,    29,    20,   -10,    11,    25,    47,    48,    17,   -65,   -67,   -62,   -21,   -49,   -34,     5,    -8,     7,    -8,   -42,   -37,   -69,   -25,   -50,     0,    45,    20,   -24,   -44,     9,    12,    26,    16,    -3,    60,    38,    46,   -14,   -21,    26,     8,   -17,   -34,   -60,    -4,    -9,   -46,   -34,   -47,   -55,   -69,   -58,    -1,    16,     9,   -23,     1,   -37,    -5,   -23,   -15,    -4,    -1,    16,   -22,   -41,   -47,   -12,    10,    28,   -40,   -21,   -31,   -38,   -19,   -15,   -16,   -51,    13,   -11,    20,    49,    31,   -12,   -12,    -7,   -22,   -12,    -8,   -17,     6,   -26,   -67,   -54,   -61,   -35,    18,    -7,   -46,   -16,    -7,   -37,    19,    57,    57,    23,    27,     0,    22,    53,    -7,    -8,   -16,   -26,   -27,   -31,    15,    40,    38,   -19,    -9,   -20,   -53,   -81,   -47,   -66,  -106,   -40,     4,   -49,   -43,    32,   121,    66,    71,    44,    10,    11,   -16,   -20,    16,   -20,   -21,    17,    88,    71,     8,   -24,   -27,   -18,   -37,   -27,   -32,    17,   -31,   -19,     6,   -96,    -8,     3,    65,    68,    63,    10,   -34,    -7,   -10,    11,   -12,    29,    44,    26,    98,    67,     5,   -49,   -26,    -7,    24,    21,     7,    54,   -13,   -28,     7,   -24,    14,   -21,    49,    39,    54,   -15,    -5,   -12,   -17,    -6,    -4,    20,   101,    71,    41,     8,    15,   -15,    19,    -7,    12,    18,   -26,   -33,   -38,   -26,    -4,   -27,   -16,   -26,    37,    57,   -10,     1,   -24,   -27,   -13,     9,     3,    75,    92,    98,    45,    12,    20,   -23,     2,    16,    24,    12,    -4,   -15,   -31,   -14,     2,   -33,   -41,   -30,     7,     8,    36,     6,     7,    12,   -11,     9,    35,    90,   103,    72,    68,    22,    28,    30,    24,    -2,   -25,   -42,   -31,   -31,     4,     4,     8,     8,   -69,   -26,   -13,   -16,    23,   -10,   -38,   -18,   -16,    -3,    30,    96,    96,    56,    59,    19,    56,    31,    47,    19,   -31,   -64,   -66,   -28,    -7,   -17,     5,   -14,   -64,   -55,   -17,   -32,    40,    15,    28,   -26,    33,    23,    44,    46,    83,    59,     6,    28,    57,    50,    74,     3,   -18,   -36,   -85,   -62,   -16,   -24,    -5,     1,   -60,   -11,   -25,   -55,    42,    53,   -11,    18,     6,    68,    49,    31,    76,    28,    13,    31,    45,    30,    51,    -2,   -14,   -36,   -82,   -32,   -49,   -19,    26,    -5,   -63,   -26,   -62,   -65,    49,    60,    56,    37,    27,    10,    -5,    13,    11,    18,     6,    79,    31,    52,    35,   -23,    -4,   -51,   -96,   -46,   -50,   -49,     0,    -1,   -83,   -21,   -73,   -66,    29,    59,    40,    46,    25,    13,   -13,     4,   -36,     7,    67,    49,    28,     5,     2,     3,    21,    -7,   -26,   -17,   -23,   -20,     2,    -9,   -77,   -31,   -73,   -45,   -35,    13,    45,    10,   -21,     3,    20,   -20,   -37,   -11,    29,    16,    -2,     1,   -10,   -23,   -21,     1,    -9,    25,   -27,     5,     1,     4,   -70,   -30,   -60,    -4,   -25,     6,   -39,   -15,   -29,     6,    17,   -32,   -35,    30,     4,     2,   -42,   -30,   -15,   -19,   -35,   -15,    17,    -2,   -63,     1,    -6,    -1,   -49,    38,   -39,   -60,   -19,   -29,   -30,   -12,   -11,     6,     8,   -53,   -15,     8,   -46,   -52,   -59,   -30,   -26,   -57,   -40,   -32,    13,   -45,   -18,    -4,     0,     5,   -34,    11,   -25,   -37,    -9,   -49,   -55,   -51,   -47,    -5,    15,    -6,     5,   -30,   -58,   -44,   -43,   -36,    38,   -39,   -43,   -57,     9,   -13,   -34,    -5,    -8,     6,   -44,   -59,   -18,    13,   -49,   -46,   -21,   -23,   -19,   -18,     6,     1,   -26,   -70,   -56,   -36,   -46,   -42,   -26,   -24,     0,   -24,     2,    -6,    -4,    -5,    -3,     6,    34,   -21,   -10,   -16,   -53,   -79,   -46,     2,   -30,   -26,     0,   -18,   -20,   -67,     6,   -18,   -13,   -43,   -26,   -25,    -1,    35,   -18,     2,   -13,     3,    -8,    -6,    -2,    57,   -27,   -58,   -42,   -47,   -38,   -31,   -36,    -1,     8,    -4,     0,   -15,    45,    29,    25,   -54,    -3,     9,    -8,     9,     9,     7,     8,    -6,    10,    -5,    -5,    -6,    -5,   -16,    27,    33,    15,    22,    13,     6,     2,    39,    17,   -12,    -8,   -34,    -1,     1,   -17,   -35,   -14,   -34,     0,    -1,    -1,    -5),
		    30 => (    9,    -9,    -4,    -2,    -7,    -4,     7,     4,     0,     2,     0,    -8,     5,    -2,   -18,    -1,     0,    -3,    -6,    -4,    -9,    -3,    -8,     5,     3,     9,    -9,     8,   -10,    -6,     0,     1,     8,    -1,    -5,   -43,   -39,   -63,   -40,    32,    14,    10,   -26,    40,    55,    42,   -23,   -13,    -7,   -13,   -12,    -7,    -2,     3,    -3,     2,     1,    -1,     6,    57,    51,     1,    -7,    -7,   -38,   -50,   -75,   -97,   -55,   -83,   -71,  -122,  -105,  -113,   -73,   -62,   -56,   -48,   -68,   -41,   -23,   -21,     0,    -5,     5,     5,     2,    36,   -18,   -37,   -34,   -58,   -53,   -19,   -64,    11,    33,    44,   -24,   -83,   -28,   -20,   -74,  -100,   -25,   -44,   -40,   -44,   -57,    -7,   -31,    -2,     8,    -4,   -33,   -68,   -15,   -85,    10,     2,   -11,     6,    19,    -7,    13,    10,   -32,   -36,   -70,    -3,    -1,    31,     3,    -2,   -25,   -44,   -81,   -97,   -40,    -7,    -9,    -4,   -16,   -49,   -11,   -19,    31,    20,    -2,   -26,    18,   -16,   -53,   -54,   -20,   -37,   -47,   -11,    22,    23,   -36,   -34,     6,   -59,    -5,  -122,   -74,    -9,    -7,     1,   -12,    -3,   -13,    -1,     4,    33,    17,   -86,    -3,   -29,   -61,     8,   -19,   -12,   -20,    -4,    -1,     8,   -22,     1,    18,    -3,    26,  -103,   -29,    -4,     8,   -22,    -3,   -32,    -9,   -10,    -1,    -1,   -43,     3,   -10,    51,   -16,    37,    -5,   -29,    12,    -2,    27,    41,    15,    50,    28,    67,    14,    -1,   -63,     0,    85,   -64,    42,    12,   -26,   -69,   -55,   -25,   -13,    -1,    45,     0,    17,    -8,     6,    57,    52,    61,    13,    51,    53,    50,    51,     3,     6,   -53,   -91,   -30,    -8,    -4,    68,   -51,   -47,   -31,   -39,   -46,    -3,    22,    15,     2,    -2,    -6,    30,    24,    35,    25,   -26,     9,    66,    31,    -8,     1,    17,   -75,   -41,   -12,   -17,   -12,    60,    31,   -61,   -32,    25,    -3,    -9,    -9,     7,   -18,   -23,   -14,     1,    45,    20,    48,     6,    -2,    25,    27,     9,   -40,   -34,   -79,   -99,    -6,    -7,    68,   -51,   -14,  -112,     3,    17,    15,    18,   -33,   -22,   -49,   -43,     8,   -25,   -37,   -22,   -19,   -26,   -31,     3,    56,    12,   -64,   -83,   -78,   -65,    -8,    -2,    12,   -46,   -12,   -22,    12,    38,    28,    -3,    16,   -10,   -62,   -23,   -12,   -62,   -35,   -12,   -23,   -29,   -20,    -3,    38,    46,     0,   -43,   -21,   -36,   -26,    -6,    17,     0,    34,    51,    18,    72,    41,     2,    32,     0,   -36,   -14,   -55,   -25,   -60,   -17,    27,     8,    18,   -54,    22,     2,    -3,   -47,   -21,   -43,   -42,     5,     0,    -3,   -10,    86,    96,    98,    46,    33,    45,    52,    18,     0,   -40,   -47,    -6,   -49,    -4,     4,    26,   -19,   -65,    -2,   -28,    24,   -62,   -86,    -1,     2,    -1,   -40,   -32,    62,   110,    30,    63,    73,   106,    64,   -20,    52,   -36,   -36,   -20,   -30,     1,    -7,   -21,    -8,   -45,     7,    15,    -3,   -48,   -94,   -46,    -6,    -2,   -23,   -75,    67,    70,    44,    44,    86,    93,    37,    75,    54,   -32,    11,    21,   -27,   -18,    -3,   -30,   -21,   -55,   -63,    36,   -68,  -103,  -132,    71,     5,    -6,   -23,   -96,    26,    28,   -18,    39,    21,    42,    58,    62,     2,   -31,   -14,    -9,    -5,     5,     4,     2,     1,   -64,    19,   -20,   -70,   -77,   -68,   100,    -7,    -7,   -16,  -107,     0,   -13,   -14,     2,    45,    21,    31,     7,    25,    -6,    -8,     4,   -18,   -33,   -29,   -26,   -27,   -25,     1,   -24,   -34,   -62,   -69,   -25,     2,    24,   -27,   -75,   -34,   -11,   -15,   -10,   -17,   -55,   -28,   -10,    44,    10,    -6,     0,   -21,   -42,   -12,     2,   -29,     2,     6,   -32,   -30,  -108,   -58,   -25,     3,    35,   -25,   -89,   -22,    -4,   -15,   -33,   -51,   -61,   -21,    17,   -10,    14,    39,    19,    -7,   -29,    -1,   -29,   -26,   -18,   -18,   -22,   -38,   -97,     1,    -8,    -8,     6,   -77,   -52,   -56,   -13,    29,    10,   -25,   -25,   -18,   -14,    20,    57,    42,    51,    48,    12,   -22,   -66,   -56,   -22,     7,   -22,   -29,   -28,    63,    22,    -1,     6,  -105,   -32,   -98,   -31,     0,    20,    61,    -4,    24,    24,    83,    33,    66,    56,     7,    -6,   -30,   -35,     4,    21,    35,    38,   -43,   -27,    37,    18,     3,    -7,   -26,  -105,   -85,   -21,    22,   -14,    -2,   -24,    13,    13,    21,    23,    39,     9,    32,   -31,   -28,   -26,   -24,    25,   -16,   -35,   -44,   -31,   -77,     1,    -4,     1,   -11,   -23,   -13,    32,   -28,   -47,   -58,   -93,   -90,   -59,    24,    68,    64,    58,    52,    -7,   -24,   -94,   -67,   -30,   -47,   -57,   -32,     2,    -7,     9,     5,     8,    -1,   -31,  -164,  -130,   -31,   -11,   -13,  -103,   -81,   -55,    -8,   -23,   -31,   -47,   -14,    -7,   -65,  -106,   -78,   -74,   -42,   -19,     4,    -2,     6,    -4,     2,     2,     7,    -4,   -83,   -72,  -104,   -35,   -50,   -83,   -78,   -41,   -46,   -50,   -85,   -70,   -50,  -115,  -113,   -52,   -71,   -79,   -36,   -44,   -14,    -5,    -1,    -4,     2,   -10,     2,    -4,     4,     1,   -11,    -6,   -30,   -20,     6,     5,     5,   -27,    -1,     2,   -17,   -18,   -26,   -25,   -11,   -37,   -39,   -34,    -3,     7,    -9,    10),
		    31 => (    7,    -9,    -3,    -4,     2,    -8,     4,     5,    -5,    -6,     4,    -9,     5,     9,    -6,     7,    -9,    -9,     8,    -3,    -2,   -10,    -8,    -8,     2,     6,     7,     9,    -4,    -3,     5,     7,     6,    -6,    -4,   -10,    -4,     0,   -14,   -14,   -12,   -39,    18,    21,     3,   -22,   -11,     6,    -4,     5,    -1,     1,     8,    10,     5,    -4,    -9,    -7,    -3,     0,    -9,     4,    -7,     9,   -30,   -47,   -32,   -32,   -65,    25,   -16,    -4,    23,     5,    15,    52,    51,   -88,   -73,   -44,   -16,   -18,     9,    -9,     2,    -2,    42,    32,    -1,   -42,   -59,    29,    44,    44,    -5,   -59,   -25,   -34,     3,    42,     7,    -2,    -3,    46,    38,   -21,    -8,   -26,   -40,    -9,   -10,     2,    -5,    -6,    48,    40,    32,    50,     0,     3,    29,     9,    34,    -5,    -4,    27,    -4,    -5,     4,    52,    71,    49,    -6,   -10,     9,    -7,   -27,   -50,   -65,   -47,     7,     8,    24,    14,    53,    62,    45,    48,   -20,   -48,   -20,   -23,    -2,    -9,   -30,    -2,   -15,   -19,     3,    52,    22,   -16,   -16,    30,   -17,   -70,   -50,   -48,     3,    -9,   -41,    16,    59,    51,    58,    39,   -24,   -27,    -3,   -14,   -36,   -22,   -25,   -36,     9,     2,    10,    20,    14,   -33,   -31,     3,    -4,   -30,   -70,    -8,     3,   -25,   -68,   -26,   -95,     7,    52,    56,   -37,   -26,   -34,   -13,     3,    18,    18,     4,     6,   -45,    -5,    20,    20,   -13,    -1,    36,   -12,   -58,  -127,   -73,     3,   -65,   -72,   -92,   -89,   -39,    19,    -1,   -45,   -31,    -5,    -9,    51,    44,    54,    -7,   -12,   -20,    19,     8,   -40,   -21,    27,     6,   -12,   -52,  -178,   -36,     7,   -19,   -59,  -101,   -81,   -41,   -51,   -21,   -46,   -34,    -9,    14,    60,    62,    43,   -16,    -2,   -22,     2,     9,   -29,   -56,     2,   -20,   -45,   -51,   -80,   -45,     0,   -18,   -57,   -29,   -76,   -58,   -58,   -31,   -40,   -71,   -38,   -19,    72,    62,    37,    -6,   -13,    18,   -21,   -29,   -37,   -42,   -55,   -58,   -50,   -33,   -27,   -11,    -7,    12,    -6,   -44,   -48,   -61,   -80,   -76,   -71,   -49,   -56,   -46,     0,    53,    19,    31,   -25,   -12,   -19,   -38,     8,   -35,   -19,   -67,   -68,   -37,   -40,    53,    -1,    -9,   -85,   -26,   -11,   -52,   -47,  -102,   -71,   -58,   -30,   -29,     6,    56,   -12,     3,    39,     8,   -19,   -17,    20,   -50,   -48,   -28,   -49,   -14,     7,    45,     5,     3,   -72,    24,   -22,   -61,   -34,   -60,   -48,   -37,   -32,   -45,     2,    -8,    20,    24,    62,    43,    -5,   -17,   -18,   -91,   -71,   -69,   -66,     8,     7,    -5,    -9,    -2,    18,     8,   -34,   -41,   -51,   -33,   -47,   -27,   -50,   -44,    14,   -10,     4,    16,    14,    11,   -22,   -57,   -18,   -64,   -49,   -36,   -49,   -47,   -18,    -6,     2,     1,    12,   -34,   -66,   -54,   -56,   -64,   -44,    -9,   -10,    -7,    -3,    21,    17,     7,    26,    25,    12,   -26,   -56,  -104,   -88,   -67,  -169,   -83,   -46,   -32,    -8,    -1,    20,   -72,   -64,    -6,   -24,   -45,   -25,    14,   -19,   -28,   -14,     8,     7,    -5,    24,    -1,   -12,   -14,   -41,   -72,   -41,   -31,    14,   -54,   -32,   -40,     9,     0,   -28,   -77,   -35,   -25,   -42,   -79,    14,     2,    26,    28,   -24,   -23,    48,    36,    28,    14,    -4,    -1,   -17,    23,    21,   -14,    18,   -28,   -44,   -43,    -6,     5,     7,   -87,   -55,   -56,  -117,   -77,    -2,    33,    38,   -18,   -45,   -27,    14,    59,    48,   -18,    13,   -57,   -31,   -15,   -13,    17,    18,    -5,   -39,     3,    -9,    -2,   -17,   -91,  -101,     5,     4,    -5,    30,    42,    41,   -13,   -27,    14,    24,    22,    21,   -23,   -32,   -69,   -52,    -1,    38,    39,    52,    23,   -50,   -12,    -7,     4,   -33,   -92,   -18,    51,    60,    82,    15,    54,    49,     5,    25,    34,    21,    13,    13,   -34,    13,   -17,    17,    25,    51,    44,    51,     6,   -16,     0,    29,    18,   -12,    -4,   -17,    29,    44,    56,    75,    74,    35,     1,    30,    67,     2,   -28,    11,   -22,    12,    -5,    27,    35,    40,     9,    12,    23,   -32,     5,    13,    16,   -26,    -9,   -11,    46,    54,    54,    44,    72,    34,    31,    30,    61,   -63,   -41,    -8,   -15,    11,    28,    52,    37,   -38,   -16,    28,     2,     7,     1,     2,     5,   -14,   -14,   -24,    16,    16,     2,    16,    73,    44,    40,    46,    -4,   -54,   -30,   -46,    18,   -18,   -16,    23,     3,   -16,   -45,   -52,   -39,    64,    -9,     3,    -7,    10,   -12,   -41,     5,   -20,     6,   -13,    25,    22,   -52,   -14,    -5,   -59,   -56,   -56,    11,   -12,   -53,   -19,    27,    -6,   -65,   -64,     6,    10,    10,   -10,     2,     0,   -16,   -45,   -74,   -42,  -100,     9,   -41,   -10,   -43,    33,    -1,   -51,   -63,   -74,  -103,  -117,   -89,  -162,   -59,   -39,   -28,   -14,   -16,   -18,    -3,    -2,    -6,    -2,   -13,   -51,  -108,  -153,  -165,  -116,  -107,    16,     3,   -66,   -65,   -62,   -66,   -43,   -84,   -44,   -14,   -30,   -33,    -8,   -11,    -2,    -3,    -5,     7,    -8,    -2,    -2,     6,    -7,   -13,    -1,     7,     5,    -8,   -63,   -52,     5,   -15,   -46,   -17,   -20,    -5,     1,     1,     9,    -8,    -5,     7,     3,    -9,     7,     9),
		    32 => (   -1,     8,     2,    -6,    -5,    -1,     1,     5,     1,    -4,    -3,    -9,   -20,   -15,    10,     0,     0,    -8,    -2,     1,    -6,     6,     8,    -3,     3,     5,     7,     3,     0,    -9,    -3,     9,    -2,    -1,     8,     3,   -39,   -25,   -21,    -9,   -15,   -17,   -60,     3,     9,   -15,    -9,   -48,   -24,   -15,   -27,    -3,     8,   -10,    -4,    -2,     4,    -7,    -3,   -11,   -13,    -5,    -4,   -29,   -12,    10,    13,   -14,    10,   -14,    -9,   -23,   -30,   -37,    13,    -3,   -41,   -16,   -14,     3,    -1,    16,     9,     1,    -6,    -9,    -5,   -17,   -34,    27,    17,    13,   -29,   -28,   -52,   -31,   -57,   -72,   -43,   -23,   -75,   -90,   -62,   -18,   -58,   -62,   -23,    -6,    -1,    -5,     4,    -4,   -10,    -5,   -17,   -14,    37,    45,    61,    46,    48,    34,     1,    13,    23,   -25,   -29,   -15,   -15,   -55,   -18,    -9,   -46,   -43,   -60,   -29,   -22,   -15,   -29,    -2,    -8,   -10,    13,    12,    16,    -3,    13,    11,    22,    38,    25,    22,    -9,   -33,   -48,   -66,   -14,    -9,   -38,   -31,   -26,   -15,   -43,   -32,    -6,     2,   -21,   -19,     5,    -3,   -25,    38,    36,    37,    59,    -3,   -12,     3,    -4,     5,   -25,   -20,   -24,   -26,    -5,    -1,    -4,     2,   -35,   -15,   -12,   -41,   -17,   -30,   -16,    -1,     5,    -1,     6,    59,    59,    20,    59,    28,    57,    -4,   -26,    -3,    28,    -8,   -41,   -13,   -12,   -38,    -2,   -14,   -19,   -17,   -33,   -87,   -54,   -27,   -34,   -14,   -25,    15,     2,    22,    29,    20,    51,    40,    29,    32,    10,    -8,    25,   -14,    27,   -14,   -62,   -26,   -38,   -14,   -19,   -52,     3,   -31,   -61,   -33,   -52,   -18,     8,   -12,    -7,   -17,     5,    30,     8,    11,   -11,   -19,   -64,   -36,   -24,   -29,    10,     3,   -16,   -44,   -16,    -5,    -2,   -13,    14,   -15,   -55,   -27,    16,    -5,     0,    -9,     5,   -59,   -32,    -1,    24,     2,   -18,   -55,   -46,  -106,  -101,   -46,    -9,     0,   -15,   -20,   -16,   -15,    17,   -35,   -39,    -3,   -24,   -22,   -27,    -5,     9,    -9,   -25,   -35,   -43,   -36,   -12,   -15,   -20,   -54,   -14,   -30,   -96,   -48,   -25,   -13,    -3,   -33,   -22,    -5,   -16,   -35,    -4,   -17,    -2,     6,   -67,   -15,     5,    -3,    -9,     2,   -54,   -97,   -71,   -63,   -53,   -53,   -36,   -15,   -31,   -51,   -28,   -50,   -22,    -9,   -36,     2,   -27,   -22,    30,     9,    58,    18,   -11,   -10,    -7,     0,    -4,   -16,   -16,   -91,  -110,   -96,   -68,   -64,   -42,     4,    -3,   -10,   -21,   -59,   -35,   -40,   -27,    -1,    22,   -13,    42,    60,    83,    47,     5,   -19,     9,   -19,   -19,   -11,   -42,   -75,  -108,   -76,   -60,   -34,    31,    13,   -24,   -52,    -6,   -31,   -42,   -61,   -15,    48,     7,    14,    40,    26,    18,     9,    23,    39,    10,   -26,    29,    27,   -32,   -71,   -61,   -12,    -2,    15,    34,    -6,    14,    34,    29,     2,   -17,     8,    12,    78,    61,    31,     6,    37,    52,    49,    35,    60,    -5,   -13,    38,     5,   -25,   -75,   -10,     5,     1,     2,    14,     7,    10,     4,     0,   -18,   -55,     8,    44,    63,    12,    43,    46,    49,    13,    80,    24,    30,     8,    -8,    52,   -12,   -42,   -16,    14,    39,    21,    48,    -4,     0,   -32,   -30,    18,   -12,   -66,    40,    63,   -12,    -6,    28,    -9,    -7,   -54,    48,    -8,    36,     3,     7,    10,    41,   -59,     6,    27,    22,    22,    -9,   -30,   -21,     9,   -36,     3,   -23,    19,    51,    34,   -35,   -46,   -15,   -25,   -23,    22,    61,     9,    85,    -7,   -40,   -24,   -20,   -59,     1,    14,    40,    13,   -23,   -32,    -6,   -17,     2,   -18,    -3,    34,    41,     4,   -31,   -49,   -60,     7,   -36,   -54,     3,    56,    64,    -9,   -37,    -3,    -5,   -42,     0,    23,    22,    17,   -31,   -43,     2,     7,    28,   -21,    -2,    11,   -10,   -10,   -32,   -47,   -49,   -37,   -46,   -67,    -9,    12,     5,    -1,    10,    13,     9,   -62,   -38,   -12,   -36,    24,   -10,   -13,    12,    -1,    13,    -2,    27,    38,     1,     7,   -25,     0,     8,   -27,     6,   -40,   -10,    17,   -10,    -1,     5,    -4,    27,   -47,   -76,   -38,   -40,   -32,   -30,   -17,    38,     8,    46,    41,    -3,     1,    15,    -2,   -23,    10,     4,   -50,     5,     3,    -6,   -27,     0,     1,     3,    -6,    33,   -46,   -67,   -47,   -34,   -34,     3,    21,    18,    57,    35,     8,     6,    17,    26,   -21,   -17,   -22,   -12,    11,    20,    11,    20,   -31,     2,     2,     4,   -50,   -38,   -77,   -52,   -68,   -28,   -51,   -66,   -59,   -45,   -41,   -44,   -16,   -21,   -60,   -16,     8,    19,    12,   -21,    -2,    20,    33,    -5,     5,     4,    -4,    -6,     3,    -5,   -14,   -14,   -12,    -7,   -32,   -72,   -98,   -72,   -68,  -122,   -10,    -7,   -35,     3,   -21,    27,    29,    22,   -29,    -7,    12,    10,     6,    -1,     4,    -9,     5,    -6,    -3,   -34,   -33,   -29,   -26,   -59,   -10,   -17,   -31,   -30,   -42,   -27,   -52,   -66,   -53,   -31,   -30,   -22,   -32,     4,     1,     2,    -6,     1,   -10,     3,     7,    -9,    -9,     3,     6,    -2,   -10,    -2,   -21,   -16,   -21,   -37,   -28,     8,     0,   -17,    -9,    -9,   -13,   -28,   -26,    -2,    10,    -1,    -5,    10),
		    33 => (   -7,    -2,     0,     9,     5,     7,     1,     8,     7,    -4,     7,     0,     1,    -6,   -10,     1,     3,   -10,    -9,     4,     6,     8,    -8,     3,     2,    -6,     2,    -4,     0,     5,    -3,    -8,    -8,    -3,     2,     3,     7,   -10,   -11,    -3,    -8,   -13,    -8,    -9,    -4,   -18,    -6,     8,     1,     0,    -2,     6,    -4,    -5,     7,     0,   -10,     3,     0,     2,     0,     8,    -7,    -2,   -25,   -32,   -13,   -13,   -39,   -35,   -59,    -1,   -20,   -11,   -20,   -16,   -34,   -15,   -17,   -20,     0,     6,   -10,    -9,     4,    10,    -1,    -6,     3,     3,     5,    -6,    -3,    -1,     4,     3,    -3,     0,     3,   -10,   -24,   -20,   -12,   -24,    -9,    -5,    -8,   -26,   -31,   -22,    -4,     0,    -5,    -3,     1,    30,    -9,    -8,    -3,    -3,    -9,    -2,    -1,     1,   -17,   -16,   -10,   -10,    -2,    -5,   -26,   -17,   -24,   -14,    -3,    -1,   -67,   -32,   -19,     4,     2,     0,    -1,    13,    31,    -4,    10,    -7,   -21,   -35,   -28,   -32,   -39,   -14,   -34,   -12,     2,    26,    32,    21,     1,   -18,   -24,   -20,   -16,   -55,   -14,     2,    -3,    -5,    25,    -9,    24,    23,     8,     8,    -3,     6,    13,     7,    18,   -11,   -17,   -17,   -30,   -43,     4,    10,   -12,   -40,   -33,   -23,    -4,    -4,   -38,    -7,     1,     8,    42,     4,   -11,    23,     3,    25,    24,    27,     8,    23,    -2,   -28,   -21,   -37,   -33,   -15,   -31,   -69,   -38,   -28,   -29,   -28,   -22,   -11,   -56,   -13,    -9,    15,    37,    31,    22,    -4,    27,    32,    27,   -17,     9,   -19,   -30,    -5,    10,    14,    -2,    18,     3,     0,   -33,   -20,   -11,    -7,   -11,   -29,   -46,     2,     8,   -41,    86,    20,    26,    -2,    46,    17,     1,    26,    20,   -39,   -27,     4,    29,    -4,   -56,     8,    22,    -6,     1,    19,   -24,     0,   -49,   -53,   -23,     0,     9,   -35,    78,    23,   -10,   -23,    22,     0,   -26,   -48,   -35,   -31,     0,     6,    41,   -40,   -52,   -10,    10,   -11,    11,    17,    -6,    -6,   -44,   -20,    -5,    -5,     2,    -6,   -32,   -26,   -14,   -29,   -49,   -40,   -49,   -58,   -22,     1,    13,   -21,   -38,   -37,    -8,    -4,    11,     3,     9,    15,    15,   -10,   -21,   -44,   -15,     1,     9,     1,   -39,   -17,   -17,   -48,   -58,    -2,   -13,   -18,    -9,     0,   -23,   -71,   -32,    -2,    -3,    21,    24,    -8,    -3,     4,    -1,   -14,   -17,     7,     1,    -7,     4,     5,   -25,   -15,    -4,   -25,   -34,     0,     8,    11,   -24,     3,   -21,    16,    -8,    -8,   -17,    23,   -14,   -16,   -33,     0,     9,   -16,   -24,   -20,   -26,   -19,    -4,    27,   -12,   -19,     3,    -5,   -16,   -36,   -19,   -25,    -2,    -8,   -26,     9,    27,    18,     7,   -29,   -45,   -27,   -40,   -15,   -15,    -7,   -18,   -56,   -28,   -20,    -5,    12,   -10,   -23,    19,   -24,   -25,   -11,     2,   -18,    -2,    -1,     6,    12,    15,   -15,     4,    -3,   -27,   -40,   -21,   -20,    19,    -1,   -14,     0,    -8,     0,    -6,     1,   -13,   -17,     3,   -24,    -6,   -21,    -6,    37,     6,   -10,   -10,     5,     3,   -16,     2,   -39,    -4,     0,   -12,    -3,    19,     1,   -11,     6,   -39,   -27,    -9,    13,    -9,    32,     5,    -8,    -3,   -13,     1,    29,    -8,    15,    13,    -8,   -15,     3,   -11,   -45,   -40,   -23,   -13,    -2,    20,    -3,   -25,   -10,    -5,   -12,   -14,     3,     2,    25,    25,    19,    -1,   -30,    -1,    23,    49,    -8,     8,    38,    -6,   -15,   -19,   -43,   -43,   -22,    -8,    21,    33,     9,   -21,   -15,    -6,   -21,   -10,    -4,     8,     6,    32,    20,     7,   -14,    -8,    -3,    19,   -18,    17,     4,   -23,   -16,   -28,   -24,   -25,   -23,    14,    11,    44,    34,   -24,   -11,   -18,   -14,    -3,     3,    -9,    10,    12,    14,    20,   -13,   -25,     7,    -3,   -56,    -5,    27,    -1,   -28,    -7,   -16,   -24,     5,   -11,    15,    41,    34,   -35,   -28,     1,   -10,    -1,     0,     4,    17,    20,     5,    -5,   -34,   -49,   -10,   -26,   -52,   -51,   -33,   -45,   -10,    14,   -21,    -5,     4,    -3,     3,     1,    34,   -25,   -27,    -2,     7,   -14,     1,     3,    13,    37,     9,    -1,   -21,   -51,   -27,   -20,   -56,   -75,   -44,   -68,   -47,   -19,   -15,    37,    46,    19,   -18,    -3,    34,   -10,   -25,    -7,     8,     2,     6,    22,   -10,    -7,   -12,   -10,   -11,   -32,   -55,   -16,   -12,   -38,   -34,   -45,    -7,    31,    13,    21,   -18,     2,     9,    17,     3,   -19,   -27,     8,   -10,    -3,    -1,   -19,    -1,   -16,   -16,   -11,    14,   -30,   -39,   -50,    -8,   -58,   -20,    27,    63,    39,     1,   -19,   -11,     3,    -8,   -22,    14,   -39,   -20,   -11,    -5,    -1,     1,    15,   -17,   -44,   -48,   -15,     7,    27,     0,   -17,   -16,    11,    62,    89,    14,    28,   -22,    -3,     3,    23,    -2,   -37,   -94,    -6,    -1,     1,     3,     2,     6,    -4,   -33,   -36,   -35,   -57,   -41,   -39,   -60,   -32,   -28,    34,    61,    43,    -8,   -21,   -19,   -17,   -21,   -32,   -25,   -49,     8,     7,    -2,    -2,     8,     0,     9,    -2,    10,     2,     2,   -10,     8,     8,   -34,   -34,   -14,   -19,   -19,   -15,   -35,    -1,     3,   -12,    -8,   -18,   -20,    -3,    -2,     3,     2,     7,     0),
		    34 => (   -7,    -6,    -5,     4,     0,     2,    -9,     7,    -3,     8,    -9,    -6,    -2,    -6,     2,     7,     4,     8,    -1,     4,    -4,    -5,    -2,    -1,     7,    -7,    -6,     6,    -7,    -9,    10,    10,     5,     0,   -10,   -20,   -19,     5,    -9,     3,     5,   -38,   -30,    -9,    -6,   -16,     1,     5,    -3,    -8,   -14,    -8,     1,    -7,    -5,     1,     8,    -6,    -8,    -7,   -22,     3,   -17,   -32,   -14,    -6,   -17,   -17,    -7,   -24,   -30,   -14,    -8,   -26,    -6,    -2,   -30,   -11,   -11,    -6,     5,    -1,     2,     8,     6,    -6,    -2,    -9,   -13,   -10,   -45,   -23,   -36,   -19,    -7,   -13,   -18,   -35,   -57,   -57,   -35,    13,    -2,   -24,   -11,    -2,    -7,    -7,     2,   -11,    -1,    -3,     5,    -3,    -2,   -12,   -19,    -6,   -21,   -17,    -7,   -13,   -17,   -19,   -25,   -46,   -66,   -34,   -19,   -21,   -53,   -42,    -9,   -32,   -40,    -9,    11,    -5,    -9,   -11,     5,    10,     7,   -11,   -15,    -3,   -19,    -8,   -25,   -31,    -9,   -41,   -65,   -38,     0,    26,   -14,   -82,   -73,     3,   -25,   -12,   -16,    29,    33,     4,   -29,    -7,    -6,    -2,     7,   -24,   -15,    33,   -26,    -5,   -26,   -24,   -38,   -26,   -12,     0,    60,     3,  -123,  -147,   -48,     8,    55,     2,    34,   -31,    13,   -13,    33,   -52,   -10,   -55,     1,    -8,   -11,    47,   -10,    -8,     6,   -23,   -64,   -38,    25,    22,    22,  -100,  -132,  -102,   -17,    27,    12,    -7,    32,    22,    14,    14,     2,   -27,   -18,   -48,    12,    -9,    -8,     7,     6,    26,    -4,   -19,   -68,     9,    31,    36,   -46,   -55,  -113,   -29,     8,     4,    14,    -5,    30,    10,    22,    -4,   -18,   -41,     7,   -40,    16,   -10,     4,   -19,   -31,   -12,   -33,   -46,   -39,    49,     6,    -2,   -29,  -100,   -75,    -9,    14,    26,    18,     4,    11,     6,     7,   -21,    -4,   -20,    -9,    -7,   -31,    -3,    -3,   -47,   -41,   -10,   -41,   -44,    -9,    49,    -1,   -33,   -66,   -31,   -22,   -15,   -10,     3,   -10,   -47,   -71,     5,   -47,    -3,   -17,   -18,    -7,    -5,   -33,   -19,   -31,   -36,   -21,   -43,    -9,   -16,    13,    25,     1,   -25,    -2,    29,   -16,     3,    -1,    37,   -19,   -21,   -40,   -50,   -33,   -15,   -36,   -48,     9,     1,   -58,   -39,   -58,   -29,   -44,   -25,   -29,     4,    21,   -14,     3,     0,    12,   -12,     3,   -14,   -14,     7,   -10,    18,   -20,   -43,   -30,   -27,   -76,   -52,    -9,    -6,   -41,   -37,   -63,   -31,    -1,   -16,     0,     3,    58,    16,   -18,    15,    25,    25,    30,   -11,   -36,    23,    25,    11,   -41,   -51,   -48,   -65,   -76,    -9,    -4,    -8,   -26,   -60,   -60,   -22,   -27,    -9,   -27,     6,    22,    -5,   -13,    12,    -8,    34,    29,   -34,     3,    22,    51,    18,   -39,   -14,   -30,   -32,   -36,    -5,    -3,     2,   -15,   -11,    10,   -26,   -39,     5,    -8,    10,    -8,   -15,    -9,    -6,    -2,    49,   -26,    -4,   -21,    42,   -33,     7,    -2,    14,   -31,   -21,   -12,    15,    -9,     7,   -16,     2,    -2,    14,   -27,     1,    20,    27,   -25,   -28,   -13,    14,     2,    -7,   -22,   -42,   -70,   -24,   -38,   -31,   -23,    10,    10,     1,   -14,    -9,     9,     4,   -33,    -7,   -21,   -24,     5,   -21,    21,    -8,   -38,   -12,   -25,   -33,   -22,    -6,    23,   -48,   -56,   -44,   -32,    -6,   -14,    15,    -6,     3,     1,   -16,   -11,     7,   -33,    12,    24,     1,   -11,    -4,   -54,   -58,   -44,    -4,   -21,   -19,    -7,   -11,     1,   -49,     0,    -6,    10,     2,   -14,     2,    -5,    -7,     5,    -9,     5,   -38,   -42,    12,    38,   -18,   -51,   -44,   -53,   -31,   -55,     1,    -1,   -16,   -12,    -8,     0,   -33,    -6,    15,     1,   -22,   -33,     1,    -6,     9,     4,   -13,     1,    -9,    -6,   -17,     8,   -31,   -75,   -46,   -73,   -25,   -20,    16,   -25,   -27,   -37,   -59,   -24,   -44,   -22,   -19,   -25,   -25,    -8,    12,    10,   -23,   -10,     6,     2,     7,   -21,   -33,    -2,   -27,   -94,   -59,    -6,    -1,     1,   -17,     0,   -18,   -32,   -38,   -70,   -38,     5,     4,   -22,   -34,    20,    14,    17,   -56,   -16,     3,   -10,     9,     7,   -24,   -29,    -1,   -35,   -49,     5,     4,    14,    35,     7,   -17,   -50,   -19,   -36,   -21,    14,   -30,   -21,    -3,     9,     4,     9,     1,     3,    -9,    -7,    10,   -20,   -16,   -15,   -42,   -28,   -32,    12,   -16,    10,    -1,   -34,   -58,   -36,   -10,   -18,   -12,    42,    27,   -45,    -3,     7,    28,    17,     9,     5,     0,     7,     6,     1,   -11,   -43,   -22,    -6,   -10,    11,    14,    32,    14,   -46,    -5,   -10,    20,     0,   -19,    50,    45,    29,    16,    25,    20,    -6,    44,    -3,    10,    -1,     0,   -24,     5,   -37,    -9,   -44,   -23,   -43,   -36,     8,     6,    17,    12,     5,   -21,   -37,    -2,    37,    44,    13,     6,    36,    13,    16,    -6,    -9,     9,     2,     1,     4,    -8,   -34,    -7,   -24,   -29,   -30,   -41,     6,   -18,    16,   -13,   -50,   -21,    -6,   -21,   -50,   -24,   -25,   -76,   -70,    -3,   -14,     0,    -1,    -9,     8,    -4,    -3,     9,     5,    -1,   -16,    -5,    -3,   -15,   -61,   -60,   -43,   -37,   -47,    -6,   -26,   -53,   -17,   -35,   -26,   -21,   -16,   -12,    -9,     4,     7,    -4),
		    35 => (    9,    -3,     8,     6,     0,     2,    -5,     2,     3,     7,    -8,    -4,    -8,    -7,    10,    -2,    -1,     4,     4,     1,    -3,    -5,     1,     3,    -5,     8,     8,     3,    -5,     0,     5,    -4,     6,    -1,    -8,    -3,    -6,    -5,     4,   -16,   -13,   -10,    -9,   -19,   -31,   -27,   -10,   -21,    -4,   -13,    -9,    -7,    -1,    -3,    -9,    -5,     8,   -10,    -8,   -15,   -16,     8,   -26,   -23,   -21,   -43,   -49,   -40,   -55,   -51,  -119,   -80,   -47,   -25,   -18,    15,     3,   -55,   -23,    10,   -24,   -17,     2,     3,     8,     6,    -4,     4,    -9,   -50,   -40,   -33,   -78,   -85,   -65,   -17,   -20,    -5,   -17,   -20,   -35,    21,    55,    24,   -33,   -17,   -20,   -33,   -33,    -7,     5,    -8,    -2,     4,   -17,    14,   -31,   -16,   -52,     3,   -17,    -5,    28,   -17,   -53,   -18,    25,    34,   -11,   -25,     4,   -34,   -37,   -19,   -42,   -62,   -70,   -49,   -15,   -10,    -3,     0,   -10,   -10,   -33,     4,   -29,   -69,   -51,   -28,   -29,   -11,   -52,   -46,   -23,   -47,   -45,   -82,   -89,   -14,    17,   -37,   -38,   -11,   -47,   -61,    20,    12,    -4,    -3,    32,   -46,   -51,    24,   -27,   -39,   -12,   -37,    10,   -16,   -44,   -19,     3,   -24,   -40,   -32,   -14,   -11,    -4,    -7,     1,   -10,     0,   -57,    -9,     3,     6,   -13,    34,   -24,   -58,    23,   -54,   -24,   -10,    -8,    68,    15,   -21,    -3,    -4,    13,   -43,   -46,   -77,   -80,   -24,    -8,     7,     9,   -24,   -14,    -1,    37,    -8,    -2,   -40,     5,   -20,   -12,   -29,    -5,    -3,     6,    16,    23,   -17,   -16,    24,    20,    28,    22,    -2,    34,    34,    35,    51,    52,    48,    34,   -30,    24,    -2,    -4,   -43,   -30,   -21,   -71,    16,    24,    -6,    -8,   -11,   -37,   -20,    -7,    26,    23,    55,    88,    63,    72,    48,    58,    50,    36,    84,    68,   -49,     9,    -3,    -7,    -9,   -33,    -4,   -15,    19,    17,   -18,    -3,     4,    39,   -22,    -5,     9,    15,     8,    33,    73,    64,    63,    79,    54,    25,    92,    66,    33,    49,     9,   -11,    -4,    -9,    14,     1,   -19,   -45,   -17,   -31,    19,   -11,   -19,   -34,   -70,   -61,   -51,   -54,   -39,   -65,   -45,    12,     8,    32,    10,    77,    69,     4,     0,   -11,    -4,     9,   -15,   -26,   -34,   -11,    -2,    25,    33,    46,    24,     0,   -35,   -47,   -77,   -67,  -137,  -221,  -140,   -93,   -94,   -56,   -46,    46,    70,   -22,     0,    -1,   -11,    15,   -15,   -47,   -55,    21,     3,   -11,    57,    19,    35,     8,    11,    -1,   -39,    -2,   -49,   -93,  -124,   -78,  -107,  -110,   -39,   -16,    48,   -23,    17,     5,   -13,   -16,    24,    -4,    21,    14,    39,    36,    -3,     3,    -8,    -8,   -11,    -3,   -21,    16,    -1,   -75,   -83,   -63,   -54,   -38,   -40,   -51,   -15,   -10,    11,     2,   -40,    38,    66,    29,    12,    50,    32,    38,    -8,     5,    14,    -5,   -31,   -37,   -61,   -16,    23,    -2,   -34,   -31,   -59,   -26,   -42,    21,   -14,   -30,     1,     3,   -37,     6,    25,    69,    -9,    36,    -1,    22,    -2,   -24,   -20,    -9,   -58,   -23,   -34,   -15,    18,     0,    -4,   -28,   -23,   -32,   -20,    20,   -36,   -40,     7,    -8,   -69,    10,    18,    18,    12,   -27,   -15,    17,     8,   -11,   -45,   -45,   -41,    -4,   -21,    -4,   -28,    -2,   -23,   -41,   -14,   -13,   -68,   -74,   -71,   -70,   -17,   -11,   -38,   -73,   -34,   -22,     1,   -20,   -24,   -38,   -77,    31,    39,   -20,   -39,     9,   -31,     6,   -18,     3,    22,   -42,    -9,    36,     7,   -26,   -76,   -47,     2,     1,   -11,   -62,    28,    42,   -14,   -26,   -15,   -55,   -67,   -67,    -3,    27,   -44,   -35,   -15,    12,     9,    33,     4,   -48,    16,    63,    61,    71,   -66,   -53,    -2,     3,   -11,   -42,    33,    -1,   -30,    -7,   -29,   -27,   -36,     3,    14,    26,   -84,   -26,    10,    -1,     4,    26,    19,   -35,    12,    10,    72,    81,   -55,     0,    -1,     7,   -13,   -29,   -15,    21,   -35,   -37,   -11,    -5,     9,    11,    18,    12,   -24,    44,   -13,    -5,    -9,    -5,    12,   -24,   -40,     1,    56,    94,    46,    -9,     0,    -4,   -30,    -6,   -15,    22,    23,   -33,   -51,    -5,     6,    14,    36,    10,    -2,    29,    14,    28,    -1,   -35,     8,    -7,   -34,    65,   110,   109,   108,     9,    -8,    -3,    34,    -7,     0,     1,   -19,   -47,   -44,    28,    44,   -21,    -1,   -28,    11,    15,   -17,    -5,    -3,   -36,     3,   -32,    -5,   103,   109,    97,   126,    -7,     9,    -8,    -8,     1,   -50,   -70,   -52,   -34,   -20,   -27,     6,    16,    34,   -14,    34,   -12,   -11,   -15,   -25,   -21,     4,    29,    71,    37,    28,   -76,   -24,     7,     3,     5,    -4,     4,   -69,   -77,   -46,   -66,   -50,   -28,   -36,     7,    71,    37,    -8,   -43,   -30,   -26,    12,    -2,   -38,    31,    41,    53,    56,    -8,   -12,    -8,    -4,     0,    -4,     1,   -40,   -84,  -115,  -107,  -101,   -95,   -86,   -58,   -60,   -91,  -145,   -38,    -6,   -23,   -12,    11,    -2,    18,    -3,   -45,   -22,     6,     7,    -2,     5,     4,     8,     5,     1,   -19,    -9,   -23,   -21,   -12,    -7,   -19,   -22,   -16,   -79,   -41,   -17,   -32,   -44,   -29,   -19,   -34,   -74,   -53,    -7,     7,    -5,     0),
		    36 => (    1,     6,     2,     6,     0,    -3,     6,     1,    -8,    -7,    -6,    -3,    12,     6,     0,    -4,     6,    -8,    -4,     8,     6,     5,     5,    -5,    -6,     2,    -7,    -1,    -7,    -6,     6,   -10,     4,     7,    30,    33,    31,    23,    46,     7,    -2,    21,   -30,     2,     6,    20,    44,    28,    86,    35,    33,    32,    10,     4,    -3,     8,    -6,     2,    27,    16,    43,    38,    43,    54,    31,   -17,   -24,   -32,   -44,   -44,     6,    24,    37,    73,    40,    19,    14,    79,    73,    54,    36,    51,    -9,    -4,    -4,    -2,   -59,     9,   -20,    28,    53,    51,     2,   -24,   -27,   -76,  -101,    -3,    46,    30,   -38,   -25,    13,   -24,   -24,    -4,   -39,    12,   -59,   -30,   -46,    -7,     3,     5,   -80,   -10,    26,    65,    47,   -21,   -52,   -43,   -57,  -100,  -130,   -55,   -69,   -37,    -2,   -28,   -14,    86,    56,    12,   -67,   -76,  -121,   -89,   -34,    24,     1,     1,   -37,   -47,    23,    50,    23,   -17,   -24,   -22,   -35,  -110,   -76,     3,    11,   -37,   -21,    -1,    24,    25,    45,    31,   -24,     3,   -57,   -85,     4,     7,    -9,    -6,    37,    13,    13,    48,    46,    -5,   -15,   -57,   -62,   -44,   -28,   -37,   -30,    44,    31,    10,     4,    -6,     3,     4,    17,   -32,   -26,   -68,   -33,    -9,     0,    -5,    -5,   -17,   -16,     7,   -22,     2,   -37,   -68,  -116,   -86,   -29,   -34,    19,    30,   -32,   -45,   -15,   -80,     7,   -10,    35,   -44,   -99,   -93,   -19,   -38,     2,     1,   -40,   -31,   -18,     8,    31,   -36,   -57,  -110,  -109,   -18,    -4,    -9,   -13,    13,    -1,   -37,   -94,    -1,   -34,   -42,   -40,  -107,   -92,   -42,   -36,   -50,     3,     0,   -36,   -26,    55,   -16,    -8,    -7,   -60,   -56,   -30,    -5,   -16,    11,    32,    16,   -42,   -71,   -97,  -121,  -148,  -139,  -130,  -119,   -93,   -51,   -55,   -17,     8,     5,   -34,   -17,   -35,   -39,   -47,   -45,   -95,   -26,    12,    -1,    10,    16,     2,    -9,   -40,   -14,   -19,   -84,   -86,   -83,  -105,  -118,   -83,   -68,   -49,   -38,    -4,     2,     9,   -59,   -25,    -9,   -13,   -23,    11,     1,    12,    15,    27,    25,   -11,   -58,   -51,   -22,   -39,   -13,   -23,   -42,     0,  -101,  -104,   -95,   -62,   -53,     9,    -8,   -12,   -41,   -38,   -13,    -7,   -40,    -5,    10,    36,    27,    14,    61,   -21,     7,   -43,    27,    -9,    -1,   -18,   -35,    16,    12,   -42,   -96,   -97,   -49,    -7,     4,   -12,   -50,   -40,   -21,   -38,   -49,    10,     7,    18,    65,    15,    33,     2,     6,   -14,    19,    66,     0,    10,     3,    66,    56,   -56,  -110,   -53,    -2,    -4,     5,    -5,   -61,   -42,    10,   -55,     1,   -19,    24,    37,    12,     1,   -23,   -18,    -3,     2,   -83,    17,    31,    -4,    57,    41,     4,    15,   -39,   -49,     1,     3,    10,     2,   -52,    -6,    13,   -32,    -1,    24,    21,    23,   -44,   -16,   -19,    -1,   -58,   -48,   -60,    16,    44,    22,    69,    26,    11,   -51,   -72,   -87,   -50,     0,     6,     0,   -20,   -16,    21,    -7,    37,   -11,    26,     4,    26,    44,    33,    27,     1,    15,    -1,     3,    -7,    29,    61,    34,    -6,   -68,   -79,   -82,   -65,     1,    -4,    -5,     3,    11,    19,     5,    12,    46,    -3,    16,    26,   -25,     3,   -15,   -26,   -25,    -9,    -3,     2,    24,    54,   -18,   -16,   -63,   -53,     0,   -67,    -2,   -10,     5,     1,    48,   -13,   -30,   -14,   -11,    49,    30,   -26,   -15,   -22,    -5,    53,    -9,    23,    36,    21,    13,   -11,   -97,   -75,   -57,   -48,   -10,   -28,     1,   -22,   -28,    11,    34,   -35,   -14,     0,   -29,    12,    23,    41,    -3,   -77,   -27,    20,    -7,    -9,    32,   -21,   -17,   -37,  -103,   -41,   -21,   -21,   -35,   -11,    -7,   -25,   -20,   -62,    41,    16,   -14,   -13,   -11,   -25,    11,    39,    38,   -21,    -7,   -13,   -56,   -38,   -55,   -15,    -3,    -6,   -15,   -50,   -27,   -32,   -43,     7,     4,    -7,   -31,   -30,   -28,   -37,    -1,   -11,    -6,     0,   -17,    42,   -20,   -10,   -22,   -51,   -18,   -30,   -20,   -36,   -13,     7,   -41,   -34,   -33,   -34,   -32,    -8,    -7,    -3,   -11,   -22,   -41,   -56,   -62,   -31,   -38,   -20,     3,     7,    20,    29,    -3,    12,   -18,   -44,   -20,   -37,   -67,   -58,   -15,   -38,   -77,   -35,     8,   -10,    -1,     6,     7,   -11,   -24,   -35,   -40,   -66,   -45,   -58,     0,    26,    20,    -5,    19,    33,   -39,   -77,    40,    59,    36,    -6,    -6,   -13,   -16,    -9,   -17,    -9,    -9,    -8,     5,     8,   -17,    -5,    -7,   -25,   -42,   -63,   -72,   -73,   -34,   -15,    14,    48,    60,     1,    -7,   -75,   -46,   -14,   -17,    -1,    -4,    -5,    10,     9,     5,    -2,    10,    10,     9,    -7,   -22,   -32,   -21,    -9,   -32,    18,    42,     8,    -7,     0,   -11,    -9,    -1,   -14,   -32,    -9,     5,     1,   -10,     9,    -5,     9,     4,     1,    -9,    -9,     0,     1,     4,    -1,    -1,    -2,    -5,    -5,     6,    -8,    -1,   -13,   -14,     2,     2,     7,    -1,   -15,     0,   -11,     1,    -6,     8,     2,     5,    -5,     8,     1,     2,     3,     9,    -8,     4,     6,   -11,    -2,   -10,     1,   -11,     0,     3,   -11,   -12,     5,     3,     2,     6,     1,    10,     1,     8,     0),
		    37 => (    0,    -8,    -2,     5,     3,     4,     5,     2,    -1,     2,    -2,    -9,     0,    -5,     9,     1,     2,    -3,    -5,    -7,     4,     4,    -8,     3,     5,     8,   -10,    -9,     1,    -9,     3,     5,    -3,     1,     5,    -6,    -6,   -11,    -4,   -34,   -42,   -27,   -20,   -33,   -39,   -32,   -11,     3,    -3,    -2,     9,    -6,     4,     8,   -10,     4,    -8,     4,    -2,   -25,   -25,     1,    -8,   -28,   -49,   -19,    -5,   -42,   -18,    -4,     1,    -4,    -1,   -13,   -12,     6,    -3,     2,     3,    -8,     6,     0,     7,     3,    -9,     9,    -9,   -18,   -15,   -10,   -27,   -72,   -69,   -22,   -39,   -33,   -25,   -30,   -15,   -19,   -20,   -49,   -21,   -34,   -11,   -12,   -17,    -2,    -7,     4,   -10,    -3,    -8,    -2,     7,   -12,   -47,   -37,   -27,   -42,   -77,   -73,   -73,   -84,   -83,   -41,   -73,   -59,   -40,   -38,   -42,   -14,   -23,   -28,   -34,   -33,   -34,   -14,     3,     8,    -5,     8,     6,   -58,   -93,    14,   -29,    26,    84,    27,   -52,   -75,   -43,    31,   -25,   -14,   -90,  -107,   -75,  -112,   -92,   -48,   -48,   -49,   -14,   -44,    -6,    -7,     4,     3,    15,    17,    -9,     3,    -6,   -39,    -1,   -16,   -66,   -38,   -44,   -53,   -21,   -38,   -86,    -8,    23,    -7,     1,    51,     5,   -44,   -68,    -8,   -71,   -22,     4,    13,    13,    29,    26,    10,    24,    34,     5,     0,     8,   -51,   -29,   -16,   -26,   -61,   -50,    -9,     0,   -98,   -57,   -15,   -13,   -28,   -62,   -30,   -31,   -17,   -23,    13,   -35,     8,    31,    39,    64,    23,     7,    55,    -6,     9,    22,     5,   -46,   -27,   -28,   -24,    26,   -47,   -19,     2,   -21,    10,     1,   -31,   -56,   -17,     4,    18,     1,    14,    86,     1,    12,    -3,    -9,    10,   -40,    20,    54,    28,    41,    26,   -32,   -30,    -6,   -19,     6,    42,    34,    72,    13,   -45,   -34,    40,     1,    49,    27,    34,    91,    40,    41,   -34,     4,    29,    -1,    33,     8,    -1,    33,    40,    -8,    -2,   -11,    -2,   -15,   -14,    79,    30,   -57,    -6,   -29,    41,    -6,    30,    77,    65,    80,    13,   -29,    -6,   -24,    -3,    12,    30,    -4,    11,    13,    17,   -33,   -25,   -19,     6,   -39,    25,    25,   -23,   -89,   -75,   -18,    63,     8,    11,    10,    88,    38,    16,   -12,   -13,   -17,   -15,   -11,     8,     7,   -18,    15,    16,     8,   -30,    22,    13,    -8,    33,    44,   -51,   -46,    20,   -18,    48,    10,    32,    37,    80,    32,    21,   -28,   -23,   -45,   -34,    26,    21,   -12,   -56,    19,   -39,     4,   -14,   -17,   -21,    67,    44,    16,   -13,    -6,    52,   -25,   -24,   -13,    19,    82,    82,    -8,    34,   -25,   -45,   -32,    -7,    34,    27,   -37,  -101,   -18,   -21,    -2,    28,     1,    46,    34,    36,    21,    70,    69,   -30,   -37,   -11,    -5,     8,    48,    41,   -34,     5,    12,     1,   -18,     5,    39,     1,   -53,   -62,    -5,   -37,   -36,    12,    11,    70,    26,    12,    43,    31,    25,   -48,   -22,   -17,     1,     1,    20,    13,    57,    20,   -23,    22,    21,    56,     5,   -13,   -98,   -45,   -32,     3,   -15,     5,     7,    28,     2,    59,    84,    75,    32,  -120,   -51,     4,   -10,    -3,   -20,    -5,    33,    16,   -31,     3,    26,    23,   -37,   -52,   -82,   -72,    24,    18,    10,   -14,    -8,   -14,    21,    32,    83,    40,     0,  -115,   -33,   -75,    35,     7,    27,   -88,    -1,     6,   -29,    17,    26,    10,   -32,   -70,  -157,   -59,    45,    32,     8,    -1,    -7,   -34,    10,    23,    43,   -10,   -61,   -28,    -4,   -25,     2,    32,   -10,   -79,   -18,     9,    35,    11,     4,   -15,   -95,  -175,  -145,   -46,    54,     2,   -25,    11,   -34,   -17,   -27,   -75,  -113,   -56,   -45,   -50,    -3,    -4,    -4,    21,    -7,   -17,    17,    52,    39,    39,     5,   -94,  -132,  -180,   -49,   -20,     4,     2,   -11,   -23,   -32,   -39,   -48,   -56,   -82,   -76,    -9,   -39,     3,     5,    -1,    -8,    -9,   -18,   -42,    32,    11,    15,   -49,   -92,  -111,   -90,     0,   -40,    11,    24,    33,   -30,   -33,   -35,   -52,   -27,   -42,   -70,   -71,   -25,    -7,     2,    -1,     3,    -7,   -12,     0,    -3,    11,   -21,   -62,   -58,   -94,   -47,   -14,   -21,    20,     0,     0,     5,     9,    14,    14,   -24,   -38,   -45,   -32,   -28,   -44,     6,    -9,     3,   -20,   -19,    12,    16,   -10,   -26,   -62,   -56,   -82,   -48,    11,   -10,    41,    21,    -5,     5,    50,     2,    -5,   -36,   -42,   -63,    -2,   -19,   -32,    -8,    -6,     7,   -13,    -2,     7,    -7,    -4,   -29,   -50,   -54,   -70,   -33,    12,   -24,    -1,   -12,   -12,    17,     8,    30,    -4,    -7,   -16,   -66,    -2,    -1,    -9,     9,    -2,     5,   -18,    -1,    -4,   -10,     6,   -11,   -39,   -45,   -85,   -42,   -48,   -28,    30,   -10,    37,    35,    26,    37,    10,     8,    17,   -80,    -5,   -24,     5,    -7,     5,    -1,   -10,     1,     2,   -11,    -3,    11,    19,    12,   -16,   -84,   -54,   -27,   -77,   -31,    29,    22,    29,    56,     8,    16,    17,   -17,   -18,     9,    -1,    -6,    -2,   -10,    -9,     5,     5,    26,   -32,   -30,     4,    41,    35,    -1,   -12,   -51,   -63,   -28,    34,    40,     9,   -44,     7,    48,    30,    41,     7,     6,    -5,     2),
		    38 => (   -3,     0,     1,     4,     8,     7,     6,     1,    -3,    -7,    -3,     2,     4,     3,     1,    -4,     3,     9,    -9,     0,    -7,    -4,    -7,     3,    -3,     7,     7,     6,    -7,     8,     1,     9,    -8,     7,    -6,    10,    -8,     5,     4,    -8,     8,   -11,   -18,   -38,   -45,   -23,   -20,    -1,   -17,    -6,   -15,    -9,    -7,    -4,    -9,     5,     2,     4,   -15,    -5,     0,   -10,    -2,     2,   -17,   -20,   -39,   -33,     4,   -10,     2,   -23,   -13,   -25,   -12,    -7,   -34,   -38,   -47,   -22,    -6,   -17,    -2,    -5,     6,     5,   -16,    -5,    -4,   -35,   -14,   -50,   -49,     5,    -5,   -33,   -31,   -36,     4,    32,    33,    26,    10,   -18,   -23,   -12,    -5,     7,    -7,    -4,   -26,    -6,    -7,    -9,    10,   -20,   -57,   -25,    -5,    -3,     5,    -8,   -16,    -8,   -25,   -34,   -10,    13,    18,     6,    11,    10,    39,    28,   -30,   -15,   -58,   -26,    -9,   -22,   -10,    -3,   -14,   -48,   -56,   -19,    -4,   -17,   -29,   -38,   -34,   -40,   -44,   -44,   -34,    17,   -12,   -10,    20,    26,    30,     4,    -3,   -38,   -21,     0,     2,   -31,    -3,     3,   -21,   -27,    -3,    12,   -24,   -13,   -19,   -41,   -61,   -63,   -50,   -32,     6,    11,     1,    -1,   -14,    28,   -20,    31,     8,     2,   -37,    -8,    -7,    -2,     7,   -36,   -26,   -17,    11,    -5,    -4,     4,    15,    -7,    11,   -14,   -13,    27,     8,    19,    -5,   -30,   -19,    -5,    -4,   -30,    -2,   -12,   -26,    22,    37,    14,   -15,   -23,   -14,     5,     4,     7,     4,     9,   -14,    24,    23,     0,     4,    -5,    56,    50,    12,     5,   -26,     2,   -28,   -15,   -32,    -9,    39,    72,    51,    22,     8,   -20,    -6,     8,   -12,   -18,   -19,   -10,   -42,   -40,    -6,   -28,   -12,    -3,    19,    37,     6,   -35,   -41,     2,   -24,    -7,    10,    45,    47,    46,    18,   -66,     4,   -10,     0,    -3,   -18,   -24,   -28,   -24,   -24,    12,   -25,   -51,   -42,   -26,     6,    -9,   -13,   -21,   -52,   -27,    -7,    47,    42,    17,     0,   -67,   -36,   -61,    -1,    -4,   -10,    -5,   -15,   -23,   -33,   -20,   -37,    -9,   -10,   -46,   -23,   -25,    19,   -16,    12,   -30,   -10,    12,   -31,    -8,    46,     1,   -20,   -38,    21,   -40,     6,     5,    -5,   -31,   -13,   -31,   -22,   -45,   -59,    -6,     9,    -2,    10,     7,    -9,    21,   -13,    11,    20,     7,    31,    23,    -2,     0,    -3,   -56,   -32,   -63,     2,    -8,   -31,   -53,   -14,   -19,   -62,   -48,   -32,   -24,   -35,   -11,   -21,    13,     4,     6,    20,    37,   -18,   -13,   -37,   -33,     8,    -4,     3,   -28,    -9,    14,    -5,    -4,    -9,   -64,   -24,   -39,    32,    20,   -29,   -81,   -64,     8,    -3,    32,    22,    11,    26,   -31,   -34,   -70,   -20,     7,     4,    11,     0,     5,   -17,   -22,   -10,    -9,    -1,    -8,   -17,    -7,    58,    22,   -36,   -36,   -11,    19,    26,    19,     2,   -10,    -7,   -43,   -80,   -38,   -25,    -9,     4,   -34,   -40,     3,   -31,   -19,     6,    -4,   -13,   -18,   -13,    20,    29,     7,    17,    41,    25,    33,    14,   -34,   -55,   -41,    -4,   -58,   -88,   -56,   -38,   -14,   -27,   -47,   -37,    -1,   -59,   -28,     7,   -15,    -3,   -14,    -4,    18,    50,    84,    64,    48,    31,     0,   -43,   -27,   -40,   -27,   -50,    -7,   -43,   -31,   -31,   -58,   -33,   -36,   -22,   -12,     5,   -12,     5,    -7,     2,    -7,    -6,    30,    54,    49,    45,    26,   -25,   -44,   -69,     2,    34,   -33,   -44,    -7,     5,   -11,   -34,   -52,   -50,   -18,    -9,   -18,     0,   -29,    -1,     3,    -8,   -37,    15,    62,    29,   -11,     8,   -31,   -72,   -41,   -24,    14,     3,   -11,   -32,     6,    15,   -46,   -27,   -52,   -42,   -27,    -8,     0,   -27,   -20,    -5,    -8,    -5,   -41,   -15,    55,   -12,    17,    11,   -41,   -50,   -38,   -45,   -22,   -23,   -17,   -22,   -21,   -24,   -49,   -58,   -47,   -45,   -11,   -15,    -5,   -27,    -4,   -26,   -21,   -16,   -35,    -5,    44,     6,     6,    25,   -31,   -14,     7,   -35,   -31,   -27,   -45,   -37,   -26,   -55,   -70,   -67,   -56,   -18,   -12,    -4,     1,   -28,    -3,   -26,   -19,    -8,   -23,    10,    -6,     5,    10,    29,   -17,    -7,     5,   -42,   -38,   -20,   -49,   -10,   -34,   -45,   -36,   -57,   -47,   -22,   -12,   -19,    -6,   -27,    -6,     2,     2,     4,   -34,   -16,   -30,   -35,    11,     1,    20,     8,    -2,   -19,    -8,   -28,     1,    11,   -29,   -65,   -46,   -51,   -31,    -4,   -12,    -9,   -13,   -48,     0,     0,     3,   -13,   -11,   -38,   -14,    33,    49,    42,    60,    23,    12,    12,    -9,   -38,     6,   -25,   -33,   -34,   -26,   -14,     0,    -1,     2,   -21,   -16,   -15,     0,     2,     1,   -14,   -11,   -19,   -41,    -5,    28,    23,     7,   -11,     3,    19,   -15,    26,     6,   -13,   -23,   -14,     2,     3,     4,     6,    -3,     0,   -10,   -24,     3,     0,    -1,     3,   -39,    -9,   -33,   -42,   -40,    12,     4,     9,     0,    10,   -18,   -27,   -30,    -6,   -13,    -6,    -6,   -40,   -19,   -26,     4,     2,    10,     9,   -10,    -8,    -5,    -4,    -6,     0,   -19,    -9,   -10,   -10,    -7,    -4,    -4,     2,   -16,    -1,    -7,    -4,    -7,   -11,     3,     5,    -2,    -6,     8,    -7,     7,    -4,     3),
		    39 => (   -5,    -3,     2,    -1,     6,    -7,    -2,    -6,     3,     0,    -6,     6,   -10,    -2,     3,    -9,   -10,    -6,    -6,    -8,    -4,     8,     2,    -8,     0,    -5,    -3,     3,   -10,     8,    -8,   -10,    -5,     4,    -4,    -8,    -6,     5,    -9,    -3,   -37,   -33,    -2,   -19,   -20,   -16,   -31,   -15,    -2,   -11,    -7,    -5,    -7,     1,     9,    -5,     8,     2,     8,    -9,     6,     6,     1,    -6,   -13,   -28,   -24,   -24,   -10,     5,   -27,     2,    -2,    -6,     2,     5,   -10,   -16,   -25,     2,    -5,     7,     2,    -2,    -7,     1,     3,   -21,   -16,    -7,   -12,   -19,   -44,   -63,   -37,   -64,   -29,   -39,   -24,   -35,   -20,   -14,   -18,   -16,   -50,   -38,   -14,     2,   -23,   -13,     6,    -7,    10,     7,    -1,   -16,   -35,   -48,   -88,   -14,   -38,   -38,     0,   -12,   -26,   -48,   -59,   -74,   -36,   -38,   -12,   -19,   -23,    -8,   -10,    -3,   -10,   -62,    -8,     3,     7,     6,     7,    -9,    -1,    -6,   -30,   -33,   -54,    10,    33,     3,    -6,    24,   -36,   -59,   -30,   -49,   -92,   -40,   -34,   -51,   -11,   -19,    -8,   -22,   -15,     1,    -7,     5,    -3,   -34,   -40,   -76,    10,   -25,    30,    32,    46,    15,     6,    60,     5,   -41,   -65,   -45,   -84,   -33,   -80,   -32,    22,     8,   -46,   -11,    -5,    -9,    10,   -14,   -43,   -38,   -58,   -66,   -47,   -26,     6,    49,    20,     7,     2,    16,   -16,   -66,   -23,   -64,   -28,   -52,   -90,   -33,    15,    -2,   -28,   -21,   -23,   -12,   -22,   -17,   -42,   -39,   -43,   -33,   -42,   -26,    -7,   -20,    -9,   -33,     6,    21,    32,   -21,   -50,   -28,   -55,   -26,   -44,   -50,     4,    -2,   -18,   -26,    -9,     0,    -1,   -10,   -55,   -14,    -6,   -18,    14,    47,    21,   -27,   -41,    20,     7,    25,    19,   -15,   -26,   -15,   -30,   -56,   -33,   -62,   -36,   -37,   -51,   -47,   -13,    -9,     1,   -25,   -40,     2,    51,   -21,    32,     0,    20,   -31,    -8,    -8,   -19,   -12,   -27,    15,     7,   -17,    -8,   -51,   -38,   -14,   -93,   -99,   -52,   -37,    -2,   -28,    -2,   -56,   -23,    34,   -12,    -7,    67,    42,   -27,   -54,   -27,   -42,   -17,    15,    16,    33,    13,    37,   -27,     5,   -17,   -34,   -77,   -58,   -44,   -85,    -6,   -33,    -7,   -51,   -30,    21,    -9,    40,    46,   -24,   -26,   -11,   -35,   -67,   -23,   -12,    28,    23,   -10,    25,     4,   -20,    -5,    20,   -39,   -30,    -7,   -58,   -45,   -21,    -8,   -49,   -22,    -2,   -34,    47,     0,    -7,     5,   -10,    19,   -47,   -25,   -13,     6,   -33,   -17,    -3,    21,    -7,    25,    19,    -7,   -43,     2,   -42,   -25,   -13,   -16,   -12,   -14,    48,     2,    17,     8,    -6,   -10,    37,    40,    45,     8,    17,   -23,   -68,   -39,    10,    39,    -7,   -21,    23,    11,    -8,    20,   -60,   -25,     3,    -7,    -4,   -14,    43,    22,    30,    28,   -35,    14,    13,    -7,    19,    42,   -41,   -13,   -49,   -73,   -20,    22,    14,    15,    -9,   -10,    -2,    16,   -62,   -38,   -26,    -6,   -10,   -35,    12,    56,   -40,    26,   -13,    -7,   -18,   -14,   -12,     8,   -19,   -57,   -68,   -47,     5,    50,    43,   -14,   -13,   -41,    -6,    26,    -1,   -31,   -55,     9,    -7,   -32,     7,    14,   -22,     7,   -30,     1,   -17,    -7,     3,    19,    21,   -24,   -30,   -12,    19,    -2,    41,   -13,   -21,   -69,   -20,   -23,   -47,   -41,   -47,    -7,     4,   -34,    12,   -24,    25,    24,    15,   -22,    -1,    21,    35,    -6,    -5,    32,    39,    28,   -29,     8,    21,    21,   -68,   -44,   -28,   -21,   -45,   -54,   -36,     5,    -5,   -28,    -3,   -25,   -17,    13,    29,    -5,    29,    23,    24,    56,    30,     7,    -2,    -1,   -57,   -40,    12,    11,   -21,   -20,    13,     4,   -62,   -38,   -16,    -9,   -18,   -15,    -7,    12,    -7,   -49,   -53,    13,   -31,     3,   -35,   -45,   -36,   -34,   -59,   -56,   -59,   -17,    49,    11,   -15,   -20,    15,    74,     5,   -65,     0,     7,    -6,   -33,    -8,     7,    -7,   -13,   -55,   -94,   -96,   -37,   -27,   -50,   -48,   -70,   -70,   -88,   -49,   -28,    36,     6,     1,   -23,     5,    44,   -33,   -82,    -2,   -10,     1,   -37,    23,   -10,   -16,   -18,   -26,   -59,   -75,   -23,    30,   -11,    25,   -10,   -47,   -21,   -46,    -4,    10,    21,    -7,     9,     3,    31,   -56,   -38,    -9,     5,    -9,    -3,    38,    11,     7,   -17,   -24,   -36,   -38,   -26,   -28,     3,    17,     4,   -10,   -35,   -25,   -12,   -21,    18,     7,   -11,    51,    61,   -44,   -30,    -2,     6,     3,   -30,    -3,    -9,     3,   -16,   -21,   -27,   -53,   -35,   -41,     2,     0,     3,   -27,   -14,    -3,    20,    42,    75,    15,    56,    89,    18,    20,     1,    -9,     2,    -3,    30,   -17,   -21,    13,    -8,   -28,   -37,   -33,    -9,    10,    -3,    13,   -56,   -67,   -69,   -55,   -12,    45,    26,    19,    -5,   -33,   -27,     4,   -14,     6,     3,    10,     7,    20,    -3,     4,    22,    10,    12,     4,     0,   -24,   -16,    18,    17,   -18,   -49,   -41,   -50,   -44,     3,     5,    22,    46,    32,    -6,    -2,     4,     1,    -8,    -9,    -6,   -12,   -19,    10,    -3,     5,    -5,    -7,    -3,    17,    20,    21,    -2,   -26,   -28,    22,    15,   -25,   -53,    -4,   -28,     6,     6,    -1,    -6),
		    40 => (  -10,    -1,     1,    -8,    -7,     4,     3,    -3,    -9,    -3,     6,    -6,     9,    -2,    -5,    -2,     0,     7,    -7,     2,    -5,     0,     3,     9,     5,     4,    -3,    -1,    -5,     1,     4,    -2,     4,     5,    10,    -2,    -2,    -8,   -16,     7,    21,    -3,    -6,    14,    27,    29,    -1,     1,     9,     5,    -2,     9,   -10,    -6,    -4,     0,    -4,     1,    10,    26,    19,    -4,     2,     6,   -28,   -57,   -48,   -31,   -51,   -77,   -61,   -77,   -17,   -35,   -31,   -48,   -47,   -10,   -43,   -24,   -16,    -7,    -4,     5,     4,    -7,    -9,    16,     2,   -15,   -35,   -14,   -20,    -1,    -7,   -26,   -22,     0,     0,   -12,   -21,   -39,   -70,   -82,   -18,   -22,   -48,   -38,   -28,   -11,   -35,     1,     9,    -1,    -6,   -16,    -4,   -59,   -50,   -24,   -17,    29,    -5,   -21,   -52,    -4,     0,   -15,    14,   -37,   -46,   -27,   -33,   -23,    20,   -47,   -26,   -29,   -46,     0,    -1,     6,   -22,    23,    -6,   -26,    -8,     3,    30,   -22,    -7,   -28,   -28,    17,    -8,   -28,   -11,    14,    -3,   -36,   -52,   -37,    -9,   -33,   -20,   -26,   -39,   -35,     7,     3,   -15,   -17,    34,    27,    10,     6,   -59,   -52,    -4,   -20,   -24,    22,   -18,   -33,    10,    16,   -35,    26,    -6,    33,    12,   -63,   -32,   -69,   -36,   -19,     7,    -2,   -16,   -21,    34,    33,     8,   -24,   -72,     9,   -12,   -28,     0,   -16,    -5,     2,    14,    35,    58,    55,    13,    16,    10,    24,   -46,   -26,   -72,    25,    59,   -32,    40,     3,    24,    18,   -17,     5,    -5,    -1,   -15,   -18,    50,     0,    24,    16,    26,    31,    45,   -34,     3,    24,    12,    36,   -61,   -82,   -66,   -11,    -4,   -11,    45,    -3,   -57,    -5,   -11,   -22,    14,     4,   -31,   -28,     2,   -19,    22,    -3,   -36,    12,    24,   -14,    57,   -19,    -3,    -9,     5,   -86,   -74,     0,    -3,    -5,    44,     0,   -36,   -45,     1,   -23,    -7,    -9,   -34,   -52,     7,     2,    32,    -2,   -11,    14,    -4,   -22,    46,    28,    51,   -11,     0,   -57,   -69,     1,    -9,    93,   -32,    -9,   -42,   -52,    35,    48,    13,    19,   -12,   -10,    10,   -12,    11,   -26,   -30,    11,   -38,   -15,    26,    44,    35,   -34,   -35,   -58,   -57,    -5,     7,    13,   -12,   -14,   -40,   -35,    56,    39,    20,    22,    -4,    12,     6,   -24,   -40,   -34,   -70,   -46,   -15,   -14,    20,    48,    14,     7,    -6,   -15,   -62,     4,     2,    18,    22,    30,   -17,    16,    40,    42,    67,    27,   -11,    11,   -52,   -44,   -18,   -82,   -57,   -67,    19,     5,    11,    34,    42,    31,     8,    34,   -33,   -11,    -3,     9,    -7,    12,    11,    62,    49,    88,    52,    21,     3,    11,   -19,    -7,   -44,   -52,   -79,   -36,   -11,    29,    19,     1,     4,    48,   -12,    -7,   -50,     7,    -4,     3,   -19,   -24,    -5,    40,     2,    35,    77,    32,    -6,    -5,   -21,   -31,   -50,   -54,   -24,   -56,   -11,     1,    28,    49,    37,    69,    49,    10,   -78,   -20,    -4,    -7,   -17,   -35,    33,    -4,    41,    59,    22,    15,    19,   -25,   -43,   -42,   -60,   -52,    -4,   -13,    15,   -36,   -19,    44,    29,     0,    25,   -28,   -87,    55,    -6,    -7,   -25,   -60,    13,   -25,    -6,     6,    34,    43,    -3,   -47,   -77,   -53,   -18,    27,    -3,   -14,   -37,   -30,    14,   -37,    52,   -18,    16,   -43,   -64,    61,     9,     7,   -18,   -61,   -16,   -49,   -12,    34,    80,    47,    15,   -38,   -76,   -39,    27,    12,    -1,   -14,     1,    -6,    16,     3,    29,   -32,    -5,    -3,   -38,   -26,     5,    27,   -28,   -24,   -15,   -36,   -26,   -14,    71,    28,    17,   -57,   -26,   -35,   -29,   -14,     5,   -25,    -8,   -39,    51,   -10,    23,    -8,    -5,   -74,    -7,    -6,    -3,    21,   -47,     3,   -11,     8,   -16,   -10,    28,    44,    83,   -31,    -2,   -23,   -17,   -36,   -27,   -22,   -32,   -15,   -45,   -32,   -19,   -60,   -54,   -39,    21,     7,    -2,    -9,   -65,   -29,   -15,     0,   -30,   -33,    15,   -13,    -3,   -27,   -33,   -43,   -32,    -1,    18,   -22,   -62,   -44,   -34,   -21,    37,   -19,   -33,   -30,    32,    15,     3,    -8,   -62,   -15,   -58,   -11,     5,     7,    43,    35,    27,   -33,   -14,   -13,   -17,    -7,   -41,   -52,   -40,    -5,   -32,     8,    12,   -20,   -22,     6,    32,    21,    -1,     9,    -6,   -71,   -54,   -37,     4,     5,    -5,    17,    22,    29,   -20,     1,   -21,   -21,   -27,   -32,   -64,   -33,   -62,   -16,   -40,   -37,   -43,   -14,   -30,    -5,    -9,    -9,   -10,     6,     6,    27,   -34,   -40,    -8,    40,    28,    29,    31,   -26,    -9,    14,   -36,   -63,   -41,   -43,   -37,   -43,   -55,   -45,    -9,    17,     0,    -5,    -8,     9,   -10,    -6,   -53,   -79,   -69,   -55,   -55,   -50,   -74,   -73,   -88,   -42,   -38,   -99,  -100,   -90,  -110,   -74,   -59,   -45,   -42,   -22,   -14,     4,    -2,     2,     3,     7,    -4,    -2,   -21,   -30,   -74,   -37,   -36,   -62,   -70,   -80,   -54,   -51,   -44,   -56,   -41,   -77,   -75,   -49,   -63,   -54,   -24,   -31,     1,    -3,     4,    -9,    -7,    -4,    -4,    -5,     8,    -8,    -9,     7,     2,    -4,     1,     4,    -8,   -34,   -14,   -19,   -19,   -16,    -8,     4,     2,   -31,   -21,   -19,    -3,     2,     5,     3),
		    41 => (    9,    -3,     2,     9,    -9,     0,    -6,    -2,   -10,     3,     3,     4,    -2,     2,     0,     9,    -3,     8,    -6,    -5,    -8,    10,     8,     5,   -10,    -3,    -4,    -9,    -1,    -7,    -2,    -4,     8,    -6,    -5,    -8,     7,    -1,   -11,   -10,   -21,   -25,     9,    23,     1,   -19,    -6,     6,     6,     2,     6,    -6,    -5,    -9,    -8,     0,     0,    -9,     8,    -8,    -1,    -7,     3,    -1,   -15,   -19,   -28,   -20,   -22,    51,    65,    86,    74,    43,    44,    86,    62,   -54,   -59,   -40,     5,     7,     0,     7,     8,    -6,    32,    60,    -5,   -29,   -45,    38,    26,   -10,   -82,   -81,     4,     7,    12,    35,    74,    34,    32,    40,    63,    57,   -32,   -39,   -19,   -15,     9,     9,    10,     4,     6,    38,     3,    13,   -17,   -48,   -38,   -21,    10,   -22,   -54,   -63,    11,    55,    55,    23,    41,    13,    15,    35,   -33,   -27,   -16,   -44,   -40,   -33,   -10,    -1,    28,    23,     6,    47,    18,   -52,   -36,   -39,   -18,   -20,   -59,   -30,    -9,    31,    53,    14,    -2,   -21,   -21,    32,   -34,    -8,   -18,   -37,   -35,   -19,    -6,    -4,   -40,     4,     4,    14,   -37,   -46,   -25,   -28,   -42,   -42,   -17,    10,     9,    32,    46,   -11,   -11,   -29,   -10,   -23,   -23,     3,     6,     0,   -28,   -22,    -7,   -13,   -53,   -14,   -26,   -66,   -73,   -10,    27,    23,   -23,     6,     4,   -23,    45,    11,     7,    12,   -86,   -49,    -9,   -32,   -43,   -16,    -3,    -3,   -35,   -36,    -9,   -18,   -51,     1,   -27,   -73,   -37,   -31,    13,    94,    -8,   -25,   -18,   -16,    18,    28,    -6,   -21,   -12,   -47,    -5,   -27,   -26,   -19,   -15,    -9,   -34,   -19,    -2,     0,   -58,   -13,   -26,   -40,    -3,    13,    44,    31,    13,   -32,   -33,   -14,    19,    32,    26,   -71,   -30,   -75,   -38,   -42,   -18,   -25,   -15,   -17,   -12,   -25,    10,    -2,   -61,    -8,   -42,   -64,   -36,    35,   -30,   -32,   -17,    -6,     1,   -27,     0,    -6,     0,     0,   -33,   -33,   -35,   -41,   -15,    -9,    -9,   -17,   -25,    30,    -2,    13,     5,    -7,   -24,   -34,     2,   -20,   -58,     9,    40,    -5,    -2,   -46,     1,    -6,   -11,   -34,   -74,   -39,   -42,   -20,   -28,    -5,   -26,   -13,   -38,     7,    -4,     7,    -4,    -8,    -5,   -17,   -19,   -34,   -42,    31,     0,    37,   -26,   -75,    -5,     2,    10,   -58,   -30,   -60,   -36,   -11,   -19,    -5,    -4,    -8,     5,     7,    -4,     5,     7,     0,   -32,   -17,   -16,   -34,   -13,    45,    10,    -6,   -18,  -129,     5,    21,     3,   -27,   -94,   -58,   -34,   -45,   -28,   -59,   -47,    -3,    -3,    -6,     1,     7,    -3,    -7,   -31,   -38,   -49,   -61,    42,    27,    10,   -48,  -129,   -66,    34,     4,   -22,   -60,   -89,   -69,   -61,   -48,   -47,   -42,    -9,   -17,    18,     3,    -8,     0,    11,    11,   -46,   -53,   -66,   -50,    49,    30,   -36,   -77,   -98,     9,    13,    -7,    -3,   -74,   -94,   -81,   -64,   -36,   -36,   -53,   -36,   -15,    -6,   -24,    -4,     5,     3,   -21,   -34,   -51,   -38,   -26,   -21,   -18,  -117,   -90,  -134,   -11,   -30,   -39,   -60,   -94,  -118,   -77,   -53,   -39,   -30,   -72,    18,   -36,   -45,   -17,     5,     4,    -7,   -34,    -6,    16,    58,   -13,   -38,   -30,   -12,   -74,   -94,   -32,    -6,   -44,   -31,   -52,     6,    40,    16,     3,    -8,   -63,     4,   -84,   -23,   -27,    -5,    -2,    -7,    -8,   -23,    56,    -3,   -15,    21,   -17,    -5,   -82,   -96,   -24,     4,    -9,    17,    -1,     8,    28,    48,     5,   -16,   -16,     2,   -27,   -50,    -7,     4,    -7,    10,   -16,   -38,   -15,     3,     2,    21,    23,   -13,   -19,   -52,   -14,     0,     8,    48,     5,   -19,    28,    42,   -12,     5,    24,    -7,   -38,   -45,   -32,     1,    -4,     9,    43,    42,  -103,   -16,   -39,    -8,    84,    16,    -7,     2,    25,    32,    24,    48,    20,    55,    43,    30,    17,    70,    36,     3,   -20,   -17,    10,    30,    29,   -13,    66,    58,    30,   -12,    27,    29,    36,    54,   -32,   -14,    29,   -10,    -3,    10,   -12,    23,     8,    34,    43,     3,   -18,    14,    23,   -27,    -1,    21,    18,   -28,    38,    24,    87,    56,     8,    19,    20,     1,    -6,     7,    -3,   -48,    -1,    -4,    -7,    -7,    -1,    21,    34,    30,    43,    48,    44,    18,    -4,     8,    -2,     4,   -12,    -1,    26,    64,   -30,   -51,    18,     4,   -24,     2,    -7,     8,    14,    -1,   -14,   -56,  -138,  -114,   -84,   -21,   -40,   -42,   -40,    24,     6,    -1,   -10,     2,   -15,   -13,   -30,   -19,   -26,   -15,    20,    13,   -14,     9,    -2,    15,     2,   -49,   -64,   -40,   -72,   -41,    -1,   -34,   -33,   -59,   -15,    11,     5,     3,     4,    -1,    -3,     3,    -2,   -11,     2,    15,    18,    -8,     1,   -10,   -65,     7,    16,   -38,  -121,     0,   -17,   -36,   -45,   -39,   -26,    -2,     3,     7,     7,     9,     1,     3,     5,   -20,   -31,   -11,    -8,   -26,   -30,    -4,     1,   -66,   -64,     9,    27,    33,   -37,    -8,     5,     3,   -12,    -9,     7,     9,     0,    -2,    -5,     5,     6,     6,     7,     2,    -4,    -1,     0,    10,    -8,   -25,   -23,    -9,   -19,     7,   -19,   -30,    -3,    -5,     0,    -2,     8,     4,    10,   -10,    -5,     0,     9),
		    42 => (   -9,    -8,     7,     5,    -6,    -5,     4,    -8,     9,     3,    -3,     3,   -10,   -13,    10,    15,     1,     6,    -2,    -9,    -4,     2,     0,    -4,    -8,    -1,    -3,    -5,     5,    -6,    -3,     9,    -3,    -5,     0,     0,     9,    -1,   -24,   -20,   -18,     3,   -22,   -25,     8,     2,    -9,   -67,   -23,   -19,   -16,     2,   -10,    -7,     1,     0,    10,    -2,    -6,   -25,   -15,    -2,    -3,   -12,    -8,    -2,    46,    52,     4,    13,    26,    28,    47,    55,    18,    -5,    -2,   -15,   -24,   -15,     6,     6,    -7,     1,    -8,     5,    -3,   -37,   -43,   -22,    -8,   -25,    23,    25,    60,     3,   -15,    -7,   -19,    -9,    10,    50,   -37,    -6,    -7,    27,    -3,   -25,   -11,   -17,    -3,     6,     0,    -9,   -19,   -31,     0,   -12,   -18,    -5,    43,    85,    37,    -3,    40,   -15,   -18,    -5,    28,    14,    15,   -12,   -47,   -32,   -11,   -35,   -41,   -27,   -65,   -34,    -7,    -1,   -12,    -2,   -10,     3,    12,    23,     4,     8,    27,    63,    20,    48,    46,    25,    47,   -13,   -12,    29,    17,    -1,   -42,   -38,   -34,   -11,   -86,   -32,     6,     5,    15,   -26,   -12,    28,    31,    54,    24,    14,    25,    15,    -8,   -20,    13,    31,    39,    16,    41,     0,    18,    41,   -24,   -92,   -94,    -7,   -71,   -13,     7,    -3,    31,   -17,   -11,    22,    30,    41,    20,     7,   -20,   -13,    36,    28,    -4,    32,    30,    15,     0,   -23,   -14,    10,   -44,   -54,     6,    41,  -107,   -45,   -25,    37,    39,   -13,    -5,     8,    18,     8,   -19,    -5,   -24,    16,   -20,   -21,   -17,   -38,    10,   -22,   -30,   -16,   -52,   -25,    -9,    58,    29,   -14,   -73,   -43,     5,   -44,    44,    13,     4,     6,    11,     1,     5,    24,    31,     3,   -25,   -31,   -41,   -17,   -18,    -8,   -53,   -41,   -18,    10,   -16,    37,    -8,   -58,   -26,   -17,   -10,   -18,    50,     0,    16,     4,    -3,    -6,   -25,    -5,     8,    15,    56,    -6,   -14,    -5,    -6,    15,   -37,   -32,   -26,   -21,   -49,   -44,   -20,   -33,   -16,   -35,     0,   -24,   -15,   -31,    -2,    15,     3,   -13,   -10,   -41,     2,    13,    29,   -36,     0,    20,     2,   -16,   -53,    -9,    14,     1,   -28,    10,   -21,    26,   -44,   -55,     5,   -24,   -61,   -18,     2,    -6,     6,   -23,    26,    60,    33,    18,    39,   -35,     9,     6,   -12,    -8,    -1,    45,   -17,    27,    51,    36,    -6,    -5,    -2,     1,     1,   -12,   -30,   -37,    -8,    -2,    31,    31,    43,    20,    -1,   -19,    -2,    -4,     1,   -18,     4,    19,    42,    54,    34,    36,    38,    19,   -19,   -29,    51,     4,    -4,   -31,    -9,    -5,   -44,   -51,    10,    70,    50,    10,   -25,   -12,   -29,   -35,   -48,   -24,   -20,     1,    66,    49,    31,    54,    62,    74,    61,    13,    39,    39,     9,   -22,    38,    13,   -38,   -21,    -1,    16,    53,    22,   -30,    16,   -15,   -73,   -61,   -21,   -17,    10,     8,    54,    61,    46,    29,    47,     7,     8,     4,    35,     3,    -3,    42,   -28,   -39,   -40,   -15,    37,    26,    24,    14,    24,   -35,   -50,   -42,    38,     7,    20,    70,    71,    62,    80,    43,    97,    30,    39,    55,    27,    -2,    -3,    41,   -10,   -46,   -22,   -25,   -12,    37,    58,    53,    35,    21,   -13,     2,    21,   -30,    -2,    53,    87,    49,    17,    15,    14,   -17,   -31,    42,    30,    -2,    -2,     6,   -19,   -23,   -14,    -4,     5,    20,    45,    79,    36,    -6,   -15,   -31,   -14,    -4,    45,    77,    96,    73,    25,    13,    21,    23,   -43,   -19,    48,     6,   -15,   -30,    -4,   -12,    -3,    -8,    11,    21,    55,    42,    24,    19,   -54,    -5,     8,     4,   123,   132,   114,    45,    27,    35,    13,    12,   -46,    -2,    33,     0,   -21,     9,    15,     6,   -40,   -49,     4,    28,     9,    39,    31,    36,   -12,   -32,    19,    94,    84,    91,    62,    32,    -3,   -36,     6,   -11,    -9,   -24,     1,    -5,    -5,    30,     0,    48,   -15,   -50,     4,     1,   -23,   -20,     2,     1,    13,   -10,    65,   105,    94,    72,    74,    19,   -11,   -11,   -22,   -44,   -19,     4,     5,    -5,   -10,   -13,     4,   -21,     2,   -39,   -24,    -2,   -24,   -19,    -3,    42,    -7,   -11,    64,   138,    89,   118,    41,    26,   -10,   -10,   -17,     2,    32,    -2,    -6,     1,     7,    -6,    -6,   -23,    -3,   -19,     2,    27,   -26,   -78,   -51,    -2,     9,    52,   109,   149,   120,    94,    44,    -1,    29,   -35,    -3,    21,    24,   -35,     6,    -8,     6,   -26,   -36,  -108,  -107,   -32,   -23,    -6,   -72,   -58,   -37,   -29,    48,    69,    52,   107,   103,    76,    21,    -4,     1,   -24,   -14,    23,     2,    16,     8,     8,     8,    -3,   -19,   -42,   -70,    45,    14,   -12,   -28,    -1,    51,    81,    98,   108,   100,    71,    33,    37,    19,   -13,   -21,   -65,    -7,     9,    25,    16,     1,    -5,    10,    -4,     1,   -18,   -52,   -76,   -71,   -70,   -77,   -83,   -42,   -60,   -54,   -73,   -54,   -54,   -53,   -46,   -64,   -26,   -25,   -77,    -1,    -6,    -3,     8,     7,    -7,     0,     5,     9,   -15,    -8,    -7,   -12,   -14,    -8,   -15,   -17,    -7,   -17,   -20,    -7,   -11,   -12,   -17,    -6,   -42,   -61,   -10,   -13,   -10,     6,    -8,    -5),
		    43 => (   -8,    -5,    -7,     2,    -3,    -4,    -2,     8,     9,     5,    -2,     3,    -1,     0,   -13,    -2,     5,    -1,    -7,     3,     5,     2,     6,     6,    -5,    -1,    -7,    -1,     3,    -2,    -4,    -1,    -9,    -6,     3,     2,    -8,    -6,   -18,   -22,   -16,   -35,   -28,   -63,   -87,   -96,   -36,   -10,    -2,    -8,     1,    -7,     9,    -2,    -1,     3,    -5,     5,     0,    -8,   -16,     5,   -21,   -35,   -65,   -65,   -14,     0,    -7,    -7,     0,    -2,    16,    -6,   -34,   -27,   -39,   -46,   -47,   -59,   -21,     1,     1,     0,     1,     0,    -1,   -25,   -14,    12,    -4,    16,    40,   -14,     0,    16,    57,    -7,    -4,    58,    65,    46,    20,   -36,     6,   -28,   -46,  -106,   -87,   -35,     7,    -1,     2,    45,   -69,    16,    20,   -22,   -47,   -52,    17,    33,    49,   -13,     2,    -1,    -8,     9,    34,   -18,   -27,   -46,   -39,   -10,    52,   -51,  -104,   -94,   -24,    -2,    -1,     3,   -18,    13,   -19,    -3,    15,    19,    -8,     6,    -7,     5,    -6,    20,     7,    18,    29,   -17,   -61,    -7,    27,   -18,   -28,    52,   -13,  -110,   -39,    -5,    -6,    10,   -43,   -19,   -44,     4,    40,    31,     7,     8,   -10,   -46,   -49,     2,    23,    37,    27,    53,    32,    25,    21,    43,    16,    18,    66,   -99,   -84,   -40,     4,    -6,   -10,     8,     7,     2,     5,    15,    -2,    -5,   -28,   -15,    -8,    14,    19,     4,   -21,    33,    37,    14,   -19,    13,   -12,    82,    37,  -134,   -78,   -45,   -31,   -12,    21,    33,    10,    -1,   -20,    10,    -8,   -20,    18,    -8,    39,    36,   -27,   -45,   -11,    14,    23,    51,     7,   -36,    38,    37,     6,  -148,   -96,    -6,    -1,   -56,    -1,   -17,    28,    -6,   -39,   -53,   -48,    -3,   -53,    -8,    92,    64,    25,    11,    31,    11,    -8,    13,    40,    -3,    60,    43,   -75,  -117,  -102,   -40,     5,   -55,    12,    21,   -28,   -33,   -63,   -66,   -75,   -78,   -90,   -21,    55,    83,   104,    34,   -28,   -17,   -31,   -23,     4,    22,     8,    20,   -75,   -48,   -76,   -41,    -4,   -31,   -10,    43,     6,   -36,   -90,   -82,   -36,   -61,  -115,   -24,    15,    84,    52,    46,    17,     6,    -6,   -30,   -18,   -29,   -40,   -75,  -192,   -97,   -62,    -9,     3,   -15,     6,     4,   -15,    -1,   -36,   -66,   -23,  -105,   -21,   -45,    20,    47,   119,    59,   -12,    24,    25,   -28,    -1,   -18,  -115,  -134,  -141,   -70,   -51,    -9,    -1,    -8,  -118,   -25,   -32,   -36,   -16,   -34,   -10,   -42,   -51,   -27,     8,    38,    82,    30,    74,    16,    21,    18,     9,   -34,   -79,   -33,   -83,   -83,   -56,   -10,   -12,    30,     4,   -69,   -74,   -49,   -32,   -39,   -33,   -15,   -57,   -17,    -2,    42,    32,    49,    20,    -1,   -44,   -35,   -39,   -55,   -28,     7,   -66,   -76,   -43,   -13,    -3,    17,     0,   -44,   -11,   -11,    13,    -7,    14,   -67,   -65,    16,    62,    63,    49,    61,   -17,   -64,   -74,   -33,   -21,    -8,    36,    36,    28,   -57,    11,   -30,     1,     6,    19,    35,     6,   -20,     0,     5,     0,   -30,   -11,    34,    23,    12,    49,   -19,   -77,   -44,   -21,   -10,   -37,   -34,    46,     8,    29,  -106,   -70,   -34,     1,    13,    25,    30,    19,   -39,   -16,   -16,   -51,   -35,    -7,    48,     6,    26,    -4,   -52,   -66,   -38,   -38,   -13,   -52,   -13,     5,     5,     3,   -83,   -18,   -28,   -21,     8,    33,    45,     0,   -12,    14,    33,   -27,   -15,    36,    60,     0,     2,   -25,   -30,   -19,     4,   -26,     8,    16,    27,   -23,   -24,   -44,   -72,   -15,   -40,    -1,   -31,    26,    75,    35,    52,   -27,    34,    -2,    19,    47,    13,   -42,   -29,   -58,    12,    10,    25,    25,     5,    17,    15,   -36,   -18,   -27,   -57,   -71,   -40,     2,   -30,   -51,    16,    -2,   -37,   -38,    21,    32,    10,    31,    15,   -52,   -16,   -18,    32,    35,    14,    -4,   -12,    -8,    16,   -23,    -4,   -37,   -47,   -11,    -1,    -7,   -12,   -32,    15,     4,   -57,     2,    39,    39,   -13,   -30,   -29,   -25,     7,   -13,     4,   -10,     3,    -4,     3,   -26,   -22,    -2,   -37,   -89,   -58,   -24,    -7,     2,     0,   -15,    20,   -38,   -24,    42,     3,   -36,   -20,   -14,   -16,    -6,     5,     0,    -3,   -10,    12,   -17,   -17,   -11,     8,    -2,   -64,   -79,  -105,    -9,    -2,     0,     3,    21,    61,   -14,     5,    51,    16,    31,    10,    45,    24,   -29,    26,   -36,    -1,    33,    -3,    31,   -10,   -24,   -36,   -41,   -53,    54,    10,   -33,     7,     4,    -7,    23,    60,   -12,    -1,    17,     6,   -26,   -33,     5,    84,   -46,    -5,    58,   -15,   -13,   -28,     2,     4,    -6,    -9,   -26,   -27,   -56,   -49,   -20,     9,     7,    -1,     8,   -31,   -37,   -31,   -48,    14,    22,     3,    70,    67,   104,    32,    -5,   -33,    28,     2,    12,    37,   -42,   -87,  -101,  -113,   -52,   -11,   -18,     4,    -4,     9,     2,   -32,   -71,   -34,   -38,   -17,    -8,   -20,    32,    20,    39,     9,   -61,   -35,    -5,     9,    17,   -32,   -28,   -59,   -80,   -53,    -2,     2,    -9,    -5,    -9,    -4,     5,     9,   -18,   -28,   -22,   -18,   -18,   -56,   -59,   -66,   -51,   -97,   -40,   -44,   -29,   -15,   -16,   -58,   -65,   -29,    -3,    10,    -4,     2,    -3,    -6),
		    44 => (    5,     6,     9,     8,    -9,    -5,     8,    10,     6,     9,     4,     3,     1,    -1,    -8,    -6,     1,     1,    -4,     9,     0,     4,    -5,    -5,     9,    10,     4,     8,    -3,     5,     8,    -9,    -1,   -10,   -10,   -15,    -1,    -8,   -48,   -19,   -67,   -53,    -5,   -32,   -24,    -2,    -8,    -6,   -30,    -4,   -11,   -19,    -9,    -7,    -1,     7,    -6,    -9,    -9,   -51,   -54,   -60,   -25,   -44,   -37,   -33,   -14,   -62,    15,     6,   -31,   -73,   -47,   -39,   -39,   -14,   -17,   -22,   -31,    -7,    -5,    -8,     8,    -7,    -9,    -9,    -1,   -65,  -100,   -54,   -58,   -53,   -65,   -39,    31,   -24,   -61,  -123,   -74,    -8,   -17,    -6,   -51,   -55,   -11,   -16,   -40,   -21,     1,   -23,    -3,     9,   -10,     6,   -11,   -41,   -20,    14,    17,     3,   -12,    -1,   -53,   -91,   -10,    14,   -81,  -104,  -114,  -102,   -56,   -18,    -8,     2,    18,    31,    44,    13,   -28,   -15,    -2,     7,   -12,    -9,   -11,     1,   -19,   -17,   -56,   -89,   -71,     5,    56,   -20,   -40,   -15,   -47,  -192,  -101,    11,    45,    16,     4,     3,     2,    -3,   -26,   -17,    -8,    -2,    -2,   -38,    29,    98,   -13,   -62,   -36,   -28,   -47,    16,    44,    14,   -34,   -36,  -138,  -150,   -61,    45,    31,    13,     1,    31,    41,   -93,    29,   -80,    -2,   -69,    -7,   -32,    13,    83,   -43,   -24,   -19,    -8,    14,    26,    -3,    28,   -12,   -74,  -162,  -152,   -10,    51,    24,   -16,     4,    23,   -18,   -24,    31,   -84,   -28,   -59,    13,   -19,    -1,    20,   -31,    17,   -34,     0,   -27,    -6,    29,    23,     8,   -77,  -197,   -59,    26,    25,    14,   -15,    38,   -38,     2,    54,    23,   -53,     5,   -50,     6,   -27,   -12,    14,   -27,   -19,   -22,     8,    -4,     6,    48,    50,    33,   -99,  -101,    27,    50,    18,    25,    15,    21,    16,    54,   -50,   -49,   -33,     7,   -33,   -47,    14,    29,    49,     2,   -26,    -5,    15,   -17,   -15,    -7,    64,   -24,  -109,   -73,    16,    51,    42,     6,    -8,    20,    33,    16,   -92,   -30,    -6,    -9,   -21,   -26,   -63,   -27,    21,    50,   -10,    23,   -21,    13,    -4,    48,   -22,   -74,  -108,   -64,   -25,     8,     9,   -46,    34,     1,   -11,    36,   -45,   -44,   -36,    -6,    -1,   -47,   -59,   -83,   -25,    12,    40,    33,   -32,   -12,    32,    43,    25,   -90,   -50,   -13,    -9,   -15,    32,     0,    46,    11,    35,   -55,   -47,   -93,   -54,     6,   -14,   -53,   -59,   -69,   -38,   -11,   -11,    21,    21,    34,    46,    11,    15,     4,    13,    15,    31,   -26,    32,    28,    18,    -6,   -21,   -93,   -77,   -74,    -1,    -7,    -9,   -12,   -62,   -48,    -5,    -7,     2,   -10,    28,     8,    30,     7,   -14,    32,     8,    -4,     3,   -15,    29,    12,   -21,   -26,   -13,   -45,   -52,   -60,     0,    -2,    -2,    -8,    19,    -2,     0,     2,   -10,    25,     9,    29,    23,    -1,    11,    21,     4,   -16,    -9,     2,    52,   -98,   -29,   -16,   -11,   -47,   -71,   -50,    -2,    -3,    -8,   -25,    16,    -2,   -16,   -67,    -6,     7,     5,     2,    -2,   -10,     1,   -27,     4,   -11,   -19,   -17,   -22,   -71,   -39,   -23,   -39,   -57,   -78,   -77,   -16,    -4,     1,   -32,    15,    42,    -6,   -48,   -22,   -31,   -16,   -16,   -14,    -2,     1,   -13,     4,   -26,    13,   -11,   -51,   -79,    14,   -15,   -16,   -59,     5,   -13,   -20,   -36,     7,   -41,    67,    89,   -39,   -25,   -50,   -38,   -45,   -89,    -2,   -33,     5,    10,    -8,    10,   -42,    -1,   -19,     7,    37,    18,    18,     0,    34,    -4,    -9,    -3,   -44,   -20,    56,    28,   -41,   -54,   -33,   -18,   -49,   -52,   -12,   -42,     5,    -9,   -25,    -5,     8,   -18,   -20,   -12,    16,    11,    16,    36,    23,   -10,   -18,    10,     2,   -15,   -69,   -63,   -75,   -66,   -39,   -51,     0,   -28,   -30,   -39,    -2,   -13,   -23,    12,    -7,   -24,   -25,   -66,   -57,   -39,   -20,   -62,   -90,   -16,     4,     4,     1,   -16,   -41,   -68,    81,    -7,    13,    51,    65,   -18,    -8,     4,    -7,   -20,   -14,    -9,   -68,   -58,     7,     8,    -9,     9,    25,   -34,  -120,   -40,   -10,    -8,    10,     4,   -45,   -76,    44,    50,    32,    29,     1,    32,     3,    -1,    -3,   -26,   -14,     3,   -29,   -53,   -23,     0,     8,    -4,    32,   -39,   -36,    18,     9,     7,     4,    -1,   -42,   -65,  -127,    20,    31,    26,    22,    16,    -3,    20,   -12,    13,    15,    40,   -28,   -25,   -15,   -10,    21,     9,    21,   -24,     7,    24,     7,     5,     5,    -5,   -15,   -99,   -83,   -14,   -41,     1,    14,    23,   -14,     8,     0,    -4,    37,    17,   -45,  -107,   -25,   -19,    29,    15,    29,   -40,    42,   -30,    -9,     9,    -9,   -16,    -6,    -2,   -59,   -52,     1,    -7,   -32,     2,     8,    17,    28,     2,   -38,   -42,   -90,   -55,   -39,   -10,   -17,    25,    57,   -11,   -26,    -5,     1,     4,    -5,    -2,   -50,     5,   -55,   -52,   -87,   -43,   -54,   -57,   -39,   -74,  -104,  -118,  -158,   -33,   -43,   -66,   -32,   -40,   -42,   -31,    22,     2,    -8,    -4,    -5,    -2,    -4,     0,     5,     8,    -1,   -28,   -40,   -35,   -26,   -55,   -66,    -9,   -36,   -57,    -4,   -45,   -60,   -32,   -29,     4,    -9,     6,    -1,    -5,    10,     6,     4),
		    45 => (   -2,    -9,    -3,     0,    -7,    -9,    -2,    -9,     9,    -9,     4,     7,     5,    -5,   -10,     4,    -9,    -7,     6,     6,     1,    -6,    -4,    -1,    -4,    -4,     8,    -6,     0,     0,     4,     0,    -1,    -7,    -7,    -1,     7,     2,    -8,   -18,   -17,   -18,   -26,   -39,   -45,   -35,   -50,   -49,   -48,   -39,    -6,     1,     4,    -2,   -10,     9,    -5,    -5,   -17,   -20,   -22,    -5,   -10,    -9,   -52,   -13,   -28,   -19,   -38,   -49,   -51,   -47,   -14,   -27,   -32,   -33,   -27,   -41,   -39,    24,   -67,    -9,    -3,    -9,    10,    -1,   -10,    43,    93,   -16,   -39,   -44,   -14,    20,   -14,   -61,   -50,   -81,   -68,   -33,    23,     4,     6,    -6,     4,    16,   -65,   -54,     1,    78,    70,     4,     3,     8,   -28,    74,    -3,    -3,   -44,   -39,   -35,    -9,    -5,   -72,   -79,   -55,   -41,   -28,   -53,   -48,    -3,    49,    -4,     0,   -47,     3,    62,    51,     5,   -22,     6,     1,   -51,    81,   -20,   -17,   -26,   -49,   -43,   -22,     3,     2,   -64,   -26,   -22,   -14,   -30,   -10,    -9,    34,     8,   -10,   -25,   -16,   -24,    18,    -4,   -21,    -5,    -2,   -40,   -14,   -26,   -19,   -29,   -52,   -26,    -7,    -9,   -45,    -4,     6,   -11,     2,    -7,   -38,    -3,   -19,   -22,   -40,    64,    48,    31,    64,    70,     3,     3,   -11,     8,   -21,   -16,   -38,   -29,   -37,     7,   -15,    -2,    -5,    23,    28,    30,    15,    34,    44,    -9,   -33,    -2,    24,    22,    26,    18,    -4,    82,    19,   -25,    -7,   -42,   -12,   -22,   -33,   -21,   -16,   -15,     1,     3,   -11,   -13,     3,    27,    -7,   -12,    10,     8,    74,    84,    39,    59,    47,    17,   -12,    29,    39,    10,   -18,   -81,   -58,   -27,   -29,   -41,   -22,   -13,   -25,   -28,    -4,    19,    -1,    17,     1,    -5,    13,   -19,   -44,    26,    11,    24,    40,   105,    83,    17,    20,     1,    -7,   -36,   -42,   -45,    23,   -21,    -2,     8,   -26,   -31,    -3,    34,    -6,    -3,    14,    34,   -46,  -163,  -173,   -94,   -83,   -88,   -30,    -2,    21,    10,    32,     0,     6,     0,    35,    18,    21,   -17,   -19,   -37,   -70,   -14,   -45,   -52,   -34,     3,    -8,     8,   -11,   -86,  -101,  -150,  -138,  -139,  -109,   -88,   -19,    -3,   -20,     6,     0,    -3,    45,    21,    -9,   -52,   -70,   -60,   -45,   -14,   -44,   -61,    -3,    28,   -13,   -21,    16,     2,   -17,   -64,  -115,  -102,  -181,  -117,   -58,    -9,   -33,    -4,    -9,     0,    56,    -7,   -26,   -15,   -24,   -34,    -3,   -19,    -1,    40,     9,    17,    18,    -9,    12,    27,    52,    31,    34,    -4,   -66,   -94,   -28,     5,   -38,    12,     0,   -14,    33,   -40,   -58,    -6,   -39,   -48,   -11,    -2,    22,    -9,     5,     8,    36,    30,   -32,     0,    18,    47,   -14,     0,    43,    21,   -28,   -17,   -33,     9,    -4,   -36,     6,   -32,     0,    23,    -9,   -20,   -54,   -16,   -24,   -23,    28,     3,   -40,   -24,    -5,   -21,   -15,    49,    -5,   -13,    37,    64,    -2,    -5,    -6,    -8,   -27,   -75,     3,    10,   -50,    52,    12,     6,   -77,   -64,   -70,   -43,   -14,    -6,   -27,    24,    17,    -1,    -2,    57,    42,     1,   -30,     8,    26,   -15,   -16,    -8,   -31,   -91,   -31,    39,   -11,    44,    85,    35,     5,     7,   -48,   -89,   -39,   -46,   -40,     1,     0,    -7,   -26,    34,     0,   -72,   -55,   -12,   -11,   -29,   -18,    -7,    -4,   -70,    -6,     9,    16,    26,    66,    39,     7,    15,   -22,    -2,   -26,    -2,    -2,    -6,     5,   -26,   -33,   -25,   -16,   -37,   -73,   -47,   -22,   -57,   -50,     6,   -14,    58,   -64,   -23,   -12,    29,    54,    38,    56,    25,    42,    41,    31,    14,    -5,   -15,   -25,    15,    24,   -17,   -30,   -35,   -50,   -30,   -23,   -32,   -38,     8,   -11,    48,   -83,   -57,    -5,    -1,   -36,    14,    21,    29,    21,    20,    -5,     8,     0,    -8,    -5,    -4,   -20,   -15,   -31,   -16,   -17,   -16,   -15,   -10,    -7,    -7,     3,   -27,     1,   -36,    23,   -20,    -6,   -53,   -36,   -25,    21,   -22,   -12,    16,     0,    14,    13,    12,   -22,   -38,    -2,    -6,   -13,   -15,   -15,    -9,    -7,    -4,    -5,   -80,    25,    32,    -4,   -41,     3,   -52,   -25,   -20,    -9,     0,   -15,    11,     8,     2,     1,    -2,   -33,    -2,    23,     8,    -6,   -12,    -9,    -5,     7,     4,    -7,     9,    14,    47,    61,     7,   -32,   -42,   -39,    -4,    -5,   -37,   -49,    -6,   -22,    -1,    28,    34,     3,    -2,    23,    15,    -4,   -35,   -17,   -11,   -10,    -6,     3,   -38,     0,   -12,   -14,   -45,   -84,   -73,   -28,   -84,  -101,   -36,   -10,   -28,   -41,   -54,   -34,     6,    30,    25,    -2,    20,     5,    12,   -48,   -19,    -3,     4,     9,     1,    18,   -33,   -21,     3,   -20,   -52,   -13,   -92,   -87,     7,   -23,   -27,   -12,    -3,   -14,    -8,    -8,   -11,   -33,    13,     3,     9,     6,   -10,    -6,     8,     8,     9,   -11,   -17,   -21,   -34,   -19,   -26,   -21,   -15,   -22,   -17,    33,    73,    68,    56,    28,    -5,    40,     3,   -18,     2,    -8,    -7,     7,     6,    -1,    -3,    -8,     8,     7,    -3,   -13,    -5,     2,    -5,     1,     6,    -2,    -3,     1,    -7,    -1,     0,     3,   -19,   -18,   -16,   -17,   -52,   -10,    -1,    -2,     7,    -7),
		    46 => (   -6,     5,    -8,    -3,   -10,    -6,     0,    -5,   -10,     0,     9,    -2,     3,     5,    -9,     7,     2,     2,    -6,     9,    -4,    -8,    -7,    -8,     8,     1,     6,     5,    -5,     5,    -2,    -5,    -2,    -2,    26,    38,    53,    57,    28,    19,     7,    18,    18,     7,     2,    -5,    12,    14,    68,    22,    12,    19,    -4,     3,    -5,     2,     0,    -4,     9,     6,    11,     3,    41,    57,    58,    29,   -18,   -16,   -17,    -1,    -7,    -6,   -10,   -25,    -9,    35,    31,    10,    12,    35,    32,    10,    -8,     0,     4,    -4,   -46,   -31,     3,     7,    25,    43,    17,    31,     3,   -42,   -49,   -16,    -6,    -7,    -4,    -9,   -10,    14,     2,    31,    -3,    37,    45,    -1,   -19,    -3,    -2,    -9,   -24,   -11,     4,    12,    11,     6,     8,    10,   -30,   -27,    -1,   -26,   -13,    26,    20,     1,   -10,     0,    -7,    18,    -1,    16,    11,     4,    22,    29,    -7,     6,     7,   -17,     9,   -19,    -7,    10,     8,   -23,   -41,     6,    -3,   -23,    15,   -17,   -32,     9,     9,     7,    17,     0,     7,    21,    23,     6,    49,    31,     4,     0,     2,    -5,   -10,    -5,   -19,     8,     2,   -17,     8,    -8,     7,   -27,   -29,   -41,   -51,    -6,    11,    19,    26,    38,    26,    18,     1,   -29,    15,    20,    -4,    -1,     7,   -15,    -4,   -12,   -25,   -28,    13,     7,     3,   -13,   -46,   -21,    17,     3,   -23,   -13,   -27,    -6,    -2,    -8,   -13,   -10,    20,   -17,     7,    12,     5,     6,    -5,   -33,   -11,     0,   -15,   -33,    13,    12,    -6,   -44,   -29,   -10,   -11,   -30,    15,    22,   -22,   -24,   -41,   -15,   -59,   -50,   -35,   -38,   -13,   -41,     3,     7,    -5,   -10,   -19,   -39,     2,     0,    28,     5,   -17,   -31,   -32,   -33,   -10,    15,     3,    -9,   -29,   -53,   -57,   -45,   -73,   -53,   -18,   -28,     6,   -10,    -2,    -2,     1,   -19,    -8,   -29,     0,   -14,    24,   -32,   -30,   -49,   -23,   -33,    -4,    18,    -5,   -42,   -48,   -25,   -45,   -35,   -49,   -51,   -19,   -17,   -14,   -24,    -1,     1,    -6,    -7,    -3,    12,    29,    -3,     6,   -26,   -52,   -32,   -12,     0,    22,    -3,   -48,   -54,   -42,     0,     6,     0,   -11,   -15,     8,   -29,   -20,    -2,     6,    -4,    -2,    -5,   -28,    16,     6,   -15,    -8,   -21,   -48,   -20,   -18,    13,   -11,   -30,   -30,    22,    16,    -5,    11,    21,    15,    12,    14,   -38,   -45,    -9,    -6,     4,   -12,    -8,   -16,    26,    -9,     9,    23,   -37,   -45,   -26,    12,    13,   -35,   -13,     1,    -4,    15,    18,    -9,    -9,     0,    20,    29,   -28,   -27,     5,    -8,    -8,     6,    -5,   -12,    40,   -12,    11,     9,   -32,   -32,    33,    20,   -10,   -32,    -3,     7,    36,    35,    32,    -3,   -31,    -9,    22,    25,   -10,   -18,   -22,     2,     9,   -14,   -12,    -6,    23,    -7,    -2,    -1,   -13,   -35,    -9,   -18,   -41,   -16,    16,    32,    26,    32,    40,    -7,   -16,   -13,    29,    33,   -20,   -23,   -43,    -9,     6,   -10,   -20,    -5,    13,   -10,   -35,    10,   -21,   -20,   -14,   -36,   -10,    10,     8,    15,    33,     3,   -25,    -5,   -11,    -3,     3,    -1,   -10,   -20,   -37,    -2,     5,   -19,    -3,    -2,   -30,    -1,   -41,    11,    -4,   -12,   -57,   -50,    -6,    19,     4,    -5,     4,    -7,   -19,    25,    20,    -6,   -10,    -1,     3,   -14,   -40,    -2,    -5,   -18,    -2,   -11,   -27,   -43,   -21,    22,    16,   -11,   -30,   -16,    15,     0,    11,    -3,   -22,   -16,   -17,    28,    -3,     1,   -26,   -19,    -1,   -43,   -31,    -3,    -8,     2,     1,    -5,   -29,    -3,    -8,    -9,     4,   -24,    11,    -2,   -17,     9,   -24,    -2,   -20,    -4,   -17,    19,    -9,    -9,    -7,   -10,   -16,   -17,     0,     6,    -2,     4,   -22,     8,   -15,   -19,    -9,    -3,   -20,    19,    -5,   -31,   -22,     7,   -11,   -36,   -14,    -7,     7,    26,    14,   -20,   -30,   -10,    12,   -15,    -3,    -9,     9,    -3,   -13,     2,   -20,   -24,     6,    -9,    14,    -7,    -1,   -27,   -34,   -13,   -20,   -13,   -18,    -4,    10,    19,   -14,   -37,   -17,   -25,     6,    -8,     2,     0,    -4,     5,    -6,    -1,    -3,    14,    -4,     2,   -13,    -2,   -21,    -9,   -17,   -27,    -1,     4,    -8,   -29,   -17,   -24,   -13,   -41,   -23,   -16,   -20,    11,    -5,    -7,     3,    -2,   -15,     6,    -1,   -18,   -15,    13,    14,     8,    14,    26,   -24,   -13,   -24,    18,    -9,   -28,   -43,   -25,   -37,   -15,   -10,   -19,     3,   -14,     6,    -7,    -2,    -9,     2,   -12,     1,   -15,   -24,   -18,   -23,   -18,    -2,    -3,   -20,   -18,   -28,     2,     4,    -7,   -41,   -42,    -8,    -9,   -10,    -3,    -8,    -5,     9,     1,     2,    -1,    -9,     6,    -4,   -19,   -12,    -9,     3,     3,    -2,    -1,    -2,     1,    -2,   -10,   -14,     1,    -2,   -29,    -8,   -14,   -32,    -8,    -7,     6,     2,    -5,     7,    -4,    -3,    -2,    -9,    -7,   -11,     0,     3,     3,     0,     7,    -9,     4,     1,    -8,    -5,    -6,    -4,    -7,   -22,    -4,     3,     7,     6,     7,     4,     9,     7,     3,     7,     1,     4,     4,     2,     2,    -5,     2,   -10,     5,     4,    -8,    -8,    -2,     6,     7,     7,    -4,    -9,     1,     2,   -10,     3,     6,     6),
		    47 => (   -3,    -2,     5,    -9,     5,     2,    -6,     8,     3,     1,     0,     7,    -4,     4,    -9,    -2,     4,     2,     0,   -10,    -2,    -7,    -5,     7,    -5,    -2,    10,    -5,    -9,     0,     2,    -7,     8,     9,     9,     0,    -8,     8,    -7,   -54,   -38,   -46,   -13,    -9,   -21,   -16,     5,     5,     8,     4,     6,    -8,    -1,    -7,     3,    -4,     7,   -10,    -2,    -5,    -3,    -9,    -4,    -2,     2,    -8,   -12,   -38,   -56,   -37,   -29,   -23,   -10,     5,     1,   -10,   -12,     2,   -12,    -3,    -9,     0,    -9,     8,     1,    -2,    10,   -19,   -21,    -9,   -15,   -33,   -27,   -19,     1,   -15,   -29,   -15,     3,   -43,   -43,   -27,   -19,    -7,   -17,    -3,   -36,    -9,   -12,     5,    -6,    -7,     7,    -7,    10,    -8,    -6,   -32,   -36,   -34,   -48,   -22,   -31,   -48,   -56,   -44,   -29,   -37,   -33,   -38,   -23,    -5,   -22,   -15,   -52,   -29,   -20,   -18,   -10,    -2,    -5,     7,    -5,   -27,   -20,   -51,   -64,   -41,   -11,   -13,   -49,    -8,    12,    -1,   -36,   -81,   -87,   -58,   -80,  -100,   -91,   -58,   -52,   -51,   -41,   -15,    -2,     9,    -7,     1,     7,    11,   -26,   -57,   -73,   -90,   -77,  -114,   -96,   -26,    34,    36,    12,   -30,   -57,    17,    28,     2,    19,    75,    20,    40,   -45,   -17,   -46,   -12,    -9,    42,    27,    40,    19,   -14,    39,    -3,   -37,   -99,   -90,   -85,   -65,   -17,   -11,   -51,    -2,     0,    21,   -31,   -62,   -31,   -25,   -15,   -12,     7,   -25,   -20,   -25,    48,   -21,    -3,    -7,     3,    41,    42,   -31,   -77,   -77,   -76,   -38,   -62,   -67,   -73,   -47,   -34,    14,   -34,   -40,   -64,   -24,    37,    19,     1,   -73,   -25,   -19,    43,   -24,   -21,    -1,    13,    67,    -6,    10,   -23,   -59,   -24,   -35,   -61,    -7,   -12,    -6,     4,     7,   -33,   -27,    56,    37,    77,    49,    16,   -48,     5,   -11,    25,    10,   -12,   -59,   -20,    27,     2,   -35,   -18,    -1,    -5,     4,    29,    12,     1,   -15,    42,    26,    25,    -6,    38,    34,    -4,   -34,   -11,   -54,    15,    -4,    12,     8,     4,    -1,    10,   -17,    47,   -15,     0,    -6,    67,    46,    32,    34,     0,   -27,   -23,     5,    22,    14,    22,    14,    23,   -13,   -29,   -10,    63,     0,    -2,    17,    41,    34,    34,   -34,    37,    45,     1,    10,    44,    60,    13,   -32,   -34,    28,    44,    10,   -13,    -3,   -15,    32,    -4,    54,    40,    74,    75,     5,    14,    35,    44,    34,    15,    15,   -48,   -15,     6,    31,    11,     2,   -32,   -36,   -36,    21,   -11,   -10,    -6,    44,    25,    35,   -56,    54,    52,    30,   -13,   -14,    36,    63,    46,    13,    79,     5,   -54,    21,    26,    39,   -11,   -77,  -103,   -29,   -30,   -16,   -29,    38,    12,    25,    23,    16,     8,     4,   -18,   -44,    -9,     7,    -9,     2,    65,   -45,    22,   -10,    31,    -1,    42,    40,   -41,  -126,  -108,   -59,    -9,    -5,    19,     0,    46,    36,    -5,   -13,   -61,   -53,   -13,    -3,    -1,     5,   -11,    -5,    31,    74,     5,    12,    16,    -4,    -2,   -37,  -154,  -178,   -36,   -20,    -1,    -8,     4,   -40,    14,    38,    26,    11,   -39,   -67,   -85,     4,   -36,     8,    -3,    38,    -3,    45,    -4,   -11,   -11,    -2,   -42,  -103,  -126,  -102,    -4,   -18,     9,   -33,   -11,   -22,   -31,    43,    29,    13,   -33,   -53,   -60,     9,   -52,    19,     5,    36,   -59,     2,   -13,     0,    31,    -8,   -87,  -128,   -58,   -34,     3,    14,     6,   -54,     0,   -19,   -19,    45,    22,     5,   -48,   -51,     2,     9,     0,    -2,    44,     8,   -63,   -14,    -3,    32,     9,   -31,   -94,  -109,   -39,   -21,    46,     3,   -13,    -6,    25,   -27,    21,   -11,   -26,   -21,   -51,   -45,    11,    -8,     3,    -5,     9,    -4,   -26,   -12,   -15,   -13,   -31,   -43,   -74,   -52,   -10,    12,     3,    10,   -23,   -41,    19,   -14,    -3,   -22,    -9,   -19,   -37,   -34,    -6,    -1,    -3,     9,    10,    -2,   -46,   -55,   -36,   -61,   -87,   -46,   -37,     8,    18,    -8,     4,    -4,   -28,   -32,    -7,    18,    16,     1,    14,   -16,   -46,    63,    -1,   -10,     7,     2,    -3,   -11,   -66,   -29,   -34,   -44,   -62,   -42,     4,   -14,     2,    14,    24,   -11,    19,   -17,   -34,    17,   -31,    47,   -17,    -1,   -48,     9,     8,    -5,    -2,    -8,    -3,   -12,   -46,     0,     8,   -56,   -27,   -11,   -31,    24,     8,    10,    -2,    -1,   -32,    -7,     4,   -17,     0,    22,   -38,    -8,   -46,    20,    -1,   -10,     8,    -1,     0,     1,    12,    25,     2,   -33,     3,    -5,    37,     1,    28,    16,   -51,    25,    -7,   -14,     0,   -28,   -55,    25,    10,   -16,   -59,    10,   -31,     6,     3,     3,     0,    -4,     5,   -15,    19,    17,    13,    -7,    -2,    22,    46,    31,     7,    54,    20,    35,    -2,   -15,    13,   -15,    12,    -1,   -59,    20,   -11,     9,    -6,     0,     6,    -2,   -14,    -8,   -27,     6,   -30,     0,    -2,   -42,    -1,    60,    41,   -12,   -23,     4,    13,   -24,   -40,     4,    23,    13,    12,   -11,    -7,    -8,     4,    -9,    -8,    -1,     2,    11,    24,   -12,    15,    39,    34,   -12,     3,    13,    32,   -13,   -24,    15,    42,   -50,    -9,    -2,    58,    57,    54,   -10,    -2,    -8,     6),
		    48 => (   -8,    -7,    -2,    -2,     2,     9,     4,    -7,    -6,    -5,    -2,     7,    -6,    -4,    -2,    -9,     7,   -10,     1,    -7,     6,     3,    -7,     5,     1,     3,     6,     8,     9,     1,    -1,    10,    -8,    -3,    -1,    -8,    -1,    -7,     2,    -6,    -2,    -6,   -14,    -7,   -26,   -12,   -15,    -1,     9,     0,   -10,    -6,     8,    -4,     4,    -4,     8,     7,     0,     4,     1,     0,    -4,   -10,   -32,   -37,   -54,   -42,     8,     3,     6,   -27,   -27,    -2,   -13,     7,   -39,   -35,   -32,   -15,   -21,    -7,     8,    -5,   -10,    -8,    -9,     2,   -17,   -29,   -43,   -38,   -27,   -28,   -33,    11,    29,    22,     7,   -21,    -2,   -11,    35,    12,     5,    -7,    -8,    66,     6,     9,   -16,    10,     7,    -6,     8,   -24,   -41,   -61,   -44,   -46,   -21,     9,   -17,   -10,   -26,   -37,     1,   -31,   -10,   -16,   -27,    33,    80,    91,    22,   -58,   -61,   -22,    27,    -7,     0,     2,   -22,   -14,   -52,   -28,   -24,    -9,    -8,   -25,   -18,     7,     2,   -31,    -2,   -78,   -57,   -40,   -54,    11,    48,    64,    31,   -25,   -41,   -16,     7,    -8,    -6,     0,   -20,   -67,   -11,   -25,    -8,     6,   -39,   -13,   -12,   -10,   -17,   -15,   -22,   -38,   -16,   -12,     6,   -16,   -14,    -5,    -9,   -21,   -49,   -30,     1,    12,    -1,   -16,   -12,   -41,    -3,    -1,     1,    -9,    -3,   -23,   -26,   -37,   -48,     1,     3,    13,     7,   -26,    -2,    56,     7,     1,    16,   -12,   -47,   -24,    15,    25,     1,   -36,   -13,    18,    14,    13,    12,    -3,    -7,   -28,   -39,   -60,   -54,   -48,   -15,    14,   -22,    22,    -9,   -26,     9,    53,    44,    -6,   -35,     8,    21,    48,    -1,   -23,   -31,   -18,    18,    -1,    13,    21,   -10,    10,    -6,   -39,   -58,   -87,   -39,   -23,   -21,   -10,    -2,    -9,     4,    23,    -8,   -14,   -13,   -21,   -11,    -5,     9,   -22,   -41,   -40,     4,    23,     1,    -3,   -20,    23,   -12,   -17,   -50,   -60,   -29,   -10,    22,    17,   -13,    33,    40,     3,    -9,   -12,   -15,   -51,    -2,   -21,    -4,     2,   -24,    30,   -22,     3,    15,   -14,     6,    21,    23,   -13,   -10,     1,   -17,   -60,   -13,    40,   -11,     5,    19,   -11,   -37,   -33,   -49,   -30,    -5,   -18,     2,     7,   -25,   -24,   -16,    -7,   -21,   -26,   -48,   -12,    18,    50,     9,   -36,   -51,   -49,    -5,    23,   -22,   -16,     6,     0,   -24,     2,     6,   -17,   -28,   -24,     0,     0,   -30,   -28,   -48,   -17,   -15,    -6,     0,    22,    11,    49,    25,    14,   -44,   -38,     6,   -17,   -74,   -23,   -24,   -17,    -4,   -10,   -37,   -30,     5,    -8,    -8,   -11,   -20,   -40,   -29,   -37,   -67,   -45,    13,   -33,   -12,    17,    12,    23,   -18,   -30,    10,   -40,   -51,   -56,   -51,   -18,   -39,   -27,   -51,   -18,   -61,   -24,   -12,    -4,   -16,    16,    -1,    -4,   -53,   -46,   -40,   -31,   -60,   -11,   -15,    30,    25,    26,    17,     1,   -53,   -62,   -47,   -11,   -32,   -22,   -18,    -9,   -44,   -40,   -10,   -12,   -18,    24,    -4,   -22,   -33,   -42,    -8,   -36,   -25,    -9,   -25,    18,   -33,   -12,   -12,    -1,   -48,   -23,   -35,    16,   -35,   -30,   -21,   -24,   -51,   -41,    -6,   -13,   -29,    27,    -6,   -30,   -46,   -42,   -79,   -81,   -14,     2,    23,    29,   -36,   -23,   -49,     4,     3,   -32,    21,    23,    46,   -10,   -30,    -4,    -6,   -24,   -17,    -9,   -14,   -12,   -12,   -25,   -58,   -53,   -53,   -33,    -7,    19,    52,   -17,     2,    21,   -20,    33,    10,     8,   -11,     1,    20,   -13,   -24,   -15,   -14,   -15,     5,     7,   -10,   -15,    -9,   -22,   -52,   -43,   -40,   -20,   -20,     3,    49,   -30,    -5,    25,   -42,    42,    41,    11,   -16,   -16,     7,    14,   -33,   -13,   -37,   -14,     9,     9,   -17,   -10,   -30,   -23,   -66,   -54,   -28,    -3,    28,    40,    32,   -23,   -27,     8,   -61,    47,   -25,    28,    10,    -3,    -5,     6,   -15,   -17,   -45,    -1,   -17,    -4,   -10,    -9,   -30,   -37,   -75,   -67,   -36,   -15,    23,    30,    10,   -37,   -16,    -6,     1,     1,     0,    27,    -6,     9,    15,    10,   -56,   -11,   -37,     7,   -12,     2,   -18,    -7,   -14,   -36,   -94,   -74,   -68,   -52,     3,     5,   -13,    14,   -23,     8,   -18,   -47,   -20,    -4,     6,    41,     9,   -38,   -33,    -3,   -27,   -12,     6,     8,   -21,   -25,    -8,   -24,   -39,   -33,   -57,   -40,   -11,   -38,    -2,   -12,    -4,    10,    -5,    18,   -26,    -5,    44,    12,    38,    -7,     5,    -9,   -22,     1,    -3,     4,    -4,     1,    -9,   -22,   -57,   -57,   -60,   -26,    -8,   -21,   -40,   -59,   -39,   -20,    39,   -32,    10,     6,    54,   -10,   -21,   -19,   -35,   -16,    -7,    -6,    -9,     1,   -26,    -6,   -24,   -28,   -22,   -57,   -52,   -47,   -33,   -42,   -33,   -37,    -7,    46,    56,    29,    34,    17,    17,   -20,    -8,    -8,    -7,    -4,    -2,     6,     0,    -9,     3,   -35,    -2,   -19,   -31,   -13,    -8,   -30,   -59,   -34,   -30,   -41,   -69,   -53,   -36,   -18,   -10,   -62,   -70,   -24,   -33,   -11,    -8,    -3,     5,   -10,    -6,    -5,     5,     2,    -8,    -3,    -8,    -7,   -13,   -14,   -12,   -18,     5,     2,   -23,   -14,   -28,   -31,    -1,     2,    -4,   -10,    -1,    -9,     9,     6,    10,    -4),
		    49 => (   -6,    -5,     2,     2,     3,     2,     7,    -8,    -4,     4,     0,     5,     1,    -2,    -1,    -3,     3,     7,     4,     4,     7,   -10,    -2,     5,    -8,     8,    -1,     6,     5,     1,     3,     4,     0,     0,     7,    -2,   -10,    -7,   -12,   -26,   -26,   -23,    -3,   -72,   -66,   -57,   -22,    -9,     6,   -13,    -1,    -9,    10,    -2,    -4,    -8,   -10,     5,    -5,   -17,   -12,     2,   -10,   -30,   -29,   -17,   -17,   -44,   -20,   -23,   -56,   -24,   -52,   -14,    -4,   -13,   -37,    -9,   -10,   -24,    -7,     9,     3,    -1,    -5,    10,    -4,   -81,   -24,   -23,   -11,   -42,   -50,   -64,   -59,   -58,  -114,   -80,   -94,   -90,   -85,   -41,    12,   -43,   -45,   -33,   -20,    -9,   -16,   -15,    -9,     6,     1,     5,   -24,   -26,   -26,   -60,   -82,   -58,   -46,   -79,   -60,  -110,  -129,   -30,   -74,   -52,   -31,     7,    25,  -134,   -70,   -89,   -51,   -13,   -11,   -56,   -50,   -13,    -7,     6,   -15,   -26,    -6,   -30,   -61,   -51,   -56,   -52,   -32,     9,   -19,    28,   -33,   -12,   -48,   -44,   -41,   -38,   -22,   -26,   -84,   -72,   -46,   -42,   -38,     3,    -8,   -14,   -19,   -73,   -86,  -177,   -90,   -11,     2,    72,    16,    30,    -9,    56,    -8,     7,    12,    26,    36,     1,    24,    20,   -54,   -55,   -84,   -76,   -48,   -32,     9,   -44,   -61,   -77,  -136,  -171,   -12,   -53,   -20,    11,    27,    32,    54,    12,   -15,    41,    -7,    25,    14,     2,    -8,     2,   -29,   -76,   -78,   -65,   -50,   -18,   -74,   -53,   -47,   -46,   -85,    -2,    -8,   -52,     8,   -22,   -13,    -1,     1,   -35,    -2,   -27,    -4,    -9,    23,   -23,    -3,    27,   -30,   -32,   -48,   -74,   -68,   -32,   -15,   -28,    -5,   -25,   -80,    -6,   -11,    -1,   -20,   -36,    -3,    16,    -4,   -13,   -25,    47,   -17,   -23,   -26,    10,     1,    26,     0,   -13,   -28,   -71,   -74,   -27,    -9,   -53,   -81,    -6,    17,     8,   -31,   -28,   -16,    19,   -13,    18,    15,   -28,   -37,   -38,   -16,    23,   -13,    17,    29,    10,    22,   -15,   -38,    94,   -75,   -51,     6,  -122,    38,   -14,    41,   -12,   -23,   -15,    22,   -12,    47,     7,     8,    11,   -32,   -16,     6,    49,    13,    15,    32,    35,    70,   -35,     8,    97,   -59,   -59,   -11,   -29,    20,    20,    74,    17,     9,    27,     5,    51,    -2,    24,   -52,   -62,    10,     2,    18,    49,    61,    67,    23,    45,    50,    73,   -78,  -149,   -89,   -17,     5,   -58,   -44,     8,    98,    76,    26,    58,    53,    32,    37,     4,    15,    16,    32,    25,    59,     0,    26,    41,    55,    40,   109,    21,  -127,   -80,   -55,     0,   -22,   -47,   -27,    17,    76,    62,    16,    25,    65,    18,    44,   -21,   -26,    16,   -13,     1,    41,     7,    29,    49,    -7,    22,   120,    -7,  -180,  -120,   -11,    -6,    -8,    -8,   -98,    21,    70,     7,   -32,    29,    77,    40,     5,   -43,   -33,    13,   -24,    39,    37,    64,    45,    41,   -22,   -43,    -4,   -43,  -160,   -92,    38,   -17,     7,    -8,   -87,   -54,    13,   -45,    -6,    -6,   -10,   -41,    48,   -41,   -20,   -22,   -20,    -4,    -9,     5,    -7,   -25,   -16,   -75,   -21,   -39,  -135,   -72,   -14,   -49,     6,     0,  -101,    -3,   -36,   -39,   -37,     9,    -5,   -23,   -21,   -60,   -14,   -29,   -30,    16,     9,    19,   -32,   -42,   -41,   -39,   -39,   -32,  -107,    -5,   -17,   -34,    44,    -2,   -94,    11,   -36,   -58,   -26,   -10,     6,    -9,     9,   -13,   -35,   -67,     0,   -14,   -11,    -4,    16,    -6,   -51,    10,    -6,   -85,  -184,   -19,   -48,   -30,     7,   -12,   -50,    65,   -30,   -69,   -58,   -63,   -42,   -49,   -44,   -35,   -53,  -113,   -19,    -7,   -30,   -26,   -14,    21,    -6,   -30,    32,   -43,   -84,    -9,   -39,   -15,    10,    -1,   -91,    49,   -27,    54,   -31,  -133,  -103,   -62,   -76,   -15,   -63,   -70,    15,   -25,     9,    10,   -29,    20,   -55,   -38,   -20,   -15,    12,    33,   -23,    -7,    -4,     2,   -91,    60,    16,    57,   -30,   -55,   -59,   -53,   -77,   -62,   -63,    -3,   -79,   -33,    10,   -30,   -49,   -29,   -63,   -17,   -30,   -66,   -32,    25,  -155,    -7,     9,   -10,   -83,    52,   -46,   -20,    14,    40,    43,    -3,    18,   -30,   -14,     0,     3,    15,   -22,   -35,   -48,   -72,   -25,   -10,   -12,   -70,     6,   -22,   -93,   -19,     4,     4,   -65,    45,   -13,   -32,   -26,    10,    -2,   -32,     3,   -38,   -28,    -2,    -2,   -44,   -36,   -28,   -26,   -16,    -4,    29,    32,   -18,    -2,    -3,   -15,     8,     1,     6,   -64,   -66,   -10,    32,   -43,    24,   -16,    -8,    15,    35,   -15,   -28,   -63,    -8,     9,   -40,     6,    19,   -29,     7,    46,    57,    -2,   -23,   -32,    -2,    -8,     6,    45,   -44,    58,    24,   -74,   -89,   -29,   -18,   -58,   -46,    16,    -7,    61,    -1,    28,    46,    44,    29,    67,    81,    15,   -12,   -24,    -2,   -37,    10,    -2,     2,     0,    35,    42,     0,    15,     3,    14,    15,   -37,   -10,    45,    12,    63,    13,    28,    68,    89,    24,    64,    62,    36,    38,    37,     9,     9,    -5,    -7,    -2,    -3,    -2,   -46,   -57,    21,    13,    29,    19,    -9,    18,     6,   -29,    43,    35,    23,   -79,   -26,    43,     5,   -49,    16,   -46,     6,    -7,     0,     3),
		    50 => (   -2,    -6,     4,     7,     7,    -4,    -1,     1,     6,     6,    -3,     5,    -5,     9,   -10,     4,     0,    -5,    -6,    -6,    -8,    -7,    10,   -10,     6,    10,     2,    -7,    -2,    -8,     9,     8,     9,     5,     4,     8,     8,    -6,    -3,     3,     6,    10,    -5,     6,    -7,    -8,     0,     6,    -7,    -9,     9,    -6,    -8,    -3,     8,     2,     3,    -4,    -2,    16,    26,   -16,   -15,   -11,   -20,   -25,   -35,   -59,   -66,   -67,   -35,   -48,   -38,   -38,   -17,     7,     9,    -2,   -42,    -9,     4,     3,   -10,     1,     7,    -9,     4,     6,    -2,    14,   -24,   -16,   -67,   -66,   -22,     1,     0,    24,    -4,   -52,   -66,   -30,   -19,    -5,   -15,    -6,   -18,   -10,    -5,    -8,    -9,     9,    -7,    -7,    -3,     8,   -17,   -56,    35,    -7,    39,    42,    23,    30,   -14,    -5,    -7,   -43,    -9,    19,    23,     4,   -46,   -65,   -15,    -3,    -9,    -5,   -19,    -2,     2,     6,     1,    17,     9,   -35,     1,   -18,   -57,   -10,    12,    27,    10,    28,    15,    -4,    25,     7,    17,   -11,   -14,   -15,    -2,    -9,   -31,   -42,   -33,   -41,     4,     5,   -27,   -14,    20,   -16,     0,   -24,   -25,   -10,    11,    14,     2,    -2,     6,    11,    41,    18,    23,   -14,   -11,   -44,   -18,    64,    40,   -50,   -53,   -12,     6,   -13,   -25,   -15,   -21,    29,    23,    15,   -11,    21,    42,    10,    10,     0,    20,     3,     1,    27,    -4,   -16,   -46,   -37,   -25,    25,    31,   -36,   -41,    17,    12,    -1,     7,   -26,   -24,    -1,    -5,     3,    36,    40,   -11,    -7,    54,    28,    34,   -20,     6,   -28,    -3,   -25,    -5,   -19,    13,     4,     9,   -39,   -56,   -23,    -5,     0,     1,   -17,   -45,    41,   -37,    -3,    -7,    16,    -3,    -1,   -16,    -5,     5,     6,   -29,   -44,    46,    44,    48,    20,    34,    -2,    55,   -62,   -53,    -7,     8,    -6,     2,   -17,   -64,     7,     0,    -7,    19,    11,    30,    -7,   -59,   -24,    -7,    -9,   -33,    21,    29,   -14,   -39,   -21,    56,    12,    49,   -41,   -35,    -8,     0,    22,   -29,   -36,   -50,    -5,     8,    -5,     4,     9,    27,   -53,   -58,   -58,   -47,   -59,   -18,    -7,     0,   -43,   -30,   -42,   -26,     8,    33,   -22,    -6,    -9,    10,     5,     3,   -23,    -2,   -37,    13,   -16,     2,   -11,   -38,   -13,   -42,   -38,   -38,   -50,   -34,   -19,   -39,     8,   -11,   -20,    -7,   -57,     7,   -19,   -40,   -18,    -1,    20,     6,     9,    46,    -4,     2,    -2,    48,    12,   -34,   -87,   -82,  -117,   -96,   -65,   -48,   -43,    -9,   -33,     1,    -6,     9,   -38,    -4,   -11,   -20,   -17,    -6,     2,    -6,   -26,   -24,    55,    27,    44,    19,    14,   -31,  -115,   -83,   -98,   -38,   -57,   -82,   -64,   -17,     6,   -27,     6,   -21,    25,    51,    -4,   -40,     2,    10,     5,    -2,   -65,    16,    48,    53,   -15,     7,    28,    27,   -70,  -130,   -76,   -25,   -35,   -51,   -50,   -35,    -5,   -12,    16,     6,   -17,    14,     0,    -4,   -31,    10,    -1,    -8,   -77,    40,    47,     6,    65,   -31,   -11,    10,   -36,   -31,   -67,    -4,   -40,   -95,   -78,   -65,   -55,    18,    50,     9,    -2,    -8,   -21,   -28,    -6,    -5,     3,   -19,   -13,    26,    38,    22,     5,   -15,   -23,    25,    50,    23,    18,   -23,  -104,  -131,   -72,   -91,   -44,   -17,   -10,   -15,     7,   -30,   -31,   -52,     7,    -1,     2,   -11,    24,   -34,    37,    59,    38,    11,    12,   -18,   -14,     3,   -37,   -59,   -84,  -103,   -45,   -19,    -8,    47,    26,    23,    12,    12,   -26,   -37,   -15,     0,     0,     6,    10,     4,    33,    -9,    10,     9,   -18,   -14,   -11,    23,   -16,   -16,   -40,    -2,    32,   -42,     2,    23,    37,    40,     2,     4,   -27,    -4,   -13,    -2,     6,    -6,    11,    54,    66,   -26,    -3,   -24,   -48,   -38,     9,    20,   -10,    -5,    -1,    13,    20,     9,    -7,    19,    25,   -22,    -8,    11,   -34,    -9,    -7,     6,   -15,     0,    48,    71,    14,    42,    12,   -41,   -13,   -29,    -6,   -30,   -14,    33,    33,   -24,    -3,    -2,    -5,    -1,    30,    42,   -11,   -13,   -11,     1,    22,     0,    -2,    -9,   -11,    12,    34,    35,    52,    37,   -10,    10,   -15,    -5,     0,    14,    12,    15,    17,    -1,   -17,     6,   -10,    18,    11,   -31,     2,    -1,    13,     1,    -9,    -8,   -48,   -48,    10,   -20,   -33,     2,    -3,    13,     5,    35,     2,   -12,    26,     0,    37,     6,     0,   -43,   -43,   -19,   -17,   -74,     3,   -17,     2,     6,   -10,    -3,   -13,   -26,     3,    20,    17,    -9,    39,    49,    10,    17,    35,   -29,    19,   -10,    38,    24,    37,   -42,   -49,   -49,   -22,    18,    18,     2,    -8,    -8,    -5,     4,    -5,    -4,   -16,   -11,   -11,   -18,    -3,   -12,   -48,   -36,   -33,   -50,   -78,   -88,   -90,  -114,   -74,   -57,   -69,   -38,    -5,   -20,    -8,     9,     7,     8,    -9,    -7,    -6,   -11,   -19,   -24,   -18,     6,   -25,   -20,   -26,   -12,   -53,   -44,   -80,   -57,   -47,   -66,   -69,   -52,   -61,   -37,   -42,     9,   -10,    -6,    -8,     3,     0,     5,    -6,    -9,    -7,    -6,     6,    -8,    -4,    -4,    -2,   -12,     7,    -4,    -5,     0,   -13,    -9,   -10,   -10,   -40,   -34,   -44,    -9,    10,     8,    -9),
		    51 => (   -9,   -10,    -4,    -6,    -3,    10,     4,    -2,     3,     5,     4,     1,     5,    -7,     1,     0,    -1,    -3,     1,     2,     7,     2,     6,    -5,     9,    -6,    -9,    -3,    -9,     0,     9,    -6,    -6,     1,     7,   -10,    -9,   -10,    -7,    -5,     1,    -8,    15,     8,    -8,    -5,   -13,     6,     0,    -4,     5,     1,     5,    -3,    -6,    -4,     1,    -4,    -3,     2,     2,    -6,    -8,    -6,   -17,   -30,   -60,   -54,   -38,    12,   -42,   -14,    57,    15,   -57,   -57,   -16,   -35,   -29,   -17,    -8,     8,     1,    -8,    -3,    -3,    91,    52,     1,   -40,   -25,    -8,   -24,   -30,   -53,   -78,   -43,    -8,   -34,   -49,   -18,   -26,   -12,    72,    60,   -54,   -10,   -29,   -11,    -7,    10,    -8,     2,     3,    80,    83,    -6,   -43,   -26,   -19,   -22,   -56,   -70,   -26,    -7,    43,    40,     0,   -46,   -71,    38,    15,    22,   -22,   -10,   -18,     1,   -11,   -34,   -32,    -6,     1,    77,    41,    13,    -7,    -4,   -34,   -89,  -100,   -22,     7,   -26,    20,     6,     6,    27,   -57,   -29,   -17,   -45,   -31,   -19,    -6,   -10,    -9,   -30,   -32,     0,    -3,   -30,     9,     3,   -16,   -34,    -6,   -83,  -107,   -54,     1,    14,    52,    18,   -31,     7,   -65,   -19,   -63,   -57,   -15,    -8,     7,    -1,     1,   -24,   -25,     3,   -10,   -35,     9,    -5,   -44,   -52,   -19,  -117,   -71,     3,    18,    35,    53,    14,   -15,   -38,   -50,   -22,  -112,   -48,   -28,     2,    -7,    -4,   -15,   -64,   -30,     5,   -13,   -32,    13,   -18,   -31,   -47,   -43,  -113,   -55,     4,     0,    10,    37,    63,    38,   -48,   -42,   -29,  -111,   -32,   -26,    24,     1,    -9,    -5,   -40,   -13,     5,   -15,   -37,   -16,   -13,     4,   -27,   -21,   -58,    -2,    21,   -11,   -52,     1,    69,    53,   -42,   -77,     1,     8,   -43,    -5,    18,    -6,   -33,   -20,   -34,   -54,    -1,   -14,   -16,   -14,   -30,   -10,   -57,   -26,   -23,   -54,    47,    -5,   -21,    25,    36,    -7,   -22,   -61,   -47,    -3,   -17,   -77,     8,    29,   -44,   -21,    11,    47,     2,     8,    -5,   -15,   -13,   -31,   -69,   -38,   -65,   -43,   -12,    25,   -22,     5,    55,   -14,     0,   -38,   -60,   -22,    30,    -8,    25,    31,   -39,   -25,   -20,    80,     9,     0,   -75,    30,     2,    -3,   -24,   -25,   -19,    46,    14,    -8,    12,     5,    32,   -23,    -7,   -67,   -73,   -37,    61,     6,    11,    38,   -44,     6,     5,    61,     5,    -6,   -73,     4,     5,   -11,    -7,    16,    49,    30,   -76,    14,    16,   -33,   -21,   -27,   -12,   -40,   -49,    19,    69,   -26,   -33,   -59,   -48,    43,    33,   -10,    -2,     1,    -5,     8,    -7,   -39,     3,    25,   -18,   -27,   -67,   -44,    17,    -4,   -10,   -31,     8,     3,     0,     6,    18,   -28,   -55,    -8,    -6,   -13,    50,     9,    -7,     0,     8,    26,    -1,   -46,   -38,    -1,   -17,   -29,   -27,    60,    35,    49,    19,   -51,     2,    -7,    35,   -17,    43,   -19,   -48,   -15,   -47,   -28,     5,   -26,     2,    -5,     9,   -29,    -4,   -25,   -16,     2,   -17,   -38,   -23,    30,    16,    -2,    14,   -37,   -36,    -9,    13,   -39,     7,   -23,   -35,   -37,    -1,   -43,     1,   -13,    -5,    10,     3,   -14,   -12,   -47,   -34,   -48,   -15,   -29,   -31,   -20,    10,     8,     8,   -20,   -28,   -40,    10,   -42,   -52,   -33,    21,    22,   -25,   -42,   -12,    10,    -7,     2,   -11,    -9,   -25,    -2,   -34,   -18,   -47,   -30,  -100,   -21,   -33,    58,    28,    -4,     7,   -12,    28,   -65,    19,    -9,   -55,   -50,   -49,     4,    -1,    41,    -8,    -6,     7,    -9,   -10,    -4,   -12,   -30,    18,   -53,   -52,   -20,   -11,    26,    50,    26,    -1,   -36,   -21,   -85,   -26,   -28,   -72,   -45,   -20,    25,    31,    46,    10,     9,     0,   -27,   -26,   -15,   -30,   -61,   -16,   -21,   -16,   -11,    44,    15,    21,    17,     6,   -14,   -21,   -37,     2,   -60,   -93,   -34,    -1,    -9,    45,    -7,    17,    13,     6,   -23,   -25,   -11,   -42,   -91,    -5,    -1,   -26,     1,     4,     7,   -10,     3,   -16,   -57,    41,   -15,    18,   -20,   -69,   -61,   -28,    15,   -17,    -4,    23,    10,     8,     8,   -17,   -12,   -17,   -74,     6,    -4,   -13,   -33,   -24,    -6,     7,   -14,   -16,   -22,    22,     9,    37,    -5,   -57,   -24,   -49,    40,    31,    -2,     6,     1,   -11,   -26,    -9,     9,    37,   -26,    10,    58,     4,    33,    -9,     3,    -2,     4,    12,    57,    47,    15,    32,   -21,   -11,   -32,   -36,   -10,    75,     7,    -8,    -7,    -7,   -13,   -11,    -9,    48,     8,    -7,     9,    42,    58,    -9,   -51,   -48,   -67,   -87,   -33,   -65,   -41,   -38,   -22,   -60,    -5,   -36,    50,    42,     8,     7,    -2,    -8,     1,    -5,    -7,    -3,    -9,   -14,   -29,  -127,  -103,   -72,   -62,   -17,   -80,   -76,   -85,   -70,   -73,  -120,   -46,   -36,   -34,    -2,    -4,    -9,     5,     7,    -9,    -4,    -3,   -29,   -59,   -43,   -38,   -37,   -32,   -26,   -36,   -60,   -63,   -67,   -64,   -47,   -47,   -12,   -27,    -5,   -31,    -3,    -3,    -6,     4,    -2,     3,    -8,    -3,     9,     0,    -9,     7,     1,     2,    -7,    10,    -5,    -6,    -3,    -7,   -14,   -10,    -2,     2,     6,    -6,     1,     3,     2,     1,    -7,    -9,    -6,   -10),
		    52 => (    3,     6,    -6,    -8,     5,     2,   -10,     7,    -5,     0,     7,    10,   -14,   -12,     8,    18,     3,     8,     8,    -3,     2,    -8,     6,    -7,     2,    10,     4,    -3,     3,    -3,     8,   -10,     9,     9,    -9,    -6,    -5,     6,     8,    -6,     6,     8,   -19,   -14,    10,    14,    -6,   -42,   -21,    -3,     2,     5,     6,     6,     4,    10,    -5,    -2,   -14,   -15,   -14,     9,   -12,   -18,    39,    60,    71,    36,    30,   -20,     0,   -27,   -72,   -54,    -2,    19,     2,    20,   -21,    15,    30,    18,    -8,     2,    -8,    -6,   -16,   -60,   -49,   -55,   -17,   -29,    20,    21,    -9,   -10,   -23,    13,    27,   -13,    -4,    -7,   -12,    48,   -15,   -11,   -17,   -73,   -38,    17,   -19,     1,     0,    -6,   -10,   -17,    44,   -11,    -8,     8,     1,    11,   -18,     1,    28,    11,    -4,    20,   -31,    17,   -37,   -13,    25,   -38,   -20,   -66,   -71,    31,   -53,   -24,    -6,    -7,     1,   -23,     8,   -58,   -63,   -85,   -41,    -7,    42,     5,   -29,    24,    14,    11,   -25,    12,    -9,    -2,    -1,    13,    -4,    34,   -58,    59,   -43,    -6,    -6,     1,     2,    60,    47,   -51,   -40,   -21,    19,    39,    39,     3,     6,    46,    10,    -1,   -18,    10,     4,    -7,   -16,   -42,   -15,    -9,     5,   -46,   -46,    -6,     2,     0,   -15,    77,    58,    41,   -15,     9,   -13,     3,   -10,    18,    13,    24,     6,    30,    36,    33,    11,    28,   -17,   -29,    49,     6,   -40,   -47,   -38,   -32,   -28,    56,    -9,    56,    37,    31,   -41,   -16,   -19,    30,     2,    -8,   -15,   -29,   -12,     7,    29,    42,    -7,    48,   -34,    -1,    45,    41,  -110,   -68,   -47,   -34,    10,   -19,    16,    12,   -17,    11,   -27,   -29,   -14,    39,   -39,     4,    22,   -54,   -16,     9,    23,    13,    -9,    47,     2,   -27,   -29,    42,   -90,   -58,   -28,   -13,     1,    -2,     5,    32,   -62,    68,    35,    -5,   -14,     3,   -36,   -45,    -2,    25,   -16,   -17,   -13,   -21,    -6,    12,    25,    -6,   -21,    43,   -19,   -21,     9,   -12,     2,   -29,    -8,    41,     8,    15,    33,     3,   -16,   -40,   -87,    -2,   -29,   -50,   -60,   -49,     3,   -18,   -47,    -9,   -23,    -4,   -22,    20,    -7,     3,   -45,    -9,    -7,     0,   -56,    -4,    12,   -61,   -24,   -45,   -56,   -41,   -49,   -47,   -18,   -76,   -94,   -24,     1,   -10,   -52,   -11,   -34,   -16,    -9,   -29,   -13,    23,    -4,   -24,    -2,     6,     4,    -7,   -10,   -23,   -86,   -76,  -128,   -76,   -58,   -73,   -96,   -55,   -43,   -22,   -17,   -41,   -36,   -45,   -37,   -42,    16,   -34,    -9,    25,    42,   -22,     7,   -30,   -38,   -14,   -50,   -91,   -99,  -102,  -159,  -101,   -52,   -54,   -17,   -30,     1,   -21,   -57,   -20,   -19,   -17,   -44,   -69,    -8,   -78,    -8,     3,    53,    28,     8,   -26,    -6,   -23,   -96,   -52,   -46,   -67,    12,    -6,   -24,    25,    -1,    32,    10,   -49,     7,    -8,   -59,   -68,   -67,   -40,   -74,   -39,    18,   -23,    60,    84,     1,    -2,   -37,   -61,  -109,   -38,   -44,   -31,   -16,    17,    20,    21,   -35,    14,    18,   -21,   -31,   -13,   -29,   -62,   -43,   -17,    28,   -23,    25,    58,    77,    51,    -8,    -6,     3,   -43,   -37,   -47,    -5,   -13,    -3,     4,    24,    10,   -34,    57,    36,     1,    -9,   -14,    -8,   -54,   -33,   -18,   -15,   -19,   -42,    99,    57,    47,    -6,    -7,   -15,   -84,   -29,   -23,    27,    39,   -16,   -25,     7,    -3,    18,    -6,    -8,   -12,    -8,    25,   -31,   -40,   -50,    31,    39,    38,    73,   120,    -7,    63,    -5,   -18,    17,   -42,   -50,   -17,    39,    25,   -26,   -39,    19,    11,     4,    75,    66,    19,    32,    -7,   -15,   -31,     5,    40,    17,    36,   -11,    34,    31,    65,     3,    -9,    38,    -5,    -5,   -26,    91,    30,    22,    28,    63,    53,    38,   103,    36,    28,    57,    -6,   -11,    -9,    62,    57,    23,    17,    12,    48,    22,     1,     7,    20,    20,    48,    16,    13,    46,    30,   -12,    26,    21,    24,     3,    77,    61,    47,    30,    40,    19,    29,    34,    27,    47,   101,    47,    47,    46,   -13,     5,    -3,    -2,     0,    -6,    50,    70,    37,     9,    41,    10,    16,    10,     6,    25,    20,   -19,   -44,    -3,   -42,    16,    44,    75,    88,    71,    -6,   -66,   -21,    -8,    -8,     7,   -47,   -25,    14,    52,    28,    20,    46,    19,    66,    49,    35,    12,   -13,   -42,   -27,   -30,    -1,    36,    52,    93,    65,    52,     8,   -34,     3,     4,    -1,   -51,   -35,   -12,   -29,     3,    28,    69,   -21,     6,     5,    45,   -22,    29,    13,   -49,   -15,    -2,     1,   -56,   -30,    -5,    53,   105,    59,    33,     3,     7,    -2,   -33,    -4,   -42,  -102,    47,   -15,   -53,  -103,  -134,   -40,   -20,    -9,    45,    33,   -33,    12,   -69,   -89,    -8,    14,   -74,   -33,    18,    55,    38,    -4,     6,    -8,    -6,    -2,   -34,   -62,   -70,   -46,   -44,   -66,  -115,   -93,   -54,   -59,   -60,   -37,   -89,   -83,   -66,    -6,   -29,   -38,   -23,     3,    -9,    -1,    -9,     6,   -10,     8,    -8,     5,    -5,     0,   -12,     1,     8,    -2,   -31,   -51,    -4,   -21,    -5,    -2,     2,   -11,    -6,     4,   -19,   -34,   -17,    -4,    -5,     2,     0,    -1),
		    53 => (   -3,    -4,     2,    -5,    -3,    -6,    10,   -10,     6,     2,     2,    -7,   -10,    -9,    -3,    -2,    -6,    -4,    -4,    -4,     9,    -7,    -8,    -3,     6,    -4,     0,     1,    -5,    -1,     7,     1,    -5,    -3,     6,    -5,     9,   -10,     2,    -3,    -8,    -7,   -19,    -5,   -23,   -10,     1,    -6,     0,     1,     9,     3,     8,    10,     2,    -9,     7,     9,     3,    -7,     3,     6,     6,     1,   -39,   -47,    33,    41,    28,   -18,   -39,   -40,   -58,   -60,   -41,   -20,    -8,   -28,   -32,   -44,   -13,    -9,    -3,     0,    -6,     1,    -3,   -23,   -10,    -2,   -14,    19,     9,   -11,    31,    33,    23,    25,     6,   -25,    14,    32,    38,   -17,   -15,   -23,    -9,   -73,   -33,    -8,    -3,     1,    -7,    18,     5,     0,   -13,     9,    10,    26,    12,   -10,   -18,   -32,   -45,   -49,     0,   -21,   -24,   -61,   -28,     2,   -39,   -32,    39,   -81,   -67,   -36,   -11,    -3,     0,     5,     9,   -15,    -8,    28,    39,    66,     6,   -45,   -65,   -31,   -23,   -28,    -1,   -11,    -8,    -9,   -11,    10,   -10,   -27,   -38,   -30,   -30,    -9,   -29,    -9,     1,    14,    -2,    18,     6,    -1,     7,    -9,   -53,   -38,    31,    -9,     4,   -18,   -29,   -19,    -9,    -1,     1,   -41,   -33,   -15,   -14,   -11,   -12,   -63,   -36,   -14,     9,    19,    27,   -39,   -90,   -37,     2,   -28,   -46,   -19,   -18,     7,   -16,    -1,     6,     5,   -10,    21,    -4,   -41,    10,   -26,    -6,   -35,   -22,   -50,   -37,   -16,     1,   -10,    24,   -55,   -75,     1,   -25,   -40,   -23,    15,    15,   -10,     3,   -30,     7,   -23,     5,     3,    34,     9,    17,    53,    31,   -70,  -118,   -38,   -51,     1,    -7,   -46,   -38,   -43,     8,     4,    27,    -5,   -14,   -17,    23,    37,    55,    29,    25,   -17,   -28,   -19,   -31,   -20,    35,    22,    22,   -55,  -141,   -56,   -57,    -9,    -1,   -48,   -22,    32,    15,    12,    60,     5,    82,    38,    44,    35,    -1,    -3,    -9,   -25,   -70,    -5,    30,    32,    22,   -10,    27,   -17,  -130,   -13,   -41,     4,    -5,   -50,   -22,    74,    67,    63,    15,    40,    24,    55,    21,   -39,   -83,   -80,   -68,    23,    16,    21,    34,    42,    65,    12,    15,    -4,   -78,   -73,   -16,   -10,    -4,   -50,   -44,    75,    43,    30,     1,    17,   -49,   -46,   -63,  -142,  -104,   -23,    35,    62,    22,     8,    31,    -3,   -14,   -34,   -22,   -48,     1,     7,     1,     7,     5,   -33,   -94,    32,   -48,   -32,   -24,   -30,   -65,  -133,  -137,   -87,   -18,    23,    47,    10,    12,    -6,   -28,   -36,   -25,   -14,   -71,   -54,    43,   -25,   -23,    -7,   -16,    14,   -15,   -25,   -63,   -76,  -110,  -101,   -99,   -51,   -22,   -39,    22,    35,    19,    15,   -11,    10,   -51,   -33,   -43,   -31,   -76,   -15,    63,   -17,   -36,   -23,    -5,    33,    15,     8,   -22,   -39,   -84,  -111,   -82,    -4,    21,   -17,    26,    54,    88,    -1,    29,   -11,   -13,    -4,   -17,     3,   -37,   -20,    49,   -20,    44,     8,    -1,     8,    24,    48,    11,   -31,   -45,   -31,   -66,   -44,   -47,   -91,   -11,     8,   -17,   -43,    29,    21,   -27,     5,     6,    57,   -13,   -41,    28,   -52,    18,     3,    -2,     5,    11,    11,     4,    -5,   -18,   -43,   -85,  -110,  -137,  -151,  -184,  -149,   -95,   -58,    36,   -10,   -46,    34,    28,    55,    18,   -38,   -16,   -68,    -9,    -3,   -19,     7,    57,    15,    71,     6,   -32,     0,   -13,   -72,   -66,  -100,  -144,  -111,   -68,   -64,    -5,    45,    33,    36,    12,    -9,    24,   -16,   -89,   -25,     5,   -23,    -2,   -29,   -36,   -31,    18,    30,    -2,     1,   -24,    19,   -10,   -32,   -24,     1,     3,   -20,   -18,     3,   -22,     0,     9,     3,    42,    -1,   -28,    16,   -13,   -21,     6,    -7,   -35,    -5,    18,    33,    38,    27,     8,    45,    39,    56,    24,     1,   -18,   -53,   -21,   -38,   -31,     8,    38,    -7,    13,   -32,   -42,   -29,    -8,   -10,    -6,    22,   -16,     2,   -15,    21,    10,    39,    45,    14,     3,     1,     7,   -19,     3,   -38,   -36,   -54,   -13,    17,    26,     0,   -21,   -29,   -47,   -20,   -18,    -1,   -10,     6,   -25,     5,     6,   -13,   -24,   -33,    -5,    -8,     9,     6,    13,    13,    17,   -10,    -5,     4,    -5,    35,    -4,     8,   -54,   -50,   -43,   -21,   -14,     7,     2,     4,    28,    40,    45,    30,   -12,   -19,   -13,    -9,   -50,   -20,   -37,   -14,   -17,    29,     7,    26,    29,     1,    13,    22,   -55,   -44,    39,    24,     2,     2,    -5,    -5,    -2,    33,    40,     0,   -36,   -19,     6,    26,     2,     8,    22,     5,     4,   -18,    36,    33,   -20,   -56,   -14,   -18,   -40,   -64,   -41,   -25,   -12,     0,    -2,     8,     2,   -43,   -34,    13,    24,    14,   -23,   -21,   -72,   -61,   -48,   -91,   -60,    -3,    -2,   -48,   -48,   -49,   -27,   -33,   -30,   -56,    -2,     1,     6,     2,    -6,    -1,     2,   -31,   -75,   -70,   -51,   -57,   -76,   -67,   -96,   -82,   -70,   -36,   -26,   -29,   -41,   -99,   -91,   -77,    -4,   -32,    -8,    -2,     6,     4,    -1,     3,    -3,    -6,    -6,    -9,    -6,   -15,   -13,   -18,   -15,   -48,   -36,   -44,     0,   -33,   -31,   -41,   -32,   -33,   -31,   -45,   -20,   -11,    -7,    -2,    -5,    -3,     9,     3),
		    54 => (   -4,    -5,    -5,     7,     3,    -5,     5,    -1,    -3,   -10,     4,     1,   -12,   -12,   -12,    -9,     7,   -10,    -9,    -2,    -9,   -10,     3,    -7,    -9,    -6,     4,     7,    -3,     9,     6,     8,     8,    -4,   -42,   -35,   -10,     2,   -19,    -2,   -17,    12,    38,    -9,    -9,    -5,    -9,    -5,   -21,   -14,   -13,    -8,    -9,    10,    -1,    -1,    -9,    -2,    -5,   -17,   -59,    -4,   -26,   -42,   -63,   -21,   -14,   -10,   -19,   -40,   -32,   -55,   -75,   -30,   -19,    -9,   -48,   -40,    -4,   -12,    -8,   -29,    -2,     1,     1,     1,   -18,   -27,   -47,   -16,   -34,   -45,   -20,    -9,   -22,   -12,     5,   -22,   -39,    -6,     7,    29,   -36,   -26,   -36,   -13,   -22,     1,    -6,   -19,     4,     1,     6,     2,   -16,   -11,   -19,   -28,   -47,    26,    60,    31,   -24,   -74,   -94,   -59,   -49,   -45,   -80,   -99,  -103,   -66,   -30,   -23,     8,    84,    62,    38,   -74,   -14,    -8,    -8,   -22,     8,   -27,    -2,   -25,    21,    87,    25,   -54,   -94,   -64,   -37,    94,    54,    39,   -17,   -96,  -118,   -42,   -39,    -7,    26,    16,   -26,   -12,   -11,     3,     5,    -9,   -35,    36,    49,   -18,    36,    38,   -38,  -109,  -127,   -21,    13,    16,    45,    40,    12,   -91,  -175,  -158,   -17,    53,    56,    35,   -81,    20,   -57,    -3,   -32,     2,   -36,    24,    38,    19,    27,    -8,   -20,   -61,   -39,   -58,    -5,    45,    45,    29,    26,  -132,  -183,   -84,    23,    77,    84,     8,   -99,     6,   -70,   -21,   -32,    -4,   -44,    -3,    45,    28,    33,   -12,   -14,   -43,   -60,   -76,     6,    32,    71,   -25,   -89,  -163,   -85,   -13,    41,    24,   -11,    -7,   -35,    20,   -50,    -6,   -13,   -16,   -49,    14,     3,    28,    65,     1,   -30,   -40,   -76,   -28,    -2,    55,    30,   -14,   -86,   -81,   -34,    29,    31,   -13,    15,   -12,   -23,    21,   -44,     4,   -18,   -45,   -52,   -19,     1,    12,     8,   -50,    16,   -15,   -62,    23,    -4,    48,    15,   -13,   -51,   -53,    -2,    20,    -3,     5,   -32,     8,    24,    -9,   -39,    -8,     4,   -44,   -26,   -38,    18,   -12,   -16,     7,    27,    -4,    13,    15,   -47,     4,     4,   -28,   -53,   -37,   -12,    -1,     6,    14,    -1,   -36,    -3,   -30,   -69,     2,    -3,   -30,  -106,   -32,    24,   -18,     4,    13,    10,    27,   -41,    13,    11,    -7,   -27,   -33,   -29,   -50,     8,    20,    10,     8,   -44,    -8,   -30,   -79,   -58,    -4,    10,   -33,   -72,   -48,    -8,    -1,    19,    -3,    23,    62,     2,   -45,    28,   -44,   -32,    20,     1,   -13,    25,     3,     5,     2,   -11,   -47,   -64,   -74,    -4,     7,    -3,   -31,   -65,   -19,     1,    36,     3,     3,    22,    32,     5,     2,    35,    18,   -20,    -2,    31,   -16,     2,    10,    24,    25,   -27,    -2,   -43,   -19,     5,    -7,    -5,     0,   -63,    -6,    10,    19,    51,    40,    32,    29,    21,    23,    -2,    15,    -8,   -32,     8,     7,     8,   -19,   -24,     8,     0,   -25,   -30,   -13,    14,     8,    -4,    -8,   -49,   -29,    16,    47,    56,    27,     0,   -27,   -12,    -3,    -7,     3,    41,    19,     7,   -11,     3,    19,   -18,   -41,   -38,   -13,   -24,   -56,   -19,    -4,     3,   -16,   -29,   -17,     4,    15,     3,    31,   -23,    -2,   -23,     3,    -7,    37,    14,    10,   -14,   -22,   -25,   -24,   -13,    -6,   -26,   -54,   -49,   -30,   -23,   -28,    -7,    -3,    43,    36,   -13,   -32,   -38,   -26,    13,   -65,   -62,   -33,     6,    34,    -9,   -19,   -25,   -18,   -42,   -69,   -30,   -35,   -41,   -23,   -37,   -14,   -25,   -10,   -23,   -26,    62,    18,   -89,   -62,   -33,   -17,    -9,   -89,   -52,   -31,   -48,     3,   -10,   -22,   -17,    21,   -31,   -55,   -60,   -51,   -55,    -4,   -30,   -18,   -19,    -1,     0,     0,   -27,    -2,   -28,   -27,   -34,   -54,    13,   -41,    -6,     2,   -45,    41,     4,   -25,    -2,    38,   -38,   -89,     4,   -21,   -15,    28,   -43,   -11,     7,     3,    -3,   -21,   -80,   -43,     5,   -45,   -59,    13,    18,    -5,    10,   -14,   -76,    -1,   -24,    -8,   -21,    10,   -12,   -64,    -7,   -22,    10,     7,   -51,   -25,     3,     2,    -5,     7,   -46,   -45,     9,   -10,    18,    33,   -32,   -12,    -4,   -23,   -42,   -16,   -25,     8,   -28,     7,    43,   -13,     5,    24,   -11,    29,     5,     7,     7,   -10,     0,     1,   -26,   -35,   -69,   -20,    15,    16,     2,    57,    26,    15,   -45,   -32,   -49,   -46,   -35,     4,    15,    30,    -7,   -24,     1,    18,    28,     0,     4,    -3,    -8,     3,     0,   -58,   -52,    22,    17,    14,     9,     7,    50,    37,   -32,   -10,    -7,   -75,     1,    16,    19,    40,     5,    38,    19,    -5,    52,     5,    -4,     6,    -2,   -10,    -8,   -39,   -84,    15,     0,    -4,    -5,    27,    30,   -74,  -107,   -33,     4,   -64,    15,   -39,   -63,     3,     5,    33,     3,    -9,   -17,    -3,     6,     5,    -4,     8,   -44,   -13,   -46,   -55,   -23,   -33,   -41,   -60,   -43,   -52,   -69,   -16,     4,   -14,    13,   -52,   -67,   -69,   -79,   -58,    -4,    -8,     5,     2,    10,    -3,     3,     3,     5,    -4,    -8,   -19,   -26,   -27,   -18,   -48,   -39,   -31,   -36,   -63,    -8,   -30,   -51,   -44,   -38,   -52,   -34,   -41,    -7,     0,    -1,     3,     1),
		    55 => (   -8,     0,     5,    -3,    -1,     7,     1,     7,    -5,    -8,     6,    -3,     2,   -14,     6,     6,     8,    -8,     2,     0,    10,     4,     9,    -2,    -1,    -6,     3,     4,    -3,    -1,    -8,     1,    -1,     0,    -1,   -13,     3,     0,    -6,   -32,   -17,   -12,   -39,   -49,   -45,   -51,   -36,   -42,   -59,   -57,   -20,    -5,    -2,     6,    -4,     1,    -6,    -7,   -31,   -31,   -14,   -16,   -31,   -29,   -50,   -79,   -71,   -83,  -100,  -127,   -64,    20,    26,    38,    19,   -16,    -4,   -45,   -47,   -11,   -42,   -31,     8,    -4,     5,     6,   -15,    -1,   -13,   -48,   -92,   -59,  -120,    25,    46,    -7,    15,     1,   -31,   -56,   -47,    -2,    28,    58,    -7,    47,     1,   -43,   -23,    26,    78,     0,    -6,   -22,   -40,     1,   -52,    -9,    -3,    11,     1,   -11,    18,    -5,    18,   -26,   -12,   -32,   -51,   -31,    34,   -46,   -42,    -8,   -25,   -22,    78,    53,    12,   -25,    -4,     6,   -40,     0,   -40,   -13,   -33,     6,   -29,     2,    -1,    69,    55,   -18,    22,    44,    -6,   -37,   -91,   -17,    -7,    -1,     8,    38,    -1,    49,    17,    -5,     9,    -1,    -4,   -57,   -58,   -29,     2,    25,    24,    -6,    -1,    49,    68,     9,     8,   -25,   -35,   -45,   -47,    -7,   -18,   -15,    16,    64,    63,    77,    -8,     9,     7,   -33,     7,   -95,   -86,   -37,    27,    63,    55,    47,    50,    19,    -8,     8,    27,    -2,    37,    12,   -52,   -14,    14,     1,     5,    -1,    17,    17,   -20,    35,    -9,   -26,   -73,  -123,   -62,    39,    -2,   -45,   -10,    17,    19,    -4,    -4,     6,    36,    38,    -6,    26,   -43,   -81,   -22,   -22,     7,    -3,    88,    33,   -64,    18,     1,    -8,   -56,   -89,   -34,    35,    19,   -53,    11,   -26,     6,    66,    40,    60,    86,    53,     6,   -24,   -87,   -95,   -95,   -48,    16,    -2,    49,    53,   -33,   -24,    -1,    -4,   -71,  -148,    54,    58,    35,    18,   -26,   -19,    30,    53,    97,    68,    64,    72,     3,   -90,   -46,   -63,   -61,   -37,  -124,  -105,    39,    57,    52,   -32,     6,   -15,    -6,   -32,    15,    32,    23,   -11,   -17,   -22,    -2,    21,    43,    47,    18,    52,    23,    -9,   -30,   -77,   -44,   -35,  -126,  -142,    -6,    -7,    23,    10,    -6,    -7,   -12,   -21,    40,    16,    -2,     6,     1,    -5,     1,   -45,     8,     8,    -8,    10,   -29,   -34,     0,   -18,   -52,   -15,   -91,   -60,  -140,   -59,    54,   -59,     1,    -4,   -25,    -6,    -1,    32,   -23,     1,    -7,    -6,    -1,    21,     7,     7,    -9,    13,   -17,   -47,    -3,    24,     6,     7,   -21,   -74,  -114,   -87,     1,   -40,    10,    -9,   -10,     7,   -59,    -9,   -18,   -12,   -27,    -7,    -6,   -23,    -2,   -35,     9,   -26,    28,    -6,   -25,     8,    26,    -9,     1,    67,     5,   -56,   -34,   -22,     2,     5,   -30,   -21,     8,     0,    -6,    -9,   -71,   -47,    11,    -5,     6,   -24,    -5,     2,   -15,    -8,     5,   -24,   -36,   -73,    -3,    64,    29,   -56,   -54,   -61,     3,   -19,   -69,    60,     6,    21,   -83,  -122,   -58,   -64,   -31,    54,    -7,    -9,   -14,   -38,   -15,   -38,     0,    20,   -22,   -24,    -6,    28,   -20,  -122,   -71,   -68,    -3,   -14,  -106,   107,    23,     2,   -25,  -110,   -75,   -58,   -25,    -6,   -40,   -26,   -28,   -24,    14,    37,    12,    43,     1,    -2,    10,    23,   -68,  -122,   -98,  -100,   -13,     9,   -72,   105,   102,    58,    -7,   -62,   -87,  -121,   -17,   -52,   -31,   -50,    -3,    -6,    24,    29,    -9,   -23,    20,    31,    33,    56,    -7,   -18,  -107,   -33,    -1,   -28,    56,     6,    82,    77,    22,   -41,   -17,   -68,   -29,   -35,    -9,    -8,     1,    27,   -22,    18,    57,    -1,    65,     3,    40,    58,    63,    36,   -66,   -72,    -9,   -28,    44,   -11,    36,    42,     8,     1,     4,   -12,   -42,     1,    -7,    31,   -10,   -20,    30,    44,     6,   -37,    30,   -11,    78,    34,    33,    60,   -58,    -2,    -7,   -10,   -52,   -97,    -6,    36,   -21,   -34,    38,    36,    -2,   -16,   -21,    -4,    18,    49,    44,    22,    44,    41,    11,    45,    -8,    51,    20,    86,    30,   -12,   -12,    -5,   -79,   -32,   -61,   -55,   -32,     7,    11,    21,    24,   -10,     0,    14,   -12,     2,    15,     0,    12,    40,   -27,     0,    -2,    88,    92,   110,    71,     1,     5,     7,    14,    18,   -28,   -18,     7,   -13,   -48,     4,   -13,    -7,   -21,    16,    17,    -9,    16,    14,    35,    36,   -15,    17,   -25,    64,    62,    76,    51,    -3,    10,    -6,   -50,   -14,   -40,   -25,   -32,    20,    26,    69,    49,    42,   -12,   -29,   -53,    11,   -14,    49,    39,    52,    19,   -28,    15,    -1,    73,   -48,   -28,     3,     9,     1,     1,    37,   -76,   -95,   -33,   -15,    14,   -33,   -48,   -47,     2,   -27,   -59,     0,    54,    74,    67,    48,    11,    53,    84,    71,    71,   -27,   -10,    -6,     9,     7,   -10,   -21,   -33,   -72,   -94,   -87,   -33,    -7,    20,    15,     0,   -17,   -78,    26,   -14,    22,    20,    79,    21,    -2,   -19,   -39,   -23,     8,     8,     5,    -4,    10,     9,    -2,   -17,   -16,    -7,   -18,   -19,   -22,     9,    10,    12,     6,   -99,   -74,   -22,   -33,   -23,   -45,   -55,   -63,   -35,    -6,     6,     8,     4,     2),
		    56 => (   -1,    -4,    -1,    -4,     5,    -5,     8,    -3,    -6,     3,     0,   -10,    16,    22,    -6,     9,    -8,     8,     4,     1,     9,     4,     5,     2,     0,     2,     5,    -5,     7,     2,    -1,    -9,   -10,    -9,    22,    25,    47,    28,    22,    16,     7,    33,    -5,   -14,   -10,    -7,     1,     9,    58,    29,    19,     4,    -3,    -4,    -1,    -3,     0,    -4,    -4,    -3,    30,     1,    17,    51,    44,    39,    25,   -15,   -22,   -26,   -23,   -10,     1,    -6,    -6,    26,    32,    43,    33,    53,    21,    20,    -7,    -6,    -6,    -8,   -45,   -46,    -9,    34,    30,    23,    16,    27,    -8,   -35,   -47,   -92,   -41,   -22,    -5,   -39,    18,    56,    32,    22,    12,    52,    37,     7,    -4,     3,    10,     1,   -53,   -58,    41,    55,    35,     7,   -20,    18,     6,   -49,   -63,   -94,   -61,    -5,   -14,   -27,   -61,     4,     5,   -18,   -40,     4,    40,    33,    63,    67,    -8,    10,   -29,   -52,    82,    46,    18,    11,    13,     5,    -1,   -25,   -36,   -69,   -27,    23,   -12,    10,   -26,   -28,   -30,   -12,   -22,    13,    25,    31,    68,    47,    -3,     0,    16,   -11,    61,    18,    33,    12,    68,    28,   -30,   -65,   -68,   -73,   -16,   -20,   -56,   -24,    -3,   -53,   -32,    -4,   -10,    -2,     9,   -39,    15,    80,     1,    -3,     5,   -18,    65,    26,   -12,    36,    29,    39,   -20,   -57,   -78,   -42,     0,   -54,   -67,    -3,    -4,    -9,   -10,   -31,   -35,   -43,   -42,   -16,    29,    69,     0,     4,     5,   -22,    48,    15,   -12,    27,     7,    -5,   -44,   -77,   -85,     2,     7,   -60,   -11,    26,    13,    24,    27,     9,   -34,   -11,   -10,   -23,    30,   -42,    -5,    -5,   -11,   -42,    30,    11,   -16,    25,    -8,   -38,   -82,   -92,   -82,   -28,   -11,   -24,    18,    46,     6,    20,    34,     4,   -14,     6,    -8,   -41,   -13,   -13,    -4,    -6,   -15,   -40,    47,    32,    18,    57,     6,   -41,   -65,   -78,   -62,   -13,    -8,     9,     9,    39,   -34,   -19,   -22,    16,     2,     6,   -19,   -16,     0,    -7,     0,     5,     8,   -12,    38,    36,    26,    13,    -4,   -31,   -49,   -60,   -36,    -5,     8,    -6,   -18,   -70,   -47,   -13,   -30,     0,    18,    25,     7,     4,   -15,   -22,    -9,     3,   -10,   -21,    24,    59,    -3,    13,    -4,   -32,   -48,   -67,   -20,    70,    12,     9,    10,   -26,   -24,   -38,   -17,    20,    39,    33,    26,    -6,    -7,   -43,     8,    10,    -7,   -19,    11,    11,   -10,     2,    16,   -25,   -31,   -74,     2,    38,   -15,   -37,    -5,     3,   -28,   -26,   -17,    17,    16,    31,    26,    -2,    -6,   -10,    -6,    -2,     5,   -27,     6,    12,   -13,    15,     0,    -6,   -41,   -27,    34,    44,   -64,   -45,    -2,     6,    -9,    -9,   -36,   -12,     4,    22,    18,    -3,   -13,   -16,    -9,     0,     4,   -16,    25,     9,   -16,    -6,    -3,    -4,   -35,    -2,     0,    22,   -26,   -10,     5,   -12,    -5,   -37,   -39,     0,    19,    39,    15,    -8,     7,   -63,     6,     5,   -17,    -7,    33,     4,   -28,   -23,   -25,   -18,   -19,   -12,    24,     1,    14,    50,     4,     5,    24,   -41,   -24,    -4,    24,    20,    -8,    11,     0,   -29,     3,     5,    -2,    25,     0,     8,   -14,   -23,   -18,     3,    15,     4,   -17,    26,     1,    10,    55,     1,    20,    -8,   -36,    -3,    -5,    23,     0,    -1,   -11,   -26,     5,     1,    -6,     7,   -17,    10,   -38,   -33,   -33,    -7,    -1,    24,   -22,     9,   -22,    22,    13,     7,    39,    14,    -6,   -17,    16,    26,    -3,    -8,    -1,   -22,    -9,    -8,    -9,    31,     5,    -6,   -41,   -50,   -42,    -3,     3,    -3,   -12,     0,    11,    27,     3,     8,    38,    40,    27,    12,    -2,   -31,   -17,    11,   -43,    -5,     2,   -13,    -7,   -24,   -21,   -28,   -11,   -56,   -50,   -19,     8,   -18,   -18,    14,    11,    29,    17,    40,    36,   -26,     1,   -23,   -57,   -28,   -21,    20,   -15,     0,    -8,     7,    -7,   -23,    -7,   -28,    -3,   -28,   -23,     8,     0,    -2,     1,    32,    14,    18,    12,   -23,   -32,   -18,     2,   -14,   -34,   -27,   -26,   -21,   -11,     4,    -3,    -8,    -2,   -27,     1,   -17,   -40,   -23,     6,    -1,   -18,   -27,    -3,    25,   -18,    12,   -11,   -19,   -54,     5,    -3,   -29,   -42,   -47,   -50,   -17,     0,     8,     2,     8,     2,   -15,   -19,     0,   -15,   -27,   -19,   -21,   -10,   -28,    -2,   -41,   -25,    15,   -28,   -57,   -27,   -23,   -19,    -5,   -28,   -30,   -37,    -2,   -12,    -6,    -3,    -9,   -10,   -10,    -7,   -12,     4,    -3,   -14,    -6,   -29,   -14,    -6,   -10,   -19,    -9,    -5,   -11,   -21,   -45,   -26,   -12,    -6,    -8,    -4,     4,     5,    -9,    -7,     2,   -10,     7,   -10,   -12,   -24,   -16,   -10,   -16,     2,   -11,   -16,   -12,     3,    -1,    -5,     3,     1,   -10,   -35,   -14,    -1,    12,    -8,    -4,    -4,    -2,   -10,     8,     3,     7,    -9,    -1,    -4,    -2,    -9,     5,   -10,     0,    -3,    -2,     5,    -2,     6,    -9,    -5,     3,   -19,   -10,    -6,     3,    -2,     1,     0,    -4,   -10,    -5,     9,   -10,     1,     0,    -4,    -7,    -9,    -5,   -12,    -9,    -4,    -9,    -1,    -7,    -2,    -7,    -7,     5,     6,    -9,     0,     4,    -3,     8,    -7,     3),
		    57 => (   -3,    -9,     7,    -5,    -8,     6,    -7,    -8,    -5,     3,    -4,    -2,     5,    -7,    -6,    -8,     9,    -1,     0,    -4,     1,    -2,    -4,     0,     6,     6,     0,     9,     1,     2,     1,    -4,     6,    -7,     8,     4,    -7,    -4,    -4,   -39,   -43,   -38,   -25,   -84,  -100,  -105,   -22,     3,    -9,     0,    -7,     0,    -7,     2,    -8,     0,    -6,    -5,    -5,    -9,     6,     5,   -19,   -20,   -61,   -62,   -90,   -81,   -49,   -31,   -23,   -54,   -42,   -24,   -30,    -1,   -50,   -44,   -39,   -34,   -31,   -15,     3,     4,    -2,    -4,    -6,   -23,   -20,   -67,  -106,  -105,   -95,   -63,   -94,  -138,  -138,   -98,   -90,   -84,   -58,   -40,   -36,   -65,   -32,   -51,  -151,   -98,   -46,   -24,     1,    -9,     4,     5,    -7,   -41,   -45,   -75,  -102,  -142,  -156,  -187,  -200,   -31,    -8,   -16,   -26,   -46,  -106,  -147,  -121,   -81,   -59,   -54,   -92,  -123,  -124,   -71,   -16,     7,     9,     7,     4,   -54,   -77,   -31,   -60,   -41,   -10,    26,   -25,    23,    40,    36,     0,   -11,   -24,   -74,   -99,  -128,  -132,   -83,   -84,  -183,  -135,  -118,   -10,     3,     2,    -4,   -28,   -25,   -19,    25,    19,    17,     4,    18,    54,    51,     3,     9,   -45,   -19,    19,   -29,    -7,   -53,   -69,   -35,   -57,   -63,   -81,   -84,   -52,   -38,     6,    33,   -28,     8,    -9,    72,    44,    48,    37,    43,    55,    -2,    20,    33,    29,     6,    26,    35,    47,    25,   -17,   -10,   -13,   -24,   -61,  -129,   -80,   -51,   -35,    22,    -6,    36,     0,    61,     4,    17,    10,   -23,    31,    36,   -44,   -55,   -37,    22,    35,    22,    36,    29,    28,    24,   -15,    -3,   -58,   -73,   -77,   -35,    -8,    25,    29,    25,    36,     4,   -13,    -7,    -3,   -13,     7,    27,    -9,   -19,   -48,     4,     8,    48,    42,    11,    -1,    40,    13,    32,   -57,   -12,    72,   101,    -6,    46,    -7,   -24,    23,   -50,     7,   -28,     9,    13,     1,    21,   -35,   -47,    -7,     6,    37,    38,    50,    31,    28,   -11,    33,   -11,    -9,    38,    64,    86,    -4,    -1,     1,   -21,    31,    25,   -36,   -22,    -7,    30,    13,   -36,   -15,    39,   -11,    -3,    34,    18,    42,    27,   -27,     7,    44,    36,   -15,   -62,    -4,    55,    -6,    26,    38,     4,    41,    57,     5,   -37,    37,   -13,   -42,   -14,   -14,   -13,   -12,    45,    34,    40,    18,     3,    -5,    12,     3,    21,     7,    33,    57,    91,     1,    14,    55,     0,    41,    48,   -14,   -21,    15,     1,    -2,    -6,   -26,     2,   -27,    13,     6,     6,    -4,     7,   -19,   -10,    47,    16,    45,    49,    -9,   -25,    -2,    22,    19,     8,     2,    35,   -37,    23,    20,   -11,    -2,   -11,     6,   -24,   -18,     2,   -21,    26,    -2,    21,   -15,   -19,    12,   -19,   -13,   -97,   -89,   -14,     9,     0,   -10,    -4,   -20,   -31,     1,    11,     9,    22,    26,    13,   -12,     4,    23,    36,   -20,     3,    19,    21,    -7,    -3,   -29,   -59,   -83,   -99,   -11,   -66,     4,     0,   -13,   -47,    11,    26,   -27,   -32,   -18,    16,    20,     3,    19,    54,    33,    78,    18,    10,     4,   -23,   -36,   -23,    -8,   -19,   -36,   -90,   -67,   -65,    -8,   -10,   -35,   -68,    19,    10,    -6,   -37,   -32,   -68,   -19,   -26,    39,    47,    35,    32,    -6,   -22,   -30,   -27,   -18,   -14,     0,    -4,    41,   -53,   -29,   -70,    15,     6,    19,  -114,     5,   -11,   -45,   -35,   -32,   -35,   -29,    -4,     8,    13,    20,   -21,   -62,     4,    -2,   -28,    47,    43,    13,    46,    13,   -82,     9,   -47,     9,    12,    -6,   -43,   -32,    -7,   -22,   -52,    -2,   -29,   -38,    -9,    21,    32,    -9,   -67,    -5,     2,    -8,    -7,    16,    54,   -18,   -43,    32,   -87,   -76,   -26,    -4,    -5,   -23,   -25,   -90,   -68,   -53,   -36,   -68,   -25,   -64,   -61,   -27,    17,     8,   -35,    -9,     4,   -73,    -7,     7,    13,   -33,   -85,   -35,   -74,   -64,     7,    -6,     2,   -35,   -61,   -83,    -9,   -21,   -21,   -26,   -60,   -16,   -23,   -18,    15,   -22,   -13,    10,     1,   -56,   -27,   -33,    42,   -32,   -74,  -106,   -28,   -20,     1,   -14,   -15,   -46,   -58,    -3,    10,    -1,   -23,    24,    -3,   -23,    -9,    11,   -27,    -2,     5,    45,    -6,   -12,    15,    41,    -4,   -47,  -191,  -102,   -10,   -31,     0,     4,   -10,   -36,   -68,    13,    17,    15,    12,    43,    22,     1,    18,    54,    32,    64,    10,    33,    30,     2,     0,    31,    -7,   -46,  -166,   -89,   -46,   -75,    -5,    -8,     5,    29,   -22,    65,    64,    63,    59,    56,     3,    30,    43,    49,   102,    89,     6,    58,    41,     9,    35,    32,    19,   -13,  -116,   -63,   -66,   -49,     7,    -1,    -6,    -8,    26,    28,    37,    31,    37,    32,    43,    75,    71,    54,    46,    19,   -27,    88,    34,    24,    25,    -2,    47,    53,   -17,   -16,   -51,   -36,     6,    -2,     5,     8,   -34,   -27,   -49,     3,    36,    37,    55,    58,    61,    56,   -48,   -87,    -9,    36,     6,    16,    54,    30,    45,    56,    19,   -25,    -6,    -7,    -2,    -5,     6,    -6,    -2,    19,    21,   -14,   -24,    -3,    26,    45,     9,    -5,   -66,   -15,    17,   -26,    31,    19,    22,    14,    46,    23,    61,     5,     0,    -8,     3),
		    58 => (    5,    -3,    -2,     2,     5,    -8,    -6,    10,    -3,     4,    -7,   -10,    -4,    -9,     1,     4,     2,    -8,     8,    -3,     6,     0,    10,    -3,     1,     1,     0,     9,     2,     2,    -6,    -9,    -7,     6,     2,     3,    -3,     3,     9,   -14,   -28,   -17,   -20,   -11,   -30,   -30,   -33,   -14,     5,     6,    -5,    10,     2,     8,    -3,     5,    -7,    -9,    -6,    -2,    -4,    -9,   -16,   -23,   -61,   -59,   -85,   -42,    -5,    -6,   -33,   -33,   -50,    11,     6,   -28,   -27,   -27,   -27,   -11,   -10,    -8,    -2,    -5,    -2,    -2,   -16,   -22,   -14,   -33,   -64,  -119,    12,    30,    29,    -5,   -32,   -40,   -28,    34,   -37,   -49,     8,   -30,   -24,   -28,    28,    54,     1,   -20,   -31,     8,    -4,   -30,   -27,   -74,   -62,   -70,   -39,    41,    90,    76,    60,    31,   -10,    -5,    26,    30,    25,    63,   -12,   -39,   -53,   -64,   -30,   -54,   -70,     7,    36,   -14,     3,     8,   -52,   -61,   -51,   -74,    -7,   101,    37,    43,    25,    52,    56,    25,     6,    15,    27,    57,    -3,    60,    -4,     9,    23,   -18,   -25,   -17,   -53,   -21,     4,    -9,   -80,   -67,   -70,   -36,   -25,    47,   -20,     4,    39,     7,    -5,    15,    -7,    18,    -4,   -14,    16,    17,    39,     2,    -7,    28,   -20,   -33,   -17,   -12,     4,   -54,   -66,   -78,   -65,   -49,    -1,     6,    -9,    -3,    -9,    41,    -1,    13,   -39,    28,    14,    -8,   -13,    11,   -24,   -11,   -19,    74,    45,   -75,   -50,    24,    18,   -37,   -58,     7,    -7,    -5,    -9,    40,    17,     8,    11,     2,    -8,     9,    -4,    -8,   -12,    -4,    27,    67,   -27,    55,    43,    70,    76,   -44,    65,    71,     5,   -19,   -75,    17,    40,   -22,     2,    35,    18,     0,   -26,     1,    -6,     1,    22,   -12,   -14,    20,     9,    -8,    46,    42,    45,    32,    14,   -21,    64,   -82,    -6,    -6,   -89,   -61,    82,    24,   -29,    28,    29,    14,    39,    14,    15,   -10,    39,   -66,   -51,     5,   -10,     1,    13,    48,    22,    45,    34,   -67,    26,   -32,     6,   -10,   -41,    -1,    76,    65,    16,    45,    13,     5,    17,     0,   -20,   -20,    14,   -58,   -52,   -39,     4,    -2,    21,    30,    34,    41,    50,    17,    76,   -16,    -5,     5,   -61,    16,    74,   130,     4,     6,    46,    20,    -2,   -27,   -41,   -40,    -6,   -30,     2,    -4,   -31,   -20,    27,    29,    68,     8,    30,   -29,    39,   -70,     9,    -6,   -38,    -4,    26,    73,    24,    13,    32,     5,    -5,   -10,   -10,   -16,    -9,    11,     1,   -53,   -26,   -20,    34,    14,    59,     3,   -39,   -42,    30,    11,     2,   -16,   -16,   -47,   -70,     9,    45,   -62,    35,   -81,   -56,   -16,   -32,   -36,     3,     7,   -21,   -56,     2,   -47,   -67,    20,    -3,   -20,   -55,    -8,   -34,   -23,     6,     6,   -28,    24,  -118,   -28,   -38,   -45,    19,   -48,   -16,   -16,   -57,     6,    21,   -31,   -24,     6,   -43,   -19,   -33,   -52,   -17,   -65,   -84,   -19,   -91,   -54,     6,   -11,   -17,    33,  -111,   -47,   -57,   -92,   -50,    -5,   -59,   -40,    -7,    31,    -3,   -17,   -43,   -77,   -38,    -5,   -42,   -60,   -32,   -20,   -31,   -31,  -103,   -53,     3,   -11,   -24,   -54,   -31,   -56,   -63,   -60,    -8,   -40,   -39,   -64,   -16,   -20,   -31,   -59,   -28,   -25,   -27,   -14,     6,   -15,   -16,    -9,   -11,   -98,   -47,   -76,   -12,   -14,   -37,  -101,     1,   -56,     1,    17,     8,    -8,   -19,   -26,    11,    -4,   -36,  -107,    -4,    10,     2,    19,    -9,   -18,     4,    -1,     3,   -91,   -40,   -50,     6,     4,   -75,   -94,   -21,   -56,   -35,    17,    60,    16,    11,   -22,   -39,   -36,   -64,   -44,   -12,    45,     5,    20,    22,   -32,    14,    47,    61,  -120,   -90,   -59,     4,     2,   -28,   -77,   -60,    13,    30,     8,    53,   -21,    54,    -3,    27,     2,   -40,   -14,    47,    32,     8,     1,    39,    41,    38,    98,    23,  -146,   -92,     4,   -25,   -39,   -35,   -42,   -49,    10,    66,     8,    41,    67,    30,    26,    15,    36,    31,    79,    -3,    54,   -57,    25,     5,     6,    74,    64,   -26,  -111,   -69,    -1,   -26,   -33,   -18,   -35,    29,    67,    40,    61,    53,    53,    74,    73,    33,    54,    91,    94,    15,    12,    22,   -21,     0,     2,    63,    36,   -35,    -6,   -69,    -5,    -8,     6,   -11,   -18,    64,    -6,    24,   -14,    28,    30,     8,    10,    61,    61,    60,    67,    59,    50,    60,    84,    20,   -23,    86,    44,   -21,    -8,   -71,     0,     8,     2,   -28,   -43,   -25,   -27,   -15,   -22,    23,    43,    19,     8,    56,    18,    25,    41,    86,    -9,    -5,   -11,     9,   -43,    11,    15,   -40,   -96,   -50,    -8,     9,    -2,   -30,     3,  -119,   -95,    -6,    -8,   -40,   -70,   -37,   -39,   -24,   -20,    27,    33,   -11,   -23,    18,    -9,   -68,   -61,   -64,   -33,   -38,   -24,   -14,     1,     3,     4,     1,   -27,   -54,   -94,   -88,   -21,    16,     6,   -46,   -25,    22,    14,   -76,  -162,   -74,   -44,   -37,  -120,  -103,   -49,   -56,   -21,    -5,     4,     0,    -7,     0,     1,    -4,     5,   -24,   -20,   -25,   -16,   -33,   -29,    -7,    -9,   -40,   -65,   -77,   -62,   -33,   -51,   -26,   -28,     0,     0,   -21,     0,    -3,    -8,     3,    -3),
		    59 => (    7,    -5,     9,    -3,    -8,     7,    -5,    -7,     9,    -1,     8,    -6,     4,     5,    -4,    -9,    -6,   -10,    -6,    -4,     9,    -4,   -10,     9,     9,     7,     5,    -6,     3,     7,     1,    -8,    -8,     7,     2,     0,   -10,    -3,     1,   -12,   -17,   -22,     8,   -13,    -5,   -17,    -2,     7,     5,     8,     4,    -7,    -6,    -8,    -9,     7,    -4,    -7,     3,     7,   -10,     6,    -8,    -7,   -16,   -10,    -4,   -17,    -7,    -9,   -30,    -9,     7,    -9,     5,    -7,    -8,     5,    -4,     2,    -6,    -7,    -2,     6,    -2,    -5,     6,    -8,   -14,   -20,   -16,    -2,   -25,   -40,   -12,   -31,   -10,   -42,   -29,   -32,    -8,     6,    17,     2,   -40,   -30,   -12,   -11,     2,   -12,     2,    10,     8,    -2,     6,    -2,    -3,   -10,   -40,   -14,   -12,    -2,   -20,     2,   -57,   -76,   -63,   -52,   -44,   -43,   -21,   -55,   -61,     0,    -8,     1,    -7,   -43,   -35,    -9,    -9,    -1,     0,    -3,   -10,     4,    -9,   -25,   -79,   -31,   -38,     4,    12,    -1,    13,    -2,   -19,   -61,   -77,   -43,    -9,   -13,     1,    -4,     4,   -39,   -20,     5,    -4,     5,   -12,    -7,   -28,   -43,   -38,   -59,   -13,    27,     5,    46,    46,    37,    -4,   -21,    29,   -13,   -99,   -93,   -44,     1,     4,    -7,     0,     1,    -6,   -27,   -10,    -1,   -11,     7,   -20,   -47,   -74,   -56,    -4,   -35,    12,    41,     5,    20,   -23,   -61,   -48,   -51,  -107,  -138,   -48,     9,    -2,     1,   -18,    -1,    -9,   -22,   -19,   -11,   -20,    25,     7,   -51,    43,   -11,    36,     3,    -3,     8,   -13,     7,   -11,   -46,   -51,   -28,    14,   -34,   -74,   -13,   -13,   -18,   -23,    -7,    -4,    -1,    -6,   -36,   -33,    14,    -3,   -32,    33,    30,    13,    25,    41,   -22,   -25,    11,     7,   -40,   -62,    28,    26,   -25,   -47,   -39,   -47,   -19,   -36,   -47,   -22,   -22,    -3,   -11,   -16,    15,   -10,   -51,    43,    23,    18,     7,     4,   -85,   -74,    13,    49,    -9,    28,    -2,    -2,   -25,   -44,   -48,   -55,   -35,   -31,   -39,    -7,   -37,    -6,   -54,   -23,    26,   -23,   -57,    19,    46,    34,     9,   -17,    -8,    30,   103,    -3,    -9,    -9,    36,   -15,    -6,   -73,   -81,   -52,   -49,   -17,   -34,     2,   -33,     8,   -21,   -22,    34,   -18,    18,    17,    -8,    -3,    40,    19,     7,    33,    69,   -27,   -55,   -12,    29,     0,    -3,   -28,   -45,   -71,   -54,   -32,   -27,   -30,   -37,     6,   -22,   -17,   -27,   -35,     3,    87,    12,   -41,     7,    14,   -18,     0,   -13,   -19,   -12,    -4,    -7,   -31,    19,   -32,   -42,   -40,   -39,   -18,   -21,   -26,    -1,    -9,    -5,   -16,   -19,   -25,   -23,    56,     6,   -22,   -17,    44,    -2,   -31,   -20,    14,    16,   -12,     1,     2,    -1,   -30,   -54,   -58,   -58,   -26,   -41,    -3,    -3,   -10,    -2,   -16,   -21,    28,   -38,   -37,     7,   -11,   -28,    21,     8,   -21,   -58,   -26,    15,    17,    -2,   -15,   -14,   -90,   -80,   -55,   -51,   -15,   -10,     0,   -25,    -7,    -1,   -28,    -5,    -2,   -23,   -86,    -8,    16,   -33,    11,    95,    33,    13,     6,   -41,   -33,   -34,   -12,   -35,  -117,   -44,   -25,   -19,   -16,   -11,     3,   -41,    -4,    -5,   -36,     4,    -2,   -31,   -68,   -81,    -8,   -60,   -21,    26,    45,    29,     6,     5,   -46,   -50,   -32,   -26,   -77,   -49,   -18,   -29,   -44,    34,   -30,   -20,   -10,     0,   -33,    -3,     3,    -1,   -21,   -50,   -65,   -61,   -65,   -26,    34,   -17,   -15,   -21,   -13,    -2,   -45,   -16,   -32,   -55,     1,   -19,   -51,    -7,   -26,   -20,   -10,    -3,   -26,    -6,     0,   -16,    -9,    -2,   -13,   -11,   -53,   -83,   -77,   -74,   -55,    30,    16,     5,   -30,   -31,   -49,   -56,   -28,     0,   -35,    37,   -25,   -22,    -5,   -13,    -1,   -16,    -3,    -2,    -3,   -39,    -2,   -39,   -43,   -72,   -95,   -57,    -3,     8,    -8,   -13,   -25,   -29,   -22,   -18,   -21,   -25,     8,    24,   -33,     2,     7,   -10,     4,   -15,    -8,    29,   -12,   -14,    -5,     6,     9,   -11,   -25,    -9,     9,   -31,    -6,     1,    -1,   -53,   -20,   -34,   -18,    -9,    19,    39,   -44,   -10,    -2,    -6,   -13,    26,     0,     9,    17,    16,    19,    30,   -14,    11,    29,    13,    11,    20,    -6,    21,   -12,   -48,   -32,   -55,   -11,     0,    14,   -10,    -3,    -6,     8,     6,   -21,    13,    -9,    -8,    21,    -4,    16,   -13,     9,   -12,     1,    -3,    -6,    29,     2,    19,    28,   -20,   -22,   -26,    -6,    19,    11,    10,   -22,     1,    -2,    -2,    -3,    -4,   -10,     7,     0,   -27,     3,   -20,    24,   -25,   -68,   -52,   -16,    13,    25,    17,    19,    24,    19,     4,    -6,    15,    10,    15,    -6,     2,    -2,    -3,    17,    -5,    -6,     3,     5,   -16,   -12,    15,   -32,   -41,   -26,    10,   -50,   -40,     8,    38,    11,   -41,   -50,   -43,   -38,   -18,   -14,    14,     3,     7,     4,    -5,     7,    17,     2,    -1,     2,     5,    10,    26,   -20,   -44,    40,     3,    41,    23,    13,    91,    34,   -42,     8,     4,    -8,    13,    13,     7,     0,   -10,    -9,    -6,     0,    -7,    -7,    -9,    18,    23,    11,   -29,   -14,     9,    -3,   -30,   -38,    73,    68,    -7,   -15,    33,    14,   -27,   -22,    -6,    -3,    -2,     8,     3),
		    60 => (    3,     1,     6,     7,     8,    -1,     8,     7,    -2,     2,     4,    10,     1,    -1,    -9,     5,    -3,    -8,    -8,    -9,     6,     6,     0,    -9,     0,     1,    -3,    10,    -1,    -4,     9,     2,     0,     5,    -4,   -21,   -18,   -24,   -44,   -19,     7,    12,   -57,    55,    68,    70,     3,   -10,   -14,   -12,     6,    -1,     6,     5,    -1,    -1,    -2,    -7,     8,    59,    71,   -20,   -33,    10,   -14,   -39,   -64,   -54,   -69,  -132,   -68,   -32,    -4,   -50,   -33,   -35,   -38,   -32,   -92,   -35,   -44,    -8,     4,     9,     6,    -5,     7,    62,    21,   -60,   -70,   -60,   -58,   -47,   -32,   -74,  -103,   -49,   -57,   -62,    24,    25,     1,   -48,   -48,   -71,  -101,   -50,   -37,   -42,   -74,     8,    -1,    -1,    -6,   -18,   -24,  -122,   -45,   -52,     5,    53,    -6,    10,   -59,     0,   -23,    21,    54,    26,    -4,     2,   -44,   -44,   -18,   -26,   -83,  -140,   -57,     4,    -3,   -10,   -31,   -20,   -28,   -62,    27,   -11,    13,    77,    49,    41,     9,     6,    33,    30,    31,    33,    31,     1,    -3,    -8,   -35,   -25,   -77,  -121,   -28,   -15,     5,     3,   -43,    -4,   -80,    22,    49,    47,    43,    30,    52,    25,     6,     3,    27,   -28,    11,   -10,   -39,    14,    -8,   -47,    -2,   -93,   -52,  -140,   -40,   -13,    -1,   -20,   -38,   -43,   -47,    -3,    43,    43,   -21,    22,   -14,     8,    13,    16,   -44,   -50,   -22,   -11,   -17,   -44,   -14,   -40,    -9,    -3,   -49,   -26,   -73,    12,    91,   -57,    -4,   -61,   -57,     4,     6,   -45,     9,    16,   -23,   -44,     3,   -13,   -74,    -6,   -16,    36,    -6,   -21,   -25,    10,     0,    34,   -58,  -134,   -69,   -16,   -11,   -16,    33,    -2,   -14,    15,   -46,   -24,   -10,    21,   -18,    17,    37,    14,    16,    35,    25,    32,    16,    21,    16,   -14,    -1,    34,   -14,   -81,   -22,   -15,   -14,   -12,    42,    17,     7,   -29,   -12,   -28,     7,    28,    -9,   -13,    -2,    30,    91,    67,    62,    75,   -12,    27,    18,   -26,    14,    35,    -2,   -48,   -60,     0,    -7,    98,   -59,    -8,   -17,   -57,   -21,   -30,   -39,   -17,   -27,    -6,    24,   109,    41,    50,   120,    93,    80,    49,    38,    19,    19,    23,    59,   -57,   -61,    -5,    -7,     3,   -61,   -21,    31,   -59,   -53,   -62,   -49,   -11,   -22,     5,    58,    83,    57,    68,    48,    44,    46,    31,   -23,     3,    -4,    15,    30,   -29,   -48,   -32,     2,     9,     0,   -26,    42,    -9,     5,   -34,   -11,   -39,   -30,    17,    23,     7,    -3,    11,     2,   -19,   -10,   -16,   -21,    15,    10,    48,    17,    26,   -85,   -30,    -8,     0,   -11,   -78,   -29,   -14,   -36,   -11,    -3,   -24,   -25,     2,   -23,   -15,   -76,   -88,   -88,   -38,    22,   -15,    34,    71,    73,    40,    68,    57,   -72,    -9,    -7,     6,   -50,   -71,   -15,   -35,   -45,    19,    -3,   -53,   -47,   -36,   -56,   -54,  -119,   -68,   -47,   -14,   -27,    -4,    42,    30,     8,    31,    51,    62,   -77,   -68,    -9,     1,   -29,   -35,    27,   -18,   -51,    12,   -10,   -27,     2,   -26,   -45,   -65,   -68,    -9,   -55,   -49,   -17,    29,    26,   -16,   -26,   -45,    -8,   -22,  -109,   -24,     3,    -6,   -38,     3,    12,     8,   -31,    20,    -9,    12,    23,    37,    15,    40,   -26,   -26,   -42,    -9,    -9,    26,    -7,   -65,   -15,   -23,   -12,   -70,   -69,    19,    -5,    -2,   -33,   -23,    37,    33,    25,   -15,    10,    40,    45,    19,     6,   -25,   -52,   -18,   -18,    14,    11,    10,   -48,   -37,   -23,    24,   -60,   -66,   -54,   -38,     7,    15,   -11,   -21,     1,    53,    35,    60,    45,    12,     1,    10,    47,   -20,   -30,    -1,    -3,     6,     6,    49,   -24,   -35,   -11,    24,    -3,  -109,   -15,   -11,     2,    16,   -47,   -36,    58,    37,    28,    47,    25,    71,     0,    22,    68,    19,     5,    25,     1,    18,    -4,     9,   -44,   -54,   -26,   -15,   -37,  -127,    10,     3,     6,    -9,   -48,   -28,     5,    -7,    51,    70,    57,    42,    28,     8,    40,     4,   -12,    26,    16,     1,    17,    13,   -19,   -39,    -6,     8,   -64,   -61,   124,    -1,    -6,    -4,   -26,   -28,   -84,   -47,   -10,    67,    53,     8,    72,    34,    -8,   -23,    18,    45,    28,    21,   -18,   -16,   -49,   -50,   -20,    -4,   -44,   -26,    75,    15,     3,     8,   -24,   -57,   -19,   -53,   -44,    -6,    48,    39,    28,   -35,    37,   -11,     9,    22,    19,    50,   -11,   -54,   -85,   -58,   -72,   -23,   -49,   -66,   -64,   -10,    10,    -7,   -18,   -29,    17,    32,   -55,   -33,   -30,   -15,   -28,   -91,   -58,   -54,   -51,    29,   -10,    -3,   -33,   -78,   -44,   -80,   -68,   -50,   -43,   -22,    -5,     1,     5,     6,    -8,   -19,   -78,   -49,   -86,  -129,   -72,   -76,   -83,   -48,   -75,   -45,   -52,   -66,  -144,  -124,  -125,  -141,   -98,  -112,   -79,   -36,    -7,    -3,     9,     9,    -2,     0,    -5,     2,   -26,   -79,  -110,   -53,   -42,   -76,   -54,   -61,   -40,   -47,   -61,   -97,   -81,   -73,   -73,   -89,   -78,   -91,   -57,   -37,   -22,    -4,    -5,     1,    -1,     1,     0,     2,     0,     1,    -5,   -14,   -24,   -44,     3,    -3,     1,   -58,   -20,   -10,    -1,     7,   -33,   -30,   -23,   -44,   -22,   -34,     3,     6,    -8,    10),
		    61 => (   -5,    -6,     6,    -2,    -9,     6,    -8,     6,     0,    -3,    -9,     2,     2,     5,    -8,    -1,    -9,    -9,    -4,     6,    -6,    -1,    -2,    -7,     1,    10,    -5,    -4,     9,     0,     1,     1,     1,     4,    -1,     1,     2,     5,    -3,    -5,   -16,   -17,    13,     4,   -15,   -11,     1,     9,     8,    -7,    -1,     4,     8,     3,     5,     8,     1,     7,     5,     3,    -6,    -6,    -5,     7,    -6,    -8,    -2,    -1,   -37,   -39,   -37,   -79,   -79,   -33,   -23,    -4,    22,   -25,   -18,    -7,   -22,   -20,     5,    -4,     3,     2,    81,    54,     9,   -14,     3,    31,    13,     8,   -12,    -7,   -63,  -157,  -121,   -94,   -63,   -57,   -37,     1,    -5,   -10,    91,    16,    -5,   -25,    -3,    10,    10,    -8,    68,    56,    24,   -21,   -37,   -23,   -60,   -28,   -51,   -59,   -99,  -109,    49,    25,    38,    27,    23,    20,     5,    23,    25,   -30,   -51,   -61,   -53,   -44,     8,    -9,    52,    79,    47,    13,   -17,   -28,  -119,   -72,  -111,  -106,  -104,   -61,     3,    24,   -15,   -28,   -68,   -35,   -15,    19,    44,    -2,   -40,   -66,   -59,   -56,    -5,    -2,   -41,    34,    68,   -34,    48,    73,   -46,  -110,  -124,  -118,   -60,   -23,    -5,   -23,   -14,     6,   -27,   -16,    24,     1,     4,   -13,   -52,   -52,   -33,   -29,    -9,   -57,   -71,   -12,   -46,    52,    55,    68,   -82,   -81,  -180,  -103,   -55,   -24,    -3,     3,    28,    23,    -1,    36,    43,     8,   -36,   -23,   -61,   -43,   -36,   -25,    -1,   -55,   -59,    21,   -45,    37,    48,    16,   -51,   -60,   -76,   -88,  -100,   -49,    -5,    29,    25,    24,    11,    23,    19,     7,   -25,   -46,   -83,   -33,   -70,   -10,     6,    -5,   -53,    11,   -26,   -35,    43,    63,    36,    14,   -16,  -100,   -29,   -76,    -6,    47,    76,    20,    28,     5,    -8,   -30,   -29,   -23,   -52,   -17,    -5,   -19,    -8,    24,   -59,   -20,   -27,   -53,    -3,    48,   -18,   -11,    31,   -10,   -33,   -64,    -4,    16,    29,    21,   -14,   -28,   -72,   -96,     3,    -9,   -45,    -2,     0,    60,     4,     5,   -11,    28,    -3,    47,    32,   -67,   -90,   -33,    21,   -23,   -92,     2,    10,    22,    19,     1,   -32,   -83,   -30,   -18,     1,   -19,   -11,     0,     3,    48,    -1,     5,   -25,    46,   -13,    60,    55,   -21,   -35,     6,    -9,   -34,   -27,    21,    39,    10,    20,    27,   -49,   -66,   -20,    48,   -14,   -27,   -41,    33,    -4,    42,    -6,    -2,   -15,    31,    17,    24,    48,    14,    30,    34,   -18,   -43,   -38,     0,    42,    -4,    10,    43,   -81,  -134,   -71,    41,   -31,   -34,   -47,     2,     8,     8,    -5,    -2,    31,    19,    66,   -32,   -36,   -99,    30,    -3,     8,   -26,   -28,    16,    17,   -23,    25,   -18,     6,   -61,   -43,    67,    40,    -7,   -23,    55,    64,    -1,     4,     0,     6,    69,    31,   -78,    -3,   -12,    34,     4,   -16,    18,    -4,    15,   -28,   -27,    46,    31,   -90,   -97,   -31,     8,    -4,   -36,   -47,    29,    30,   -15,     1,    10,    30,   -14,    -4,     6,     0,   -56,     5,    -2,   -70,    12,   -24,    25,   -10,    -9,    45,     8,   -52,   -98,   -55,    25,     1,    27,    33,    14,    -1,   -13,   -10,     6,     3,   -58,    17,    -6,    11,   -17,   -25,   -32,   -47,    34,     7,    22,    -8,   -39,   -10,   -79,   -68,   -52,   -38,    12,   -23,     3,    18,    29,    -9,    -9,   -10,    -5,    -9,   -13,   -23,   -76,   -57,   -59,   -12,     1,   -11,    15,     8,    18,   -12,   -30,   -70,   -68,   -44,   -64,   -57,     8,     1,    30,    11,    34,     4,    40,    -9,    -6,    33,    17,    -1,   -63,   -20,   -38,    -8,    28,     5,    20,   -10,    25,    -2,     5,   -50,   -35,   -19,   -62,   -45,    -6,   -36,    34,    47,    55,    12,    36,    -1,     1,    32,    -5,    30,   -15,   -10,   -32,     1,   -30,     7,     3,   -20,    15,    32,   -15,    -5,   -60,    -4,   -21,    35,   -21,   -10,    22,    70,    60,     7,    -5,    37,    47,    39,    29,    15,    42,   -26,    -6,     3,   -21,    16,   -35,    -2,     2,     7,     7,   -37,   -79,    -2,    28,    65,    22,    -5,    36,    60,    32,     3,    -4,    30,    45,    30,    28,    -9,    18,     8,   -50,   -43,   -14,   -34,   -34,    -4,    -2,    39,    64,    28,     7,    70,    33,     2,   -10,    13,    45,     8,    -8,    21,     2,     9,     8,    -2,    -8,   -14,    -9,    38,    54,    68,    74,    -8,   -16,    -9,    15,    18,    78,    32,    49,    37,    -5,   -60,   -61,   -15,   -18,    24,    53,    79,    -8,     4,     2,     4,   -20,   -74,   -70,   -64,    -8,    -6,    70,   -26,   -19,   -22,     6,     5,    48,   -10,    -6,   -12,    14,    -4,    28,     5,   -30,   -23,    33,    23,     0,     7,     4,     8,   -16,   -38,   -30,   -24,  -104,    -3,    47,  -130,  -107,     0,   -13,    36,   -16,   -56,  -107,   -58,   -33,   -54,   -38,   -28,   -21,    -7,     5,     0,    -7,    -8,    -1,    -4,     5,   -15,   -35,   -79,   -98,   -87,   -88,   -34,   -48,   -85,   -87,   -46,   -24,    25,   -52,    -5,   -15,    -9,   -15,    -2,    -2,     9,   -10,    -8,    -5,    -2,     7,     8,    -1,     6,     6,    -1,    -7,    -4,   -13,   -43,   -36,    -2,    -7,   -32,   -11,   -20,     6,    10,    -7,     2,    -2,    -3,     2,     1,     3,     3,     8),
		    62 => (   -6,     3,     1,     4,     9,    -4,     3,     2,    -3,     0,   -10,    -3,    -6,     6,    16,     9,     8,    -6,     7,     9,    -1,     6,    -3,     1,    -7,    -2,    -9,    -1,     8,     4,    -3,    -9,    -1,    -2,    -9,     5,     5,    16,     8,    -4,    -1,     1,    -4,   -27,    26,    11,     2,   -41,   -11,   -10,    -1,     1,     1,     7,     0,     7,     5,     5,    -7,     1,   -14,    -8,    10,    -5,    10,    -9,    20,    73,    56,    88,    35,   -13,   -24,   -28,   -50,  -124,   -92,   -22,   -20,    -7,     1,    14,    -2,    -1,    -1,    -5,    -9,   -34,   -33,    21,    51,    -6,   -12,    39,   -19,     9,   -15,     5,     0,    14,    41,     2,   -65,   -55,   -62,   -37,    35,     5,    -2,    -5,     8,    -2,     8,     7,   -23,    20,    24,    33,    86,    83,   -22,     6,    46,    49,    34,    75,    51,    46,     1,     9,     8,   -36,    12,    19,    12,   -55,   -59,   -21,   -35,   -10,     5,     8,    13,     3,    -9,   -36,   -28,    51,    -9,   -28,    17,     7,    27,    22,     2,    26,    28,    -3,     5,    -8,   -43,    29,    65,     9,   -31,   -33,   -39,   -20,     4,     3,    24,    17,   -15,   -58,    17,    21,   -12,     2,   -10,   -21,     0,   -12,    27,    -4,    -1,   -32,    14,   -43,     6,    27,    83,    18,   -30,   -43,   -22,   -12,    -6,     1,    -8,    42,    -2,   -19,   -57,    -3,    26,   -10,    23,    -2,     8,    18,    49,    36,    -4,   -23,   -25,   -53,    15,     0,    37,   -60,   -48,   -66,   -14,   -17,   -29,    22,    20,     5,    43,   -28,   -44,   -21,    13,     0,    40,    38,    -8,   -24,   -34,     8,     8,     5,   -10,    -3,     1,    -3,     9,     1,   -31,   -39,   -46,   -12,    -3,   -23,    77,   -20,    34,    43,   -53,     6,    -5,     3,    -3,   -35,     8,   -90,  -146,   -15,    21,    16,    -3,   -10,    -1,    -2,    -3,    28,   -68,   -36,    20,   -22,    -7,   -13,    43,    17,   -13,    -4,   -21,    50,    17,   -36,   -31,   -38,   -78,  -114,   -54,   -45,     6,     0,   -26,    -5,   -39,    14,   -67,    31,   -28,   -17,    27,   -11,     2,     1,   -18,    33,    38,   -13,    -1,   -11,   -14,   -85,   -65,  -108,  -124,  -127,   -28,   -14,     2,   -38,   -48,   -38,   -14,   -22,   -32,    50,     2,     2,   -25,    -3,     7,    -5,   -26,   -15,    -3,   -10,   -36,  -106,   -83,   -97,   -95,   -75,   -93,   -34,    -5,   -36,    27,    -7,   -43,   -39,    -6,     2,   -31,    33,    -5,    17,    45,   -21,     2,     7,    32,     1,   -23,   -57,   -95,  -139,  -157,  -151,   -78,   -65,   -29,    44,   -24,   -28,    19,    -3,   -21,   -57,   -46,   -16,   -41,     8,   -19,    -4,    46,     7,     0,   -14,   -18,    -5,    -6,   -65,   -79,  -109,  -117,   -78,   -15,   -10,     4,    13,   -37,   -35,    -4,   -12,   -51,   -35,   -46,    -9,     2,   -14,   -16,     4,    30,    31,    -8,   -23,    -2,    -8,   -68,   -51,   -20,   -42,   -13,    33,    45,    28,   -22,    17,   -14,   -30,    -7,   -36,   -54,   -37,   -69,     8,    -5,   -21,    -9,    28,    31,    66,    -8,    -1,    -4,   -28,   -57,   -38,     1,   -41,   -25,    17,    12,    20,     5,     5,    11,   -68,   -13,   -42,   -80,   -43,   -69,   -19,     1,    -4,   -21,    74,    33,    27,     5,     2,     6,    -8,   -47,   -14,   -55,   -26,    -9,     4,     8,    23,    37,    21,    -9,   -23,   -37,   -63,   -93,   -56,     8,    -2,   -51,   -51,   -39,    37,   -13,    28,     9,     6,   -20,    18,    45,   -12,   -10,   -14,    47,    30,    12,    13,    57,   -13,   -12,   -80,   -59,   -45,   -13,   -21,     6,     9,    -3,   -35,   -26,    98,   -35,    65,     6,    -7,    15,    44,    40,     6,    -4,    33,    64,   -14,    30,    28,    58,    33,   -40,   -28,   -44,   -65,   -18,    -5,     2,     1,   -46,   -59,    35,    37,    56,    72,    -1,    -4,    45,    54,    55,    49,   -47,    22,    -6,    -6,    15,    28,    42,    23,    -2,    32,     5,    41,   -54,     8,    14,    20,    -1,    -9,    32,    39,    50,    10,    -5,    23,    56,    48,    35,    28,   -30,   -21,   -22,    14,    15,    -1,    27,    -9,    -3,    14,    32,   -26,     5,    48,    11,    30,    35,    33,    93,   106,    35,    -5,     2,    -5,    50,    48,    14,     0,    -9,     6,    17,   -23,    24,     9,    14,    -4,    30,    34,     7,   -76,   -17,    27,    34,   -12,    21,   -29,    -3,    14,   -42,   -22,    -7,    -4,    -8,    11,   -29,    21,    -2,    15,    49,    -4,    -9,    25,    -1,   -23,    19,    53,    13,   -49,    36,    17,    -1,    39,    27,    41,    33,    23,   -30,    -3,    -5,     0,   -33,   -17,   -37,   -58,   -98,  -142,   -90,   -39,     4,    12,    17,    19,    72,     6,   -34,    14,    46,    44,   -40,    27,   109,    64,    64,    23,    26,    -8,     2,    -6,   -15,   -11,   -15,   -31,   -23,   -48,   -90,   -93,   -18,    -5,   -17,    -1,    50,    59,    30,    84,    -9,   -82,     7,    18,    14,     2,    33,    31,    24,     7,    -5,     2,   -10,     1,    -4,    -9,   -25,   -22,   -25,   -13,    -7,   -40,    -2,   -54,   -54,   -35,   -88,   -61,   -43,   -19,    -7,    -5,   -29,     4,   -10,    -8,     2,     7,    10,     9,     5,     8,     8,     8,   -10,     6,     7,     5,    -7,    -7,    -4,    -8,     1,     7,    -8,    -9,     6,    -9,   -24,   -19,    -3,    -8,     2,    -6,     1,     9),
		    63 => (    6,     8,     8,     1,     1,     6,    -7,    -1,    -4,    -8,    -2,    -6,    -6,    -3,    -2,   -11,    10,    -3,    -9,    -3,     3,    -4,     1,    -8,     3,    -7,    10,    -6,    10,     2,    -2,    -5,     5,   -10,     3,    -6,    -3,     6,    -9,   -20,   -15,   -24,   -28,   -25,   -14,   -45,   -23,    -2,     5,    -6,     9,     3,     0,    -2,     3,    -3,     5,     1,     7,    -6,     1,    -1,    -1,   -20,   -73,   -66,    35,    33,   -26,   -52,   -71,    -1,   -25,   -18,   -10,   -13,   -52,   -40,   -33,   -38,   -17,     0,     1,    10,     9,     8,    -2,   -17,    -3,    21,    21,    55,    41,    -3,   -23,    40,    35,    30,    67,    23,   -35,   -16,   -30,   -24,    13,     1,   -86,  -129,   -65,   -47,     7,     5,    -7,    -8,   -31,    36,   -66,     7,    65,    24,    11,   -24,   -21,   -19,     9,    31,    51,    -1,    -2,   -62,   -42,   -15,   -26,    18,     9,  -158,  -143,   -74,   -64,     9,    -6,     4,    -9,    -3,   -24,   -16,    32,     4,   -30,   -52,   -10,    40,    47,     7,    18,    -9,    17,    12,    -7,    18,    19,    74,    35,    50,    39,  -135,   -25,     6,     7,    -5,    25,     9,    30,   -13,    17,    45,   -59,    -5,    19,    54,    21,    19,   -30,   -30,   -21,    13,    21,     0,    59,    68,     1,   -10,    35,   -95,   -69,   -19,     7,    14,     4,    29,    90,    27,    62,    22,     6,    -4,    16,    45,    27,     5,    34,    30,   -51,   -16,     5,    45,     0,    12,   -54,   -10,    16,   -88,  -112,   -33,   -22,    -1,     2,    12,    31,    11,   -17,   -30,     9,     6,     6,    19,    -4,   -29,    39,    23,    16,   -31,    26,    63,    30,    46,   -34,   -21,   -19,  -115,  -111,   -18,     5,   -39,    -9,   -21,    24,    23,    -4,   -18,     3,   -18,   -28,    -3,    -5,    16,    35,    18,    44,    34,    21,    19,   -19,   -26,   -21,   -29,  -132,  -140,  -130,   -46,    -2,   -50,   -34,   -33,   -10,   -39,   -44,    -6,   -18,     6,   -18,     4,    33,    27,   -27,    -1,    17,    63,    17,   -57,    -9,   -91,   -49,   -11,   -89,   -65,  -100,   -42,    -7,   -46,   -52,     8,   -19,   -18,   -15,    19,    -3,   -31,    -2,    16,     4,   -24,   -28,   -25,    -2,    94,    40,     0,   -13,   -48,   -48,   -44,  -120,  -153,   -88,    -9,    -1,   -30,   -64,     0,   -22,     6,   -11,   -31,   -21,    -6,    -2,    19,    44,    -2,   -22,   -11,    24,    53,    44,    50,    32,   -14,   -11,   -19,  -159,   -81,   -41,     0,    -6,   -19,   -47,     1,   -51,   -36,   -27,    -1,    -2,   -44,   -19,    -5,    40,    -8,   -14,   -31,    60,    51,    11,    40,    25,     9,   -35,   -19,   -12,   -99,   -76,   -26,   -15,    21,    -3,   -22,   -48,    -7,     2,    -6,   -15,   -29,     6,    20,    10,   -11,   -31,   -17,    15,    57,    42,    73,    29,    48,    -9,    -8,    27,  -105,   -71,   -12,    -1,    17,    -2,     0,   -19,    64,    59,     2,    -2,   -18,   -36,    -6,   -30,    -6,   -39,   -24,    19,    29,    22,    47,    26,    12,    21,    14,    49,   -71,   -40,   -21,    -1,    10,     3,    22,    -4,    20,    67,    34,   -16,    -1,    -5,     5,    12,   -25,   -34,   -37,    38,    58,    35,    15,    49,    41,    -9,   -28,    -1,   -99,  -107,   -37,    -3,    -3,    -5,    50,   -11,   -11,    57,    63,   -31,   -23,    -7,     4,    23,   -14,   -56,     6,    40,    39,   -11,   -26,    -7,    -7,   -16,   -21,  -108,   -99,   -48,   -11,   -26,     9,    15,    53,     4,   -10,    48,    22,     6,    16,    33,    16,    -2,   -62,   -18,    31,    33,    -1,   -25,     1,    14,    10,   -24,   -40,   -96,  -101,   -23,   -26,     3,   -41,    -9,     2,    47,    47,    31,    54,    24,    22,    32,    -5,   -71,   -78,   -37,    -3,   -61,   -65,   -20,   -11,    -7,   -26,    38,     8,   -61,   -92,   -91,   -45,    -3,   -22,   -26,   -15,    16,    59,    36,    45,   -10,    15,    20,    27,   -71,   -61,   -38,   -39,   -69,   -75,   -41,   -23,   -28,   -59,    52,    -7,   -16,   -68,   -20,    -9,    -4,    -7,    23,     6,   -14,    19,    38,     7,    -9,    -1,    26,    66,    11,   -52,    -7,     5,    -2,   -28,    -6,    12,   -13,     1,    18,    -3,   -48,   -74,   -33,     8,   -19,   -17,    31,     1,   -12,    18,    29,   -20,    14,   -13,    65,    73,    46,   -40,   -16,    40,     7,    10,    25,   -14,    -1,    -4,    46,   -21,   -96,   -62,   -51,    -8,    -1,     9,    11,    10,     0,    -1,   -12,     9,     9,    39,    64,    77,    16,    50,    37,    52,    28,    18,    40,     4,   -10,    16,   -13,   -40,   -44,   -57,   -78,    -2,    -1,    -1,   -20,    51,     3,   -13,    -1,    47,    66,    67,    71,     7,    13,    17,    34,    38,    64,    21,   -23,   -37,     2,    11,   -11,    -1,   -87,   -67,   -35,    -8,    -5,     2,     7,   -28,   -27,    47,    42,    43,    48,    60,    34,   -10,    18,    -2,    29,    40,    48,    44,    29,    38,    43,    -1,   -44,  -121,   -75,   -26,   -16,     2,   -10,     9,     0,   -29,   -66,    46,    31,    37,   -51,   -51,    12,    10,   -20,   -56,   -47,   -24,    21,    11,   -10,   -18,   -17,   -44,   -42,   -28,   -10,     3,     3,     0,    -9,     0,     5,    -3,    -2,   -19,    -7,     3,   -16,   -33,   -41,   -44,   -23,   -41,   -45,   -30,    -1,   -10,   -28,   -37,   -28,   -21,   -11,    -2,     3,    -5,    -8,    -6),
		    64 => (   -3,    -4,   -10,    -2,     5,    -6,     7,     6,    -3,    -2,    -9,    -8,   -15,   -19,    -6,    -8,     3,   -10,    -8,    -4,    -2,    -5,   -10,    -2,    -1,    -2,     2,     8,    -2,    10,    -6,     8,     3,    -5,   -36,   -28,   -21,   -14,   -40,   -31,   -10,   -36,   -15,   -25,   -18,     2,     6,    -2,    -8,    -5,    -4,   -13,     1,    -5,    -3,    -2,     6,    -2,    -1,     8,    -6,    -2,   -46,   -38,   -47,   -74,   -67,   -79,   -48,   -35,   -15,   -16,   -13,   -11,   -17,   -10,   -33,    -8,   -15,   -18,    -8,     2,    -5,     6,     0,    -7,     6,     4,   -22,   -28,   -10,   -22,   -70,  -102,   -56,    -4,   -24,   -60,   -44,     1,    -1,   -12,    47,    16,   -24,    -8,   -31,     2,    23,    -4,     9,     0,    -8,     0,   -11,   -19,   -29,     0,     7,   -11,   -23,   -38,    -1,   -14,   -27,   -37,   -28,   -36,   -24,   -33,    -2,    23,   -25,   -19,    15,    62,    24,    22,   -33,   -17,    -2,     8,    -3,   -13,   -13,   -39,    -9,   -38,    20,     0,    31,   -62,  -108,  -139,  -117,   -34,    47,    34,   -59,   -61,   -35,   -43,    -9,    44,     4,    28,   -33,   -10,     8,     7,    -9,   -45,   -36,   -12,    32,    14,    20,    42,   -44,  -107,  -125,  -187,  -133,   -23,    13,    41,   -16,   -85,   -28,     6,    40,    52,   -22,   -54,    13,   -24,    -9,   -46,     0,   -38,   -35,     1,    -6,     1,    43,    64,    23,   -65,  -157,  -215,   -70,    37,    26,    32,   -75,   -10,    24,    49,   105,    29,   -70,   -64,   -16,   -61,   -24,   -37,   -14,   -48,   -41,   -18,    22,    -1,    16,    64,    27,   -41,  -188,  -139,   -38,    14,    50,    -5,   -65,   -44,    12,    40,    11,    30,   -79,   -11,   -49,   -51,     4,   -17,    -5,   -55,   -36,   -10,   -36,    30,    46,    45,    33,   -23,   -70,   -55,   -21,    -1,    19,   -19,   -19,     1,    -3,     7,     2,    43,   -32,   -20,   -34,   -20,    -5,     9,     1,   -56,    -6,     1,   -10,    22,    31,    69,    46,     5,   -67,   -85,   -14,    35,    11,     3,     5,   -10,   -32,   -30,   -25,    -7,    25,    16,   -18,   -30,     6,   -16,   -10,   -36,    11,    20,    14,     6,    48,    66,    26,   -30,   -60,   -58,   -41,   -15,    -9,     3,   -31,   -15,     6,   -11,     6,   -23,   -10,    25,   -24,   -57,     9,   -16,    10,   -74,   -28,    -7,    26,   -14,     9,    43,    22,    -6,    -8,    10,   -12,    15,    -3,     4,    -6,    13,    37,    -7,     4,   -58,   -50,   -11,   -27,   -54,    -7,    -1,   -19,   -48,   -55,   -38,    28,    20,   -12,    47,    19,     0,    -1,    24,     8,    26,    -2,     9,    32,    57,   -12,    10,    10,   -76,   -76,    -3,   -31,     8,    -9,    15,   -58,   -14,     4,   -21,   -25,    16,   -38,   -25,    -3,    -9,     4,   -12,    16,    47,    12,    36,    31,     8,    12,    33,   -28,   -83,   -63,    11,    65,     7,     7,    -4,    39,     6,    48,    -5,    40,    -4,    42,   -29,   -21,   -35,   -41,     1,   -22,    32,    10,     2,   -13,     7,   -58,   -10,    14,    34,   -49,    23,    83,    10,     4,     2,   -29,    28,   -10,   -44,   -37,    25,    -7,    13,    -8,   -21,   -13,   -13,   -39,    13,   -11,    -5,    -3,   -31,   -87,     1,    11,    -6,    57,    72,    24,    -9,     8,    -3,   -15,     5,     4,   -33,   -29,    15,    13,     5,   -18,   -25,   -34,   -24,   -47,    15,     2,   -18,     0,   -46,   -38,    30,    -9,    14,    27,    78,    62,   -20,    -4,    -1,   -13,    -7,    -7,   -43,   -33,     8,    -4,     0,   -37,   -62,   -63,   -20,   -30,    20,   -31,   -22,    13,   -15,   -24,    -7,   -13,     6,   -29,   -14,     4,   -17,     9,   -11,   -27,    12,   -20,   -37,   -12,    18,   -24,   -22,   -33,   -58,   -52,    -1,    -8,    30,    -6,   -26,    43,   -16,   -55,   -20,    -4,   -23,   -30,   -40,     2,   -19,     8,    -1,     0,   -27,   -36,   -36,   -35,    25,   -16,   -17,   -44,   -23,   -63,   -25,   -13,     5,    13,    -8,     6,    16,    -8,    11,    21,     4,   -10,   -64,    -1,     0,     7,     8,   -33,   -39,     0,    -1,   -13,    25,    10,   -21,   -38,   -93,   -55,    -9,    41,     9,   -10,   -13,    -3,    13,     3,     0,   -19,    36,    -2,   -69,   -33,    -4,     5,     3,     4,   -24,   -37,     5,    11,    -7,    18,   -33,   -55,   -64,   -42,   -10,    10,    10,   -22,   -47,   -11,    45,     4,    14,    22,    56,   -28,   -29,    19,    -1,    -6,     6,    -8,    -9,   -22,   -28,     3,    -5,   -19,    -6,   -22,   -73,   -13,    18,    14,    -7,   -24,   -49,    22,    34,   -25,    50,     3,   -25,   -58,    21,     7,    -2,    -1,    -4,    -4,     2,   -28,   -23,   -22,   -35,     9,    -9,   -25,   -29,   -21,   -10,    21,    27,     1,     0,    15,    11,    13,    19,    41,   -28,   -68,     6,   -18,    10,    -3,     8,    -4,    -1,   -12,    -5,   -23,   -17,    19,   -12,   -36,   -34,    -2,    25,   -55,   -30,   -27,    19,    19,    10,    41,    23,   -21,   -24,   -30,   -17,   -13,     6,     8,   -10,    -5,   -20,   -10,   -20,    -9,    -3,    10,     5,   -29,   -17,   -17,  -112,  -123,  -116,   -60,    -8,   -27,   -67,   -88,   -81,  -100,    -5,   -28,     0,    -8,    -2,     7,     6,    -2,    -4,     7,     1,   -16,   -36,   -40,   -23,   -18,   -40,   -39,   -35,   -40,   -14,   -42,   -67,   -50,   -39,   -46,   -51,   -55,    -1,     5,    -3,    -1,    10),
		    65 => (   -8,     7,     3,    -3,    -7,     0,    -1,     6,   -10,    -9,     3,    -4,    -6,    -1,     3,     4,     4,    -4,   -10,    -8,     6,   -10,    -7,     5,    -8,    -6,    -9,    -5,    -1,    -1,    -8,    -4,     1,    -2,    -6,     8,     9,    -3,   -13,    -3,   -10,   -12,   -15,   -18,   -20,   -16,   -19,    -2,    -8,    -4,     6,     6,     3,    -7,    -2,    -9,    -1,     5,   -10,     8,   -10,     0,     1,    -5,   -16,    -5,   -10,   -46,   -44,   -51,   -62,   -31,   -37,    38,     3,    20,    49,   -14,    -3,   -14,   -19,   -12,    -8,    -1,     3,    -9,    -3,    -3,     8,    -8,   -20,   -16,   -26,   -39,     9,   -15,   -36,   -13,   -12,    15,   -34,    34,    27,    26,    61,    66,    41,   -47,   -37,    18,    65,     5,    -3,     7,   -23,   -13,   -15,   -21,   -56,   -27,   -50,    39,    38,    -1,     6,   -56,   -33,   -16,   -63,   -16,    34,   -27,   -27,    16,    -3,   -23,    -8,    47,    38,   -36,    -5,     8,   -33,   -24,   -19,   -32,  -104,  -111,   -25,    42,     9,    -5,    22,    51,   -10,  -107,   -40,   -29,   -42,   -23,    45,    25,    25,   -26,   -26,    30,    48,   -16,    -7,    -9,    42,   -21,   -36,   -79,  -102,  -108,   -56,   -11,    29,   -15,    54,    52,    -5,   -32,   -36,     0,    -8,    16,    51,    20,    43,    -3,     3,    88,    91,    30,     9,    -9,    40,   -47,   -27,   -27,   -91,   -88,   -51,    30,     5,    -4,    43,    35,   -30,    27,    46,    47,    53,    57,    64,    15,    40,    -4,   -24,    38,    91,     2,    -3,   -21,   -39,   -39,   -22,   -95,   -80,   -41,    -8,   -11,   -29,   -23,    -4,   -25,     4,    28,    42,    52,    91,    69,    53,    -9,    15,    33,    -4,   -11,    49,    27,     5,    -3,   -63,   -69,   -64,   -61,   -38,   -34,   -50,     0,   -14,   -17,   -33,   -22,   -51,   -50,   -26,    53,    22,    -7,   -41,   -32,    -5,   -15,   -23,    38,     7,    46,     8,   -12,    -5,   -11,    11,   -36,   -13,   -71,   -29,    22,   -30,     1,     5,   -30,   -65,  -149,  -156,  -122,   -97,  -134,  -116,   -42,   -54,  -120,   -53,     4,    52,    58,    -6,    -3,     1,   -12,    69,     1,   -70,   -44,   -25,     2,     2,   -21,     1,   -22,   -36,   -96,  -123,  -173,  -158,  -146,  -162,   -99,   -80,   -99,   -64,   -35,     9,    51,     3,    -6,     2,    18,    33,   -30,   -60,   -24,   -19,   -12,    21,     7,    -2,    50,     8,    -7,   -27,   -67,   -43,   -66,   -78,  -107,  -107,   -81,   -65,   -28,    -7,   -26,    -2,    -9,     3,    30,    16,   -22,   -11,     5,   -23,   -35,   -14,   -20,    -9,    24,    30,    23,   -24,   -27,   -32,   -37,   -11,   -85,  -139,   -83,   -67,   -22,    -4,   -27,     1,   -16,   -13,    43,    13,   -37,   -17,    21,     9,    14,    -1,    12,    16,    -5,   -18,    11,   -25,   -14,   -26,    -3,    40,   -11,   -31,   -25,   -25,   -15,    -7,    -7,    14,   -15,   -49,   -29,    19,     2,    32,   -33,   -18,    32,    -5,     2,    11,   -25,    -8,   -16,    15,   -20,    -2,   -23,    19,    51,   -23,   -13,    20,     4,   -13,   -31,     4,   -11,   -29,   -27,   -13,    -7,   -35,   -53,    -2,     6,    20,    26,     8,    26,     2,   -32,    -3,     9,   -51,     7,    -9,   -22,   -51,   -64,    -2,   -30,   -50,   -34,     0,   -10,   -39,     0,     7,   -41,   -47,   -17,   -39,   -12,    36,    32,    16,    37,   -22,   -16,   -14,   -13,   -18,     5,    22,   -28,   -40,   -78,   -11,   -36,   -10,   -44,     2,   -11,   -34,    15,    14,    -5,   -64,   -92,   -62,   -79,   -41,    28,   -12,   -11,   -53,   -45,    32,    14,    10,     0,    42,   -36,   -27,    -2,    11,    -8,   -43,   -25,     9,     1,   -26,   -43,    66,    -2,    -1,   -43,   -49,  -110,  -100,  -114,   -40,     7,   -29,   -63,     1,    29,    10,   -12,    38,   -36,   -32,    27,    29,   -22,    -6,   -13,     2,   -12,   -19,   -22,    12,    32,    11,     7,   -15,   -60,    -8,   -44,   -78,   -10,   -12,    13,   -27,     8,     9,    31,    27,   -14,    -6,    18,    -6,   -11,   -19,     8,     1,    -7,   -47,    -3,    49,    28,     5,     6,    -2,    15,    22,    -5,    -7,    24,     9,     7,   -22,   -23,    10,    42,     9,   -26,    29,    21,   -18,    -9,   -32,     2,     9,     6,   -54,    51,    21,   -31,   -15,   -25,    16,    63,    49,    39,     9,   -30,    18,   -21,   -12,    16,    -7,    -2,    11,    -3,    -5,    59,    -5,   -16,    -8,    -9,    -2,     5,    23,    63,    57,    28,    40,     6,     9,   -37,    14,    31,    13,     3,    -9,     6,   -32,   -16,    -9,     8,    10,    -1,    17,    63,   -13,   -40,     7,    -7,     9,     8,   -33,    13,   -17,   -17,    -3,     3,   -15,     5,     9,   -19,   -12,    -7,     4,     2,   -30,   -19,    24,   -14,   -35,    14,    82,    19,    31,   -46,   -25,    -4,    -9,   -10,    -9,    73,   -55,   -56,   -22,   -35,   -53,     6,   -31,   -25,     7,    41,   -13,   -12,   -89,    15,    18,     9,    26,    67,   103,    50,    30,     1,     2,     0,     1,     5,     0,    -5,    -9,   -18,   -16,   -18,   -27,   -50,   -12,    37,    43,    23,   -85,   -99,   -83,   -86,   -41,    21,   -31,    28,    24,   -10,    -8,     0,    -5,    -7,     9,     0,    -5,     1,     1,    -9,     3,    -6,   -10,   -16,    -1,     4,     9,    16,   -21,    -3,    -3,    -2,   -13,    -6,     4,   -12,   -25,   -10,    -6,    -3,    10,     2),
		    66 => (   -1,     4,     2,    -6,     7,     8,    -3,    -4,     5,    -9,    -2,     3,    34,    40,     5,    -7,    -3,     0,    -8,    -6,    -3,     7,     4,     7,     8,    -5,     1,     0,    -2,     8,    -5,    -9,     1,     2,    19,    18,     9,     3,    44,     5,    19,    48,   -21,   -19,   -10,     9,    27,    42,    46,    38,    35,    31,    -2,    10,    -2,     0,    -2,    -8,     2,   -12,    14,    31,    20,    -5,    11,    37,    34,    34,    23,    34,    29,   -14,    29,    31,    41,    66,    56,    31,    94,    63,    48,    38,     1,     3,     8,     5,   -56,    30,    -6,    56,    62,    58,    80,    81,    94,    95,   122,    78,   107,    75,    19,     8,    10,     8,   -31,   -39,   -27,    -2,    38,   -77,   -66,     2,     6,    -7,   -43,     4,    31,    51,    55,    77,    39,    83,    72,    39,    71,    12,    82,    68,    18,    31,    14,    43,    51,    27,   -14,   -21,   -25,   -52,   -21,    60,    -9,    -5,   -22,   -45,    70,    31,    43,    50,    31,    36,    64,    15,   -36,    33,    68,    35,     9,    50,     6,   -20,    12,   -43,    -8,     5,    56,    26,    53,    19,     4,     1,     1,     4,    53,    19,    57,    32,    -8,    24,   -14,   -32,    19,    16,    17,     7,     4,     1,   -64,    15,    -6,   -37,   -38,   -33,    -8,    21,    49,    69,     4,    -8,    -4,   -19,    55,    38,    21,    19,     5,   -19,   -31,   -14,   -45,   -60,    22,   -21,    -9,   -20,   -20,     6,   -19,   -11,   -14,   -12,    21,     6,    43,    47,    -6,   -22,   -28,  -105,    61,    21,    11,   -23,     2,    32,   -28,   -31,   -19,   -36,     1,   -48,   -85,   -37,   -21,    -8,    20,    21,   -20,   -38,   -38,   -85,    -7,   -66,     0,    -9,   -36,   -57,    49,   -11,   -34,   -23,     7,   -19,   -29,   -37,   -54,   -64,     0,     3,   -35,   -83,   -14,   -16,    -8,    40,    -7,    -9,   -57,  -103,   -64,   -57,    -6,    -9,   -41,   -32,    14,     5,   -36,   -38,    -9,   -23,   -14,   -53,   -65,   -30,     8,   -26,   -71,   -44,   -60,   -44,     8,     5,   -48,   -41,   -71,   -76,   -64,   -63,    -2,   -10,    -7,   -64,    14,     9,    -3,    -9,   -31,   -12,   -27,   -50,     5,    -5,   -10,   -43,   -37,   -33,   -38,   -21,   -19,     5,   -43,   -10,   -33,   -65,   -69,   -48,    10,    -8,   -30,   -60,   -10,    16,    45,    13,   -16,    15,    -3,     8,   -15,    25,   -33,   -22,   -54,   -34,   -48,   -36,    26,    19,   -30,    29,    42,    -4,   -93,   -47,    -3,     6,   -21,   -53,   -24,    20,    -6,   -24,   -23,    42,    52,    35,    34,    17,    23,     8,   -12,   -61,   -17,    25,    29,    31,   -20,    32,    22,   -30,   -97,    -1,     0,    -4,    -9,   -51,   -72,    24,   -30,   -50,    15,    18,    51,    51,    54,    28,    12,   -37,    -7,   -35,    15,    18,     9,    23,    24,   -27,   -13,    51,   -78,   -16,     0,    -3,   -31,   -35,   -80,   -29,   -27,    -9,   -24,    -8,    13,    27,     0,    62,    41,   -25,   -27,   -66,     4,    34,    -5,    10,   -47,     6,     1,    44,   -33,   -94,     7,    -1,   -46,   -36,   -18,    15,    14,    21,   -23,    28,    27,    11,   -18,   -33,   -22,   -20,   -23,   -30,    44,    49,   -20,   -16,    15,    -3,   -15,    34,   -50,   -77,    -9,     3,   -54,   -54,   -36,    46,     3,    18,   -11,   -36,   -20,    -9,   -19,   -32,     6,    19,    19,    34,    27,    32,    26,   -12,   -10,   -22,   -11,    30,   -47,  -109,     8,    -7,   -52,   -84,   -15,    -6,   -35,     8,    -4,    10,    34,   -57,    -4,    -7,     0,   -39,     4,    32,    83,    67,     7,   -26,     2,    14,    10,    51,     4,   -47,     7,     1,   -61,   -68,     8,    25,    22,    -8,     4,     3,    63,    63,    36,    15,    10,    18,     2,    46,    -2,    68,    -6,    -4,   -11,   -26,   -54,    16,   -32,    -2,     1,    -3,   -56,   -85,    -3,    -4,     2,    26,     9,    15,    54,    58,    49,   -31,    13,    14,    12,    32,    35,    31,    32,    -3,    -6,   -62,   -74,   -21,   -20,    -1,    -5,    -9,   -72,   -76,   -58,   -68,   -19,    45,    56,     0,    29,     3,    83,    39,    16,     9,    67,    42,    36,    22,    14,   -22,   -15,   -66,   -33,    -3,    -6,   -11,     1,     5,   -52,   -60,  -107,  -134,  -179,     0,     2,    33,    17,    10,     4,     1,     5,    46,    53,    77,    48,     6,    16,    15,   -55,   -47,  -119,   -31,   -13,    -8,    -2,     9,     8,   -65,   -81,   -92,   -85,   -12,   -22,     4,   -35,    10,    40,   -11,    20,    43,     3,   -36,    10,     2,     6,    27,   -66,   -82,   -79,   -54,   -64,    10,    -9,     4,    -5,   -10,   -26,   -30,   -45,   -86,  -117,  -153,  -105,  -135,   -66,   -66,   -42,    11,    22,    31,    69,  -105,   -16,   -56,   -48,   -44,   -34,   -22,    -9,     0,     5,     6,    -3,    -4,    -9,   -19,   -34,   -33,   -24,   -32,   -38,    14,    30,   -19,   -17,   -28,   -49,   -48,   -27,   -78,   -72,   -14,   -38,   -38,   -31,     8,    -4,     8,     3,     8,     1,    -2,    -9,   -14,     6,   -11,    -4,   -11,    -9,   -17,    -6,     3,    -5,   -15,    -3,   -10,    -1,   -11,    -9,     9,    -9,   -10,     5,     7,     4,     8,     0,     5,    -7,     9,     3,     3,    -1,    -1,    10,    -4,    -5,    -7,     4,     5,    -6,     0,    -4,    -9,     1,     3,    -9,   -11,    -5,     5,    -9,    -2,     3,     1),
		    67 => (   -7,    -7,     7,    -7,     1,     3,     4,     7,    -9,    -8,     7,     5,     8,     2,    -2,     1,    10,     5,     7,     9,    -4,    -8,     7,     9,     3,     8,    -8,   -10,     5,    -6,    -2,     0,     4,    -3,     9,    -5,     6,     4,    -3,   -11,   -10,   -15,   -16,   -37,   -37,   -24,    -3,     2,     2,    -7,    -4,    -6,     6,     6,     2,     6,    -6,    -6,     9,    -6,     1,    -3,   -10,    -5,   -16,    12,    -8,   -35,   -57,   -25,   -25,   -24,     8,    -3,    -8,    -9,   -11,   -12,    -3,     9,     2,    -2,     2,    -6,    -8,     7,    -7,     0,   -15,   -30,   -34,   -56,   -25,   -10,   -24,   -37,   -68,   -69,   -50,   -49,   -32,   -25,   -11,     1,    -9,     8,   -20,    -6,   -15,   -13,     7,     0,     9,     0,     0,    -7,   -25,    -6,   -42,   -43,   -60,   -73,  -106,     4,     9,     4,   -16,   -50,  -117,   -88,   -65,   -69,   -51,     6,   -33,   -42,   -45,   -28,   -12,    -8,    -5,    -7,    -2,   -27,   -38,   -15,   -78,     3,    77,    15,   -15,     1,    25,   -10,    28,     8,    11,    -1,    60,    -3,   -40,   -20,   -17,   -36,   -61,    -9,   -14,    -5,    -4,     3,    28,   -20,   -20,   -16,   -50,    21,    34,    54,    25,    -9,   -13,   -15,   -17,    24,    11,     2,    37,    15,   -74,   -33,     4,   -40,   -40,   -28,   -29,   -15,     7,    22,    31,    -1,    17,     0,    21,    19,    28,    21,    -7,   -21,   -39,   -42,   -46,    -4,    38,    39,    30,    48,    72,    13,   -30,   -32,   -54,   -31,   -28,   -16,   -41,    12,    77,     5,    31,    22,    13,    50,    45,     4,    -9,   -18,   -12,   -35,     5,    45,    12,    11,    19,    24,    48,    26,    -6,   -70,   -45,    -9,   -20,   -15,    14,    16,    18,    38,    36,   -55,   -14,     3,    16,    -4,    14,   -30,   -19,    14,     2,   -12,    15,    41,   -13,   -11,    22,   -36,   -21,   -43,   -27,    -6,   -39,    15,    12,     5,   -12,    10,    53,   -14,   -13,     8,   -21,    19,    12,   -35,   -67,    12,    -5,     8,     7,   -10,     1,    11,   -13,   -49,   -13,   -36,   -37,    -6,   -27,     2,    13,    14,    -8,   -39,     0,     7,   -19,    30,    13,   -21,     7,    -1,   -66,   -44,    -1,    59,    -5,    -2,     0,    -5,   -40,   -28,   -38,   -78,   -42,   -46,   -36,    14,     7,     7,   -31,    -9,   -31,    -8,   -32,    28,    -6,   -44,   -25,   -73,   -76,   -52,   -31,    38,   -18,   -52,   -17,   -68,   -40,   -40,   -74,   -72,   -81,   -21,   -24,     5,    -5,    26,    29,   -13,    -9,    -9,   -26,    -2,     4,   -30,   -42,   -69,  -138,   -90,   -49,   -10,   -26,    -3,   -20,   -64,   -56,   -56,   -67,   -88,   -77,   -10,   -47,   -23,    -2,    32,    10,    33,    -4,    24,   -54,   -28,   -53,   -82,  -145,  -114,   -74,   -54,   -41,     1,   -40,    13,    33,     8,   -23,    16,   -47,   -58,   -22,   -12,   -38,   -15,     7,    -4,    -1,    26,    20,   -12,   -37,  -100,   -61,   -55,   -79,     8,   -14,   -10,   -48,    -2,    -4,    37,    42,    11,    25,    23,   -11,     5,     8,    20,   -12,   -18,     4,     4,     2,   -26,   -17,     0,   -63,   -31,    55,   -19,   -17,    50,    16,    -2,   -10,    42,    17,     8,    38,   -24,    -7,   -41,   -26,   -12,    -9,   -62,   -29,    -8,     8,    -1,   -29,   -24,   -37,   -70,   -35,   -25,   -14,     3,   -43,     4,   -11,     4,   -13,    16,    12,    36,    23,     3,   -70,   -74,   -60,   -50,   -20,   -96,   -53,   -67,    12,     3,    13,   -35,   -31,   -10,   -26,     3,   -22,    12,    -4,     5,   -42,    30,    12,    52,    -5,    57,   -29,    20,    32,     6,   -49,   -62,   -37,   -74,     7,   -47,    -4,     5,     3,    -4,    -9,   -67,   -25,   -25,    23,   -19,   -18,   -48,   -22,   -21,    49,    69,   -31,   -27,   -23,    20,    34,    37,   -23,    -7,    13,   -31,   -40,   -35,    -1,    27,   -14,    -3,   -12,   -54,   -42,    -2,    14,    20,   -11,  -101,   -30,   -13,    20,    16,   -29,   -53,   -22,    -9,    30,    -4,   -25,   -83,   -43,   -23,   -42,     7,   -12,     7,   -13,   -20,   -16,   -57,   -77,   -71,    16,   -20,   -33,   -54,   -11,     3,    29,    11,    43,   -57,   -24,   -36,   -22,     8,   -28,   -98,   -54,   -53,    -3,    -3,   -15,     5,    -8,    -5,   -13,   -47,   -63,   -62,   -36,   -47,   -25,   -53,   -31,    36,     8,    30,     9,    16,   -39,   -20,   -28,   -83,  -125,   -89,   -53,   -30,   -50,     3,    -1,    10,   -13,   -33,   -69,   -72,   -63,   -96,   -81,  -112,   -77,   -66,   -38,   -18,   -18,     2,   -13,   -59,   -88,   -61,   -57,   -60,   -56,   -44,    14,   -30,   -45,    -8,    -9,    -8,     6,     0,   -27,   -71,   -84,   -83,  -121,  -115,   -85,   -57,   -15,    -1,    13,    43,    -9,   -15,   -80,   -50,    -7,   -22,    -6,   -38,   -25,   -26,    -7,    -3,    -5,     0,   -46,     0,     6,   -30,   -46,   -65,   -66,  -104,   -63,    17,   -28,   -24,    -8,    54,     5,    14,    -3,    27,    37,    26,   -17,   -31,     1,    -4,    -7,    -4,     1,    -5,     0,    -3,   -23,   -25,    -7,    30,    17,    19,   -25,   -18,    26,    39,    21,     8,    -1,    14,   113,    93,    57,    16,   -11,   -16,    -5,     0,     0,     0,    -6,    -3,    -1,     5,    19,     4,    -4,   -17,     1,    40,    56,    34,    25,    25,    10,    44,    39,    67,   100,    63,    29,    -5,   -19,     9,     2,    -8,    -5,    -9),
		    68 => (    7,     9,     7,     2,    -5,    -8,     4,   -10,     3,    -5,    -9,    -1,    -3,     4,     1,     6,     6,     3,    -3,     2,     3,     3,    -4,    -2,    -1,    -9,    10,     3,     8,    -5,    -5,    -7,     9,     6,     8,    -8,     3,     1,     7,    -3,     3,     0,    -2,    -8,   -42,   -36,     2,     0,    -5,   -10,    -9,     4,     2,    -3,     6,    -4,    -3,    -9,    -7,    -6,   -10,     1,     3,    -9,    10,   -12,   -23,    -6,     0,    -7,     5,    -4,   -21,    -3,     1,    -1,    -8,   -22,   -10,   -20,    -3,    -8,     9,     7,    -8,    -4,     1,    -3,    -8,   -18,   -11,   -21,   -16,   -15,    -1,     0,    -8,     3,   -33,   -23,    -8,    -3,    12,    -8,   -21,     4,     9,     8,    -8,     2,   -16,     6,     9,    -5,     3,   -15,   -10,   -10,   -29,   -30,     7,     2,    -6,    30,    29,   -21,    -2,   -51,   -42,    -9,    16,     3,    12,   -18,   -20,    -2,   -13,     5,     1,     1,    -9,    -9,     0,   -17,   -46,   -55,    -2,    -8,     2,     2,   -24,   -12,   -24,   -22,     6,   -12,   -33,   -13,   -17,   -21,    -7,   -16,   -25,   -14,    -8,    21,     1,   -16,    -9,     2,   -20,   -40,    -7,     8,    -8,    22,    -6,   -20,   -32,   -49,   -19,   -45,   -26,    -1,    -4,     3,   -11,   -17,   -13,   -28,   -11,    -7,    -8,   -15,    -9,     0,     5,    -5,   -15,     1,    10,    47,     9,    12,     5,   -10,   -12,   -29,     7,     3,    11,    17,    14,     9,     4,    10,   -29,    -9,     9,     1,    14,    -2,     3,    -9,    -3,   -21,    -7,    38,    58,    63,    24,    -8,   -36,   -26,    -8,    13,     6,     9,    -4,   -24,   -33,   -18,   -18,   -17,     4,     7,    11,   -12,    -9,     6,   -17,    -3,     3,   -26,   -34,    31,    49,    57,    22,   -21,   -52,   -32,    19,   -33,   -32,   -18,   -25,   -48,   -42,   -11,   -20,    21,    25,    27,     7,    -2,     3,    28,   -15,   -12,    -7,   -17,   -34,    19,    14,    45,    38,    24,   -25,     7,    22,    -6,    -1,   -17,   -19,   -26,   -21,     1,   -16,     1,    10,    -3,   -20,   -21,    -3,   -28,   -14,   -15,    -1,    -4,   -44,   -23,   -19,    -3,    37,    47,    32,    47,    34,    10,   -10,   -18,   -26,   -14,   -14,   -19,   -38,    -4,   -11,   -10,     7,   -11,   -21,   -15,    -1,   -37,     3,     4,   -26,   -57,   -44,   -10,     5,   -19,    18,     9,    31,     3,     0,   -41,   -42,     0,     0,    -9,    -7,   -28,   -27,    20,     8,   -10,   -16,   -26,   -28,   -44,     2,   -12,   -40,   -62,   -24,   -38,   -38,   -39,   -38,   -33,   -19,     5,     4,   -24,    11,    13,     4,   -27,   -24,   -45,   -35,    -7,    -5,    -9,   -26,   -44,   -27,    13,   -17,   -11,     9,   -61,   -27,   -24,   -34,   -50,   -46,   -69,   -34,   -47,   -28,    -2,   -11,   -36,   -38,    -4,     1,   -16,   -38,   -15,    -6,    -8,   -31,   -14,   -70,    -8,     2,     9,   -13,    13,     2,   -13,   -25,   -44,   -28,   -40,   -29,   -16,   -22,    -2,    -4,   -13,    -3,   -13,    -4,   -23,    -3,   -27,   -21,   -23,   -27,    13,   -25,   -29,     6,   -15,    -4,    16,    -1,   -14,   -32,   -19,    -8,   -36,    -1,     9,     1,   -19,   -41,   -44,    15,    19,   -20,   -15,    -5,     0,     1,   -19,   -19,     7,   -32,   -23,     9,    -1,    -1,    25,    -8,   -24,   -21,   -16,   -26,   -25,    26,    29,    -4,   -29,   -31,   -48,   -26,    14,     2,   -22,   -16,     9,    19,   -27,   -13,   -15,    -9,   -14,    -2,    -9,    -6,     4,   -19,   -15,   -22,   -16,   -29,   -25,    10,     2,    13,     2,   -41,   -33,   -32,    25,     9,   -10,   -37,   -17,    32,    -9,   -16,     6,    -3,   -29,     5,     4,   -11,    -4,   -23,    -9,    -8,   -15,   -56,    -3,    23,    24,    -4,     3,   -28,   -34,   -34,    -6,    28,    10,   -11,     5,    17,    20,    -1,     5,   -21,   -23,    -7,    -3,   -20,   -16,   -19,   -12,    -6,   -18,   -36,    -6,    11,    31,    13,   -36,   -44,   -29,   -42,    -9,    15,     3,    -1,    -3,    31,     9,    -9,    -3,   -26,     1,   -14,   -16,    -7,   -27,    -9,    -9,   -35,   -26,   -21,   -16,   -13,    10,    14,    -8,   -22,   -21,   -39,     5,    14,     6,     5,     7,    32,     0,   -11,   -13,   -13,    -3,   -31,   -13,   -12,   -19,   -13,   -24,   -19,   -14,   -21,   -28,    -6,    -6,   -13,    -9,   -19,   -14,   -24,    13,    -7,    -5,     1,    23,     9,    -9,   -34,   -13,    -4,     2,     8,     8,    -1,   -16,   -16,   -30,   -29,   -21,   -11,   -22,    -4,   -34,   -15,    19,   -15,     1,    13,     3,    -9,     2,    17,    30,    11,   -18,    -2,     0,   -44,     0,    -7,     9,   -12,     2,    -8,   -20,   -18,     9,   -15,    -4,     0,   -30,   -27,   -30,     9,    23,    26,   -24,   -41,   -25,    -2,   -26,   -30,   -10,   -11,   -14,    -5,     8,     4,    -7,   -17,   -15,   -15,   -17,   -22,   -26,   -18,     2,    25,   -17,   -23,   -16,     0,     9,     2,    -6,   -20,   -16,   -30,   -24,     0,    -3,   -11,    -6,   -19,    -8,     0,    -4,    -3,    -5,     0,   -16,   -13,   -27,   -13,   -30,   -27,   -25,   -28,   -21,   -37,   -32,   -10,    -1,     1,   -41,   -49,    -4,   -32,     1,     4,     5,     0,     2,    -2,     9,     8,     2,    -3,     4,    -2,    -6,    -5,   -16,   -14,    -6,     1,   -13,   -11,    -7,   -16,   -13,   -27,    -6,    -4,    -5,    -9,    -7,    -1,     8,    -8,     2),
		    69 => (   -7,    -8,     6,     7,     7,     8,     0,    10,    -9,     7,     9,     8,    -3,     4,     1,     4,    -8,    -6,    10,    -6,     2,    -4,     3,    -2,     1,    -7,    -1,     3,     2,     6,     9,    -8,     2,    -1,    -6,   -17,   -22,   -19,   -16,   -26,   -31,   -46,   -24,   -53,   -46,   -48,   -24,     2,     6,    -8,   -25,     2,     8,    -8,    -7,    -7,    -7,    -3,    -8,   -36,   -41,    -8,    -7,   -43,   -54,   -23,   -27,   -39,     3,     0,  -113,   -63,   -58,   -36,   -64,   -46,   -85,   -96,   -70,   -58,   -35,   -18,     8,     2,     2,    -2,    -4,   -47,   -61,   -54,   -34,   -58,  -127,  -159,  -215,  -192,  -128,  -166,  -153,  -166,  -217,  -188,   -60,   -81,  -133,  -117,   -97,   -55,   -48,   -30,    10,     5,     9,    -7,   -27,   -42,   -69,   -88,  -126,   -88,   -98,  -108,   -66,   -18,     8,   -10,   -35,   -35,   -30,   -62,  -115,  -225,  -144,  -119,  -118,   -62,   -53,   -86,   -61,     5,    -4,     2,   -27,   -39,   -32,   -52,   -54,   -35,   -79,    13,    14,     5,    29,    62,    20,    24,    52,    52,    -7,   -32,   -66,   -27,  -131,   -55,   -82,   -85,   -59,   -15,    -5,     9,   -26,   -86,   -63,   -79,   -41,   -25,    -3,    40,    41,   -20,   -16,    60,    26,    62,    97,    61,    14,    21,   -14,    -7,   -17,    15,     3,   -28,   -64,   -75,     1,   -30,   -55,   -72,   -46,   -84,   -11,    -8,   -15,    16,    15,   -11,    35,    73,    67,    57,   117,    71,     0,    22,    36,    -4,    19,    19,     0,     7,   -70,   -57,   -51,   -65,   -51,   -57,   -63,    -6,    23,   -11,     0,    19,     7,     5,    48,    42,    65,    98,    78,    54,    48,    59,     5,    24,    16,    38,    40,     3,   -67,   -37,    -9,   -45,   -67,   -70,    42,    16,    40,    20,    23,    43,     8,   -12,    19,    56,    52,    33,    24,    19,    16,    13,    47,     0,    -3,   -17,   -21,   -71,   -87,   -58,    -4,   -31,   -95,   -44,    42,    43,     2,     8,    -6,    -7,     3,    -3,    32,    22,    12,   -40,     1,   -24,    -1,    -2,    12,   -44,   -26,   -21,   -55,    37,   -91,   -36,    -4,  -146,    -1,   -31,    12,    49,    21,   -17,   -43,   -12,   -12,   -34,    -1,   -56,   -47,   -50,    -2,    13,   -37,   -18,    32,   -21,   -63,   -40,   -53,    -6,   -76,   -30,     2,   -15,   -11,   -29,    34,    20,    16,   -21,   -49,   -49,   -18,     1,   -42,   -54,   -26,   -41,   -22,    11,   -30,   -46,    11,   -34,   -30,    -5,   -63,  -106,   -64,   -44,   -10,   -31,   -47,   -33,    16,   -15,    13,     9,     2,   -30,    -7,   -30,     3,   -17,   -25,   -47,    11,     1,   -15,   -24,   -32,     2,   -38,   -36,   -27,   -77,   -47,   -13,   -17,   -28,   -29,    -7,    22,   -11,    -6,    13,     2,    -5,     4,   -18,    25,   -46,   -30,    18,     4,     0,    21,    17,    -5,   -31,   -44,   -89,   -40,   -93,   -55,     0,     0,    -4,   -65,   -28,    11,     8,    24,     6,    33,    21,   -33,   -47,   -40,   -13,    24,    19,    37,    19,    31,    50,    60,    23,    11,   -65,   -37,   -89,   -20,   -59,     5,   -15,   -45,   -29,     1,    37,    35,   -10,    16,     4,   -11,   -53,   -55,   -15,    43,    30,     5,    41,   -13,    30,    47,    10,    -2,   -45,   -17,  -112,   -60,   -65,    -2,    -3,   -65,     6,   -41,    12,   -35,   -17,    -1,    14,   -18,   -34,   -10,   -23,    31,    10,     7,    15,   -25,     3,    13,   -22,   -91,  -106,   -33,  -136,   -80,   -46,    23,     2,   -77,    57,   -36,   -33,    -7,    -1,   -58,   -28,   -34,   -46,   -71,    -9,   -30,   -18,    25,    15,   -59,    11,     4,   -46,   -31,   -35,   -46,  -106,   -68,   -30,     7,   -16,   -66,    27,    -7,   -35,   -49,   -19,   -61,   -24,     1,   -17,   -11,   -34,    -2,   -35,    19,   -20,   -13,     7,    -7,   -41,    -1,    36,   -21,   -70,   -52,   -20,     4,   -21,  -126,    10,   -46,    13,    -4,   -81,   -22,   -39,   -23,   -26,   -52,   -36,   -26,   -37,     8,     7,   -25,     9,   -34,   -51,     2,    70,    63,    30,   -38,     2,     8,    -6,  -106,    14,   -17,    21,    18,   -19,   -28,   -54,    14,   -10,   -38,   -26,    -5,   -21,    41,    35,    -9,   -36,   -57,    -8,    16,    51,    45,    -7,  -103,     4,     4,     0,   -82,    30,   -29,    -4,   -23,   -34,    -2,   -26,     0,   -45,    16,   -22,    39,     7,    48,    44,     5,   -37,   -19,     9,    62,    63,    49,   -74,   -74,    -4,     0,     5,   -11,    16,   -28,     5,     9,    60,    26,     2,   -23,    -7,     5,    22,    51,    42,    32,    23,    18,    -2,   -17,    -7,    24,    50,    76,   -34,   -51,     5,   -10,    -1,   -38,   -54,   -19,    25,    70,    88,    55,    38,    14,    30,    12,    23,   -46,   -28,   -35,    21,    87,    42,    45,     8,   -35,    10,    15,   -35,    -4,    -4,    -4,     1,    39,   -46,    -8,    35,    60,    79,    54,    50,     1,    20,   -13,   -35,    27,   -14,    -7,    57,    46,    22,    40,   -19,    -7,   -29,     1,     3,   -14,     5,    -3,    -8,     1,    35,     2,    21,    41,    72,   -17,    19,    -2,   -28,    23,   -19,    53,    50,    22,     2,    25,    -9,    73,    17,   -23,    45,    19,    -2,     8,    -1,     6,     4,    -5,     7,    -2,   -35,    15,    10,    14,    -1,    19,    28,    35,    20,    27,     9,    27,   -42,     1,    15,   -24,   -58,   -42,   -38,     5,    -4,    10,    -8),
		    70 => (    2,    -6,    -4,     3,     9,    -4,    -6,     2,    -3,     9,     0,    -5,     0,     0,    -7,    -6,     6,   -10,     2,     3,    -7,     8,     0,    -4,    10,    -2,    -3,    -1,     7,     9,    10,     0,     1,     1,     0,    -2,     6,    -9,    -6,    -1,     7,    19,   -12,     4,    -7,     5,     6,     1,     1,    -2,     8,     9,     0,     2,     3,     3,    -2,     0,     4,    -6,    -6,    -8,   -11,     5,   -15,   -16,    -1,   -17,   -23,   -39,   -16,     9,   -19,   -28,   -13,    -9,     0,   -10,    -3,   -11,    -5,     5,   -10,    -3,    -9,    10,    -9,    -9,    -5,    13,   -19,   -21,   -21,   -78,   -42,   -27,     5,    28,    15,   -42,    -9,    -7,     1,     5,   -18,   -43,   -42,   -20,     8,     4,    -3,    -8,     6,     8,    10,     4,   -16,   -69,   -21,    -4,   -25,    -9,   -15,    42,    56,    63,    30,    17,   -53,   -64,   -17,    10,   -50,   -57,   -29,   -18,   -18,   -33,   -18,     0,    -6,    -4,   -20,    -7,   -13,   -45,   -15,     3,     6,    -1,     7,    20,    68,    18,    18,    32,   -13,   -59,   -45,    30,   -31,   -60,     4,    12,    -3,   -47,   -39,   -25,     9,   -11,    -6,   -14,    13,    18,    24,    23,    27,     8,     1,    58,     8,    -9,     7,     1,    39,    25,   -30,     0,   -22,   -13,    -7,   -13,   -10,   -71,   -36,   -15,     0,    -7,   -16,   -38,     7,    25,    37,    30,    10,    25,     5,    30,    -5,     8,    46,    26,    53,    16,    14,    21,    28,    19,   -37,   -14,   -15,   -15,   -39,   -30,     9,    -8,    36,   -31,    28,     2,    21,   -24,    -4,    38,    30,   -10,   -24,    38,    29,   -10,   -28,   -30,    37,     2,    13,    36,    -8,     2,   -31,   -23,   -59,   -24,     8,    -2,    50,    -7,   -10,   -22,   -41,   -37,    28,    33,    41,    -6,   -14,    37,    -5,     5,   -20,    -6,   -17,    45,    -8,   -21,   -15,   -22,   -41,   -40,   -48,     8,    -2,     8,    48,    11,   -28,    -7,   -32,   -38,    24,    22,    -5,    -1,     2,   -42,   -12,    26,     4,   -23,   -39,   -33,   -44,   -25,   -23,    25,   -10,   -18,   -37,     3,     4,    51,     2,   -25,   -34,    -8,   -17,   -24,    -6,   -10,    21,   -25,   -76,  -113,   -85,   -13,   -27,   -39,   -39,   -42,   -17,   -23,   -16,   -16,    20,   -23,   -17,   -22,     4,     0,    -7,   -15,   -36,   -45,   -20,   -43,   -21,    -8,   -31,    -3,   -92,  -111,  -131,   -60,    31,   -21,   -29,   -12,     8,     6,    -7,   -21,   -48,   -35,   -34,   -24,    -2,     9,    13,    31,   -15,    -1,     7,   -26,   -20,    12,    14,     2,   -68,  -112,   -50,   -25,     1,    19,   -13,   -23,    15,    31,   -12,   -14,   -41,   -31,   -48,   -12,     1,     4,    -9,    29,    18,    -4,   -23,   -20,   -36,    26,    57,    -2,   -65,   -49,   -38,   -46,   -56,    -8,    12,    -3,     7,    28,     9,   -15,   -27,    -4,   -44,   -10,    -1,     1,   -13,    17,    29,     9,   -61,   -22,     9,    45,    74,     2,   -32,   -58,   -18,   -45,   -95,    -7,    -6,   -11,    36,    20,    36,   -26,   -34,    33,   -35,   -38,    -5,     2,    -7,    19,    20,   -32,   -46,   -25,    -7,    17,    35,    34,   -44,   -26,   -35,   -25,  -119,    -6,   -18,   -15,    29,   -16,    23,   -23,   -51,   -21,   -82,   -20,    -1,   -10,   -24,    12,    10,   -24,   -41,   -12,    -4,    19,    35,    11,   -12,   -61,   -84,  -152,   -64,    -4,   -36,   -13,    16,   -22,     2,     4,   -19,   -30,   -61,     2,     3,    -4,   -20,    -4,    -7,   -37,   -45,   -33,   -28,    19,    41,    11,   -21,   -53,  -113,  -121,   -81,   -44,    44,    -1,    30,   -17,    -5,    -1,   -27,   -30,   -41,   -14,    -8,    11,   -19,   -10,   -10,   -16,   -49,   -31,   -16,    52,    20,   -15,     9,   -26,   -52,   -38,   -19,   -13,     2,    -5,    20,    -5,   -29,     8,     6,   -77,   -17,     0,     7,     8,    -5,   -22,    18,    36,   -56,   -32,   -29,     3,    22,    45,   -36,   -13,    43,     2,   -18,   -11,     8,   -25,     4,    15,   -32,    22,     7,   -59,    23,     9,    -4,     7,    -2,    -9,   -12,    -3,   -73,   -15,   -36,   -22,     6,    28,    39,    38,    27,    34,   -34,   -25,   -13,     7,    29,     5,     4,    14,    14,    -8,    20,    27,     1,     0,    -3,   -13,   -23,   -11,   -31,   -15,   -17,    -1,   -22,    30,    -5,    22,    29,    -7,    15,   -16,     3,    23,    33,    16,     9,    19,    -9,     4,    20,    17,    -1,     4,    -7,   -28,     3,   -11,   -47,   -65,   -22,    25,    -8,   -19,   -10,    36,    24,    48,    67,    67,    17,   -36,   -31,   -14,    -8,   -26,     9,   -38,   -16,     2,    -2,    -7,   -15,     4,    25,   -14,   -33,   -28,   -46,   -20,   -17,   -24,   -18,   -15,   -24,    -1,    -5,    10,    -6,   -32,   -15,     3,     2,   -17,   -13,    -5,     4,     0,     6,     9,     8,    -5,   -11,    -2,   -20,    -4,   -10,    -6,    -7,   -14,   -12,   -17,    -4,   -73,   -53,   -58,   -31,   -40,   -48,   -32,   -29,    -6,   -10,     8,     3,    -3,     2,    -8,     7,    -2,     0,   -27,   -41,    -4,    -9,    -2,   -18,   -14,   -10,   -36,   -47,   -39,   -35,   -58,   -61,   -12,   -53,   -38,    -8,    -6,   -10,    -9,    -1,     8,     1,    10,    -9,    -3,     9,     6,    -5,     4,    -9,    -9,   -10,   -11,     3,   -20,   -11,    -6,    -8,    -7,    -9,    -1,    -6,   -19,   -15,   -10,    -5,     3,    -3,    -4),
		    71 => (   -5,   -10,    -9,    -6,    -4,    -3,     3,     1,     3,   -10,    -4,     5,     4,    -6,     7,     5,     5,     4,     9,     2,    -9,     1,    -5,   -10,    -6,     8,    -9,     8,    -6,    -5,     3,     6,     4,     4,     6,     6,   -10,     4,    -5,     5,    -6,    -4,    27,     9,    19,     0,   -12,    -8,    -8,     6,    -6,    -9,    -2,     5,    -8,     4,    -6,     8,    -5,    -4,    -7,     6,     5,     7,   -31,   -35,   -20,   -17,   -45,   -24,   -34,    -1,    45,    -4,   -13,   -11,   -30,   -74,   -50,   -35,   -13,   -17,     1,    -6,     6,    -7,    53,     4,     2,   -16,   -17,    -6,   -33,   -48,   -54,   -67,    -5,     7,   -66,   -19,    32,    36,    37,    33,    37,    41,   -16,    -3,   -12,    -4,    -3,     9,     4,    -6,    43,    44,    12,    18,     5,    -5,    17,    -1,    15,    -6,    -3,    20,   -36,   -50,    -6,    13,    25,    41,   -23,    33,   -18,     7,    -9,   -32,   -44,   -18,     9,     5,    24,     8,    12,    20,    -3,    -9,   -32,   -22,   -22,     3,    36,     2,    29,    32,    13,   -45,    -4,    25,    19,    18,    14,     9,   -11,   -35,    -8,   -20,    -4,    -1,   -30,   -28,   -10,    15,     7,    -7,   -86,  -126,   -55,     5,   -12,   -24,   -17,   -10,     4,   -50,    32,    -8,     7,    31,    20,     8,    -4,     2,   -22,   -12,     5,    -7,   -37,   -34,   -42,    17,    18,   -41,   -80,   -38,     0,   -30,   -10,   -35,    -8,   -41,   -27,   -21,    20,    10,    23,    49,    16,   -11,   -19,     3,   -41,    -9,    -4,   -14,   -51,   -37,   -53,   -16,    56,    10,   -64,   -29,     6,   -12,    39,    37,     4,   -14,   -25,   -33,   -46,   -59,     3,    25,    34,   -20,   -32,    -5,   -43,    -2,    -3,    -1,   -28,   -43,   -33,    -4,     8,    34,    22,     6,   -41,   -21,   -19,    22,     7,    -4,   -35,   -32,   -57,   -80,   -32,   -11,    14,    36,   -15,    50,    39,   -17,    -5,   -15,   -32,   -19,   -24,   -26,   -41,   -24,    29,   -19,   -49,   -16,     8,    41,    10,   -38,   -13,     4,   -41,   -21,   -54,   -66,    29,    33,   -23,    40,    34,    35,    -2,    -2,   -12,   -11,   -23,   -26,   -40,   -39,   -54,   -64,   -53,    -3,    11,     1,   -17,   -41,   -34,     3,   -47,   -39,   -22,   -29,    25,    33,   -20,    37,    22,    59,     9,     8,   -14,   -20,     2,    -7,    -1,    -1,   -41,   -21,    -9,     7,    35,    33,    -9,   -15,     6,    46,   -56,   -53,   -19,   -19,   -24,   -11,    -1,    51,    62,    74,    -6,     4,    -4,     1,    -4,    22,    16,     8,    35,    38,   -17,   -14,   -12,   -55,    -3,   -10,     9,    10,   -74,   -71,   -46,   -41,   -45,   -69,   -44,    66,    52,    -5,     9,    -6,     3,    13,   -13,    23,    25,   -12,    75,    66,    24,   -42,   -62,   -50,     8,    -9,    36,    -4,   -34,   -59,   -23,   -36,   -30,   -13,    -6,    -5,     5,     1,    -2,    -6,     3,   -16,   -25,   -19,   -39,    20,    30,    68,     2,   -23,   -18,    -6,    -8,    -5,    22,    -7,   -15,   -44,   -44,   -52,   -38,   -37,   -48,    -4,    -3,   -18,     3,     4,     3,   -24,    -3,    17,   -37,    -2,    29,    16,    12,   -40,    -5,   -10,     9,   -49,     0,   -20,   -40,   -79,   -52,   -78,   -49,   -40,    -3,   -51,   -28,    -9,     9,    -3,    -3,   -25,    -1,    17,   -20,   -51,   -15,   -37,   -49,   -89,    12,    36,    10,    -6,     2,   -38,   -76,   -62,   -28,   -50,   -38,   -20,   -13,   -28,   -34,   -53,    19,    -4,   -15,    -6,   -43,   -36,   -56,   -68,   -71,  -115,   -89,   -98,   -42,   -10,    41,     7,     5,   -22,   -67,   -35,   -31,   -27,   -27,   -29,   -42,   -20,   -35,   -14,     2,    -6,     7,   -28,   -32,   -84,   -32,   -58,   -23,   -62,   -71,   -97,   -64,   -46,    45,    35,     4,    -8,   -37,   -15,   -39,   -28,    -3,     7,   -17,   -15,   -23,    -2,    -5,     3,   -13,    15,    27,   -13,    14,   -20,   -28,    23,    22,     1,    10,   -52,    49,    36,    35,    23,    66,     9,    34,   -34,   -41,    -6,    15,   -24,   -17,    -4,    16,     0,   -23,    34,    48,    27,    43,    37,    -4,   -21,     7,   -16,   -42,   -34,    20,    23,    49,     3,    51,    17,    46,    13,   -65,   -37,   -19,    -8,   -35,     0,    17,    15,   -67,   -34,    62,    84,    51,    27,     8,   -29,   -47,   -26,     1,   -22,   -13,    80,    32,   -23,    12,     5,    20,     8,   -34,   -38,   -26,    -6,     2,    -2,     8,    10,   -14,   -29,    10,     3,    32,   -40,   -58,   -24,   -65,   -50,     9,    -5,     1,    17,     7,     2,     8,   -12,     6,   -26,    -1,   -15,   -19,   -42,    54,    -4,     5,     4,     0,   -16,     3,    -4,   -14,   -14,   -37,    38,    34,     7,   -17,   -67,   -60,    15,   -12,    23,   -40,  -103,   -48,   -36,   -54,   -37,   -50,    64,    70,     9,    -6,     3,    -8,   -11,    -2,    -8,   -21,   -10,   -12,   -23,   -30,   -55,   -43,   -89,   -41,   -66,   -50,   -99,   -68,   -49,   -73,   -21,   -14,   -17,     0,    -9,   -16,     1,     0,    -1,    -2,    -6,    -8,   -14,    -5,   -19,    -5,   -21,    -2,     0,   -68,   -50,    23,    14,    41,   -67,   -21,   -17,    -1,   -15,    -2,     3,     9,     0,     9,    10,    -6,    -2,    -1,    -1,     9,     9,    -6,    -1,    -9,    10,   -21,   -17,   -10,   -13,   -25,   -23,   -17,    -2,     8,     7,    -9,     7,    -3,     2,     3,     1,    -7,     6),
		    72 => (   -7,    -3,    -1,   -10,    -3,     9,    -5,     4,     5,    -1,     6,     6,   -22,   -21,    14,     8,     7,    10,    -9,     7,    -2,     8,    -1,     6,    -6,     4,    -4,    -2,    -5,     0,     1,     2,     2,     5,   -11,     1,   -44,   -27,   -43,   -55,   -39,   -54,   -26,   -37,   -13,   -26,   -37,   -80,   -56,   -18,   -14,   -17,     9,     2,     3,     6,    -6,     0,   -13,   -11,   -34,    -4,    -5,   -52,   -19,    46,    41,    -5,   -12,   -81,   -66,  -107,   -73,   -19,     2,   -16,   -91,   -25,   -32,   -13,    21,     8,    -6,     9,     0,     4,   -14,   -39,   -19,     9,     4,    -1,    18,    17,    30,    -1,   -44,   -99,   -75,   -85,   -83,   -68,   -75,   -66,   -75,   -55,   -35,   -15,     3,     3,     9,     4,     5,    -9,   -28,    -4,     5,   -20,    25,    23,     7,   -14,    33,     6,   -30,   -87,   -76,   -63,   -72,   -44,   -70,   -69,   -45,   -52,   -35,   -30,     3,    -7,   -33,   -13,    -9,     7,   -19,    -1,    21,   -30,    44,    41,    46,     4,    26,   -25,    20,    -1,   -34,    -6,   -87,   -88,   -63,   -39,   -23,   -44,   -57,   -19,   -34,   -11,    -6,   -17,    -9,     3,    -6,     7,    19,    50,    33,     9,    29,    35,     0,   -10,    -8,    24,    -8,   -38,   -44,   -46,   -46,   -22,   -19,   -44,   -43,   -35,   -55,   -19,   -16,   -15,    -1,    -4,    -3,   -19,    -8,    -7,   -35,   -19,     4,    11,   -42,    -5,   -12,   -11,   -29,   -32,   -42,   -11,   -46,   -54,   -49,   -66,   -72,   -79,   -56,   -35,   -32,   -20,   -32,    59,   -13,     1,   -55,   -16,    14,   -15,     4,   -20,    21,   -19,   -24,    28,    29,     6,   -17,   -16,   -36,   -42,   -83,   -86,   -70,   -68,   -77,   -32,   -44,   -21,    -8,   -28,   -17,    19,   -64,   -10,     3,   -22,    -1,    -4,    14,     5,    12,     6,    82,    24,   -12,   -36,   -48,   -40,   -53,   -50,  -104,   -26,    67,   -58,   -19,   -25,     0,   -21,   -17,    -8,   -77,    27,    -4,    -2,    -1,   -30,   -35,   -17,    10,   -13,    19,    51,    40,   -30,   -46,   -28,   -30,   -52,   -53,    11,    40,   -29,   -43,   -38,    -1,    -6,   -56,   -23,   -29,   -22,   -23,   -15,   -24,     1,    13,    56,   -31,   -50,   -10,    16,     5,   -13,    -8,   -42,   -50,   -72,   -41,     5,    -9,   -42,   -77,    -8,    -7,   -10,   -67,    -9,    -6,    18,   -43,   -76,    -9,   -26,   -40,   -25,    -5,    -3,   -21,    -9,    22,   -11,    -6,   -52,   -41,   -14,    10,   -66,   -18,   -23,   -35,     7,    -7,   -10,   -51,    -2,   -11,   -16,   -60,   -80,   -19,   -31,   -57,   -33,   -20,     3,   -25,    20,     5,     9,   -25,   -30,    16,    48,    62,    11,   -17,   -11,    41,    39,     5,    -4,   -11,   -16,   -44,    -5,   -69,   -49,   -20,   -45,   -15,   -21,    -1,    15,    10,    16,    23,    -3,   -28,     0,    20,    50,    29,    -7,   -16,     2,    81,    40,    -2,   -14,    43,   -34,   -10,    -6,   -11,   -39,   -24,    -8,    11,     1,    36,    55,    20,    25,    -1,   -12,   -11,     3,    27,     6,   -27,   -41,    -1,    14,    22,    49,     5,     2,    47,   -10,    27,   -35,     5,   -11,   -65,   -15,    13,    36,     5,    28,    23,    21,    44,    24,     5,    21,    -4,    20,    18,    22,    15,    28,   -11,    47,   -10,    -3,    69,    10,    37,   -19,    35,     4,   -17,     7,    25,    31,    -5,     6,    35,    32,    37,    26,    36,    53,    32,    40,   -15,    10,    -2,   -20,   -52,    44,    -5,     5,    30,    24,    20,    16,    54,    -6,   -29,     9,    29,    31,   -22,    12,   -16,    25,    14,     6,    31,    19,     9,    32,    26,    38,    62,    32,   -38,    30,     1,   -36,     5,    55,    -8,    34,    23,    14,    -4,    40,    11,    -9,   -31,   -24,   -11,    29,    -3,    -3,   -18,   -26,   -27,     0,    36,    61,    36,    19,    34,    71,    -4,   -17,    11,    40,     5,   -11,     8,   -18,    20,    -7,     1,    -6,    -8,     4,    10,    -2,   -49,   -72,   -62,   -59,   -53,   -14,   -27,   -14,   -16,   -50,    28,    -5,     9,    -3,    -8,    23,    17,    12,    61,     1,    -3,    -7,    36,   -31,    12,   -22,   -29,   -30,   -94,  -141,   -19,   -28,   -47,   -56,   -61,   -83,   -83,   -41,   -37,    -1,    10,     6,    -3,    -4,    -3,    21,    12,   -27,   -29,   -31,   -42,   -17,   -20,   -39,   -33,   -87,  -135,  -125,   -38,   -22,   -50,   -75,   -92,   -68,   -67,   -56,   -90,    -1,     6,   -10,     8,    -9,   -12,   -19,   -24,   -41,    -2,    -3,   -59,   -64,  -115,   -99,  -131,  -106,  -124,  -119,   -82,   -87,   -81,   -87,   -76,  -106,   -83,   -47,   -84,     8,    -1,     8,   -26,    -8,   -94,   -26,   -59,   -17,     7,   -43,     6,   -27,  -179,  -128,  -112,   -93,  -106,  -117,  -100,   -96,   -91,   -97,   -74,   -75,    13,    32,    29,     1,    -4,     1,    -3,     5,   -25,   -17,    -4,   -14,   -71,   -95,  -103,   -64,  -101,   -94,   -66,   -81,   -82,   -62,   -48,   -81,   -84,   -70,   -19,   -20,    -1,    17,    20,     4,    -2,    -7,    -9,     5,     0,   -31,   -51,   -49,   -72,   -90,   -66,   -23,   -28,   -32,   -47,   -18,   -38,   -33,   -17,   -58,   -30,   -20,   -37,    -8,    -8,     1,     2,    -5,    -6,     2,     4,    -7,    -1,    -6,   -10,    -3,     7,   -13,   -23,    -5,   -13,   -34,   -20,    -4,   -18,   -16,   -29,   -16,   -22,   -23,   -21,    -8,    10,     9,    -2,     0),
		    73 => (    8,     1,    -8,     5,    -9,     6,    -3,    -7,    -7,     1,     4,     9,   -12,    -6,   -15,     1,    -3,     7,    -7,   -10,     6,     4,     1,     3,     5,    -9,    -3,     1,    -5,     6,     6,    -3,     1,    -1,    -6,     2,     1,     1,   -11,   -10,    -7,   -14,   -26,   -21,   -14,   -11,    -3,     5,     1,     3,     5,     0,    -6,    -4,     9,    -1,    -6,    -2,    -6,    -2,    -3,     5,     3,   -11,   -16,   -28,   -79,   -78,   -78,   -15,   -16,    -2,   -11,   -11,     6,     0,   -24,    -5,     0,   -17,    -9,    -2,    -3,     0,    -6,     0,    -2,    -1,     0,   -16,   -10,    -2,    12,     2,   -12,   -45,   -27,   -41,   -56,   -62,   -58,   -24,   -19,   -10,   -16,   -21,   -31,   -41,     1,    -1,    -9,     2,    -5,    -2,     8,     5,     0,    -6,   -17,   -57,   -43,  -103,    13,    36,    -8,    -8,    33,     8,     0,    -7,    -4,    -1,   -10,    32,    64,   -42,   -44,   -37,    -5,     1,    -3,     0,     6,    -7,     2,   -34,   -24,   -34,   -77,   -81,   -30,    35,    28,   -37,   -17,   -20,     1,   -26,   -20,   -31,     4,   -38,   -14,   -29,   -26,   -93,   -29,    -8,     0,     4,    20,    14,    -1,   -28,    10,   -17,   -11,    22,    52,    13,    -7,    18,   -12,    13,    18,   -38,   -17,   -46,     4,     0,   -29,    -5,   -22,   -44,   -65,   -20,     9,     9,     6,    -4,     8,   -91,   -73,   -33,     9,     5,    -2,   -41,    12,    64,     4,   -27,   -33,   -11,     1,   -13,   -15,   -29,   -18,   -46,   -68,   -41,   -51,    -7,    -1,    -5,    -7,   -16,     0,   -65,   -45,     5,     9,     9,   -19,   -14,    32,    27,    -7,   -18,     6,   -19,   -14,    -6,    -9,   -11,    -1,   -26,  -119,   -36,   -80,     9,   -10,   -13,     7,   -17,   -38,   -36,   -15,    22,    -7,    10,    23,    48,    31,   -12,   -11,   -27,    15,    27,   -19,     5,    10,    -9,    15,     9,   -96,   -35,   -46,   -40,     3,   -23,    -5,   -11,   -20,   -38,   -14,   -37,    18,     4,    16,    50,    29,   -46,   -55,   -21,   -26,   -18,   -32,    12,    42,   -33,    11,    -4,   -91,   -77,   -70,   -31,    -8,   -30,     0,    20,    46,    30,    13,     0,    44,     7,   -46,   -52,  -177,   -68,   -28,   -35,   -26,    -9,   -25,     9,    27,    51,    -5,    24,   -75,   -51,   -33,     7,    -3,   -19,    80,    15,    56,    36,     3,   -63,   -53,   -86,   -87,  -120,   -90,   -11,     3,   -18,   -17,   -35,   -22,    -7,    15,    37,    31,    27,   -49,    12,   -25,     0,    -5,   -31,   -38,   -49,   -54,   -45,   -37,  -136,  -120,   -92,   -50,   -30,     7,    49,    47,   -30,     4,    -7,   -15,     3,    -8,   -15,   -17,    -8,   -55,   -36,   -45,   -15,     0,    11,    25,   -21,   -38,  -105,  -102,  -119,   -14,    34,    18,   -19,    -1,    26,    -3,    12,    -9,    24,     2,   -37,   -47,   -25,   -26,     5,   -31,   -73,   -45,   -14,    -9,     3,     1,   -10,   -53,  -112,  -145,    51,    48,     8,    12,    21,    42,    40,    36,    10,    -7,    -6,     7,   -10,   -57,   -36,   -68,   -29,   -31,   -42,    44,   -12,    -6,     8,    22,   -17,   -22,   -39,   -15,   -18,    26,    37,    38,    42,    35,    28,    33,    -9,    -3,   -23,    -7,   -28,   -66,   -45,   -42,     6,   -20,   -27,   -13,   -14,     8,     8,    19,    15,   -49,   -51,   -24,   -36,   -13,    16,    57,    21,    58,    52,    12,   -53,   -37,     2,   -13,    -4,   -66,   -47,   -34,   -24,   -74,   -28,    -9,    -6,   -18,   -12,     5,    19,   -46,   -87,   -95,   -30,   -46,    -3,    21,    39,    52,     8,     2,   -22,   -24,   -43,    18,    -6,     9,   -24,   -25,   -64,   -76,   -13,    -8,    -7,    -9,   -25,     4,    -5,   -73,   -67,   -80,   -72,   -96,   -69,   -86,   -33,   -63,   -23,   -44,   -23,    31,    20,    40,     6,   -34,    14,   -34,   -68,   -75,    -4,   -36,   -11,     5,   -24,    14,    51,   -19,    -6,   -75,  -122,  -129,  -193,  -256,  -189,  -150,   -53,    -7,   -24,    -7,    34,    47,    28,    11,   -18,   -34,   -89,   -71,   -46,   -12,     9,   -13,    -8,    38,    82,    50,     0,    -7,   -49,   -10,   -39,   -40,   -60,   -41,   -31,     2,    18,    -3,    -2,    25,     0,    24,    -9,   -24,   -61,   -45,   -17,   -23,     9,    -7,     3,    10,    45,    84,    79,    57,    36,    32,    19,    44,    18,   -17,    10,    11,    11,    21,    -7,   -13,    -4,   -24,   -17,   -44,   -28,   -47,   -28,    -4,     0,     6,     8,     9,   -20,    57,    56,    50,    43,     9,   -14,    22,    -2,    32,    56,    -2,    28,   -58,    10,    -5,   -39,    27,     8,   -15,   -14,   -51,   -31,    -6,     9,    -6,    -5,    12,    36,    73,   -13,    38,    31,     4,     6,    28,    33,    21,    25,    -5,   -11,   -22,    15,  -103,   -29,    21,    26,    37,    39,   -63,   -18,   -25,     1,     7,    -4,    11,   -40,     1,   108,    70,    59,    25,    34,     5,   -15,     7,   -15,   -39,   -17,   -15,   -39,  -105,   -22,   -30,   -66,   -25,   -80,   -49,   -26,   -35,     9,     4,     8,     0,   -32,   -63,    -1,     6,   -13,   -13,   -52,     0,     6,   -19,     8,     0,   -53,    -7,    24,    18,   -26,   -13,   -22,     8,    -7,    -8,    -3,     5,    -1,     9,    -7,    -9,    -1,    -6,   -23,    -8,    -6,    -7,   -59,   -53,   -41,   -28,   -35,   -37,   -38,     3,    -6,   -19,   -42,   -38,    -8,   -32,     2,    -8,    -4,    -1,    -3),
		    74 => (   -3,    -1,   -10,     1,     2,     8,    -3,     5,     9,     6,     6,     9,    -7,   -31,    -6,    -2,    -8,    -2,   -10,    10,    -6,    -7,    -3,     4,    -3,    10,    -6,    -2,     0,    -2,    10,    -7,     9,     8,   -38,   -37,   -14,   -33,   -60,   -34,   -72,   -44,    18,  -110,   -98,   -70,   -20,    -4,   -46,    -8,     0,   -16,    -9,     4,     5,    -7,    -2,    -6,   -16,   -42,   -62,   -42,   -21,   -57,   -35,   -36,   -96,  -124,   -95,   -22,    13,   -31,   -55,   -45,   -63,   -83,   -85,   -54,   -56,   -68,   -17,   -41,     7,   -10,    -8,    -2,   -26,   -78,  -127,   -43,   -49,    -5,   -87,   -99,   -60,   -84,  -143,   -48,    15,   -10,   -37,   -56,   -76,   -25,   -19,   -40,   -24,   -71,   -83,   -34,    -3,     4,     0,     0,   -14,  -110,   -12,     4,     6,    17,    -5,   -58,   -42,   -40,   -11,    29,    35,    16,     9,    25,    41,     1,   -22,     8,    83,     3,    -9,   -17,   -75,   -22,    -6,     5,   -27,   -51,     9,    24,    16,    67,    37,    28,    27,   -12,    25,    41,    64,    16,    -4,    47,    16,    56,   -11,    37,    36,    62,    63,    35,   -71,     0,    -7,     4,   -24,   -14,    42,    29,    11,    70,    57,    62,    37,    22,    12,    64,    80,   104,    62,    14,   -29,     0,    26,     3,    -6,    61,    80,    23,    16,   -42,    -1,   -41,   -35,    20,    45,    21,    43,    72,    32,   149,    95,   132,    72,    80,    73,    67,    40,    46,    16,    52,    22,   -22,   -16,     7,    32,   -32,    84,   -58,   -42,   -48,    52,    24,    24,     4,    56,    30,    -4,   125,    72,    81,    13,   -16,    -7,    20,   -24,   -25,   -24,    -9,    11,     8,   -56,   -20,    -1,    21,    39,   -64,     4,   -19,    41,   -34,     6,   -30,   -43,   -20,   -20,    -2,    22,   -53,   -20,     9,   -16,     9,   -39,    20,    -9,   -14,   -12,   -15,   -68,     0,   -14,   -39,   -38,   -34,     7,   -25,    23,   -22,   -21,   -47,   -82,   -36,   -38,    11,   -22,   -63,     0,   -51,   -43,   -22,   -21,    -3,   -52,    -1,   -65,   -34,   -16,   -41,   -88,   -25,    -6,   -51,    10,   -43,    22,   -34,   -42,   -35,    29,   -61,     8,   -26,   -55,   -17,    -7,   -18,   -31,   -11,     7,    34,   -45,   -39,  -107,   -44,   -29,   -65,  -106,   -26,   -43,   -83,    -7,    10,     8,   -34,   -58,   -17,    -7,   -41,    -8,     6,   -31,    18,    62,    31,   -59,     1,    12,    25,   -14,   -27,    -1,    32,   -15,   -42,     8,    50,   -40,   -68,    -3,   -20,   -57,   -53,   -58,    -6,     5,    58,    33,   -26,    18,    57,    72,    -7,    20,    10,    -1,    29,    34,    -9,     3,   -31,   -38,   -17,     6,    28,   -20,    -8,    -9,    32,  -100,   -69,    -1,    -2,    -2,    93,    53,    30,    52,    38,    24,   -16,   -21,    -8,    13,    12,   -17,    -8,   -42,   -53,   -12,    -9,    -3,    40,   -55,    -7,   -10,     9,    43,    10,    51,    -3,    34,    44,    53,    26,     9,    10,    47,    32,    10,    -5,    23,    48,   -13,   -23,     3,     4,    46,    27,   -19,    -5,   -36,   -56,     6,     2,   -62,    14,   -26,   -26,   -23,   -20,     2,    -3,    28,    28,     3,    -1,    11,    -7,    16,    20,    10,    22,    48,    33,    34,    -8,    22,     9,   -33,   -23,     2,    -5,   -40,   -52,     1,     4,   -28,    47,     8,   -10,   -54,   -22,     5,   -37,   -10,   -37,    40,    -9,   -17,    12,     2,    36,    14,    67,    20,   -79,   -14,   -26,   -42,    -9,   -15,     2,     7,    38,    20,     6,   -44,   -18,   -53,   -37,    20,   -24,     5,   -24,   -30,   -63,   -19,    50,    84,    51,    31,    57,    37,   -21,   -36,   -51,     3,   -38,   -56,   111,   -29,   -19,   -31,   -55,   -22,   -49,   -59,   -60,    -6,     4,    19,    27,    11,   -65,    -1,    25,    28,    21,    36,     6,    12,    -5,   -15,   -41,     7,   -12,   -29,    27,   -36,   -54,   -60,   -65,   -35,    26,     4,     6,     1,   -10,     3,    22,    35,    -9,    41,    38,    59,    38,    15,   -12,   -59,   -68,   -29,    -8,   -16,    -5,   -42,    35,    26,   -24,   -39,   -32,    10,    15,     0,    18,   -43,   -21,   -13,    26,    30,    24,    -8,    51,   111,    85,    88,    27,   -21,   -95,   -63,     3,   -16,   -15,   -18,   -54,  -116,   -62,    -1,    20,    48,   -20,    59,     7,   -12,    -2,   -44,   -26,    45,    42,    -2,    84,    97,   106,    67,    55,     4,    -2,   -18,   -12,    10,     6,    -3,   -77,   -99,  -184,    32,    51,    78,    50,    89,    67,    28,     2,   -15,   -26,    16,    -7,    40,    91,    90,    39,   -37,    40,    -1,    57,   -18,    -2,     2,     6,     4,   -29,   -96,   -16,    77,    83,    23,    60,     9,    70,   -22,    -3,    -4,   -63,   -30,   -35,    47,    82,    -1,   -27,   -14,    -6,   -50,    48,   -47,    -4,     1,    -2,   -30,    -3,    81,   112,    37,   -30,   -22,    10,    42,    37,   -40,    22,   -52,    17,     7,   -12,   -13,   -10,   -13,   -20,   -18,    10,   -20,   -53,   -39,     9,     3,    -9,     1,   -72,   124,   105,    61,   -21,   -44,   -71,  -123,   -25,   -36,   -40,   -23,   -91,   -95,   -63,   -16,    -6,   -73,  -147,  -129,   -34,     7,    -8,    10,     6,     0,   -10,     5,    -4,   -15,    -3,   -43,   -47,   -31,   -38,   -51,   -61,   -50,   -17,   -37,   -15,   -78,  -116,   -92,   -55,   -59,   -27,   -42,     4,    10,     1,     0,     1),
		    75 => (   -7,     8,    -8,    -2,     0,    -3,    -7,     5,    -4,    -8,     1,    -2,     7,     3,     2,    -8,    10,     1,     6,    -1,     7,     4,    -2,    -3,     8,     4,    -7,    -6,    -6,     0,    -8,    -2,    -9,     8,    -1,    -2,     8,     6,    -9,   -11,   -17,   -30,   -22,   -15,   -13,   -30,   -21,    -2,    -4,   -13,     4,     5,   -10,    10,    -5,     3,     3,    -3,    -8,    -8,     2,     2,   -23,   -15,   -49,   -50,   -59,   -60,   -31,   -38,   -93,   -15,    11,    11,    -8,    30,    51,     3,     0,    14,   -25,    -5,     9,     0,     3,     2,   -10,    14,    27,   -40,   -47,   -50,   -30,   -16,   -17,   -26,     6,    15,    29,    34,    28,    -4,   -34,   -26,    10,    30,     9,    26,    13,     8,    13,    10,     6,    -6,     0,    22,     0,    -4,    26,    39,    11,    39,     2,   -49,   -29,    -4,    17,    40,    45,     5,    -3,   -31,    -9,     3,    22,    28,    21,    31,   -19,   -28,   -10,    -4,     5,     5,   -27,     1,    39,    21,    25,     5,    -9,   -38,   -45,    -9,     2,   -11,    -3,    -2,    -6,    49,    36,    -1,    31,    32,    29,    23,   -22,   -25,     3,    -9,   -42,   -28,    18,    25,    54,    17,     5,    -5,    -1,   -24,   -30,   -13,    -4,    -2,   -10,   -23,    11,    52,    55,    38,    29,    17,    29,    29,    20,    10,    -8,     4,     4,   -35,     8,    63,     9,    13,   -24,   -11,   -17,    -9,   -16,   -23,    -5,   -24,    -2,    -9,   -14,     4,    24,   -10,    30,    27,    59,    33,    25,    28,    -8,   -30,   -34,   -55,    11,     2,     3,     6,   -20,     6,     1,    26,    17,    18,    -3,   -34,   -31,   -47,     9,    13,   -16,     3,    46,    60,    29,    43,    26,    15,    -3,   -14,   -70,   -49,     5,    10,     4,     4,   -22,   -14,    22,    32,    47,    36,   -17,   -20,   -41,   -38,   -15,     1,    19,    47,    58,    56,    46,     9,    38,    11,     5,    -4,   -11,   -74,    -2,    -2,    -5,    20,   -21,     7,    -3,    46,    62,     6,    28,     1,   -45,   -16,     4,    28,    54,    81,    76,    59,    55,    28,     3,   -27,     7,   -11,    -7,   -47,    16,    -1,    11,    19,    26,    -9,   -19,    45,    36,     4,    30,   -27,   -39,   -62,    49,    42,    74,    29,    35,    37,    49,    43,     8,   -33,     4,     5,     0,   -56,    16,    26,    28,    28,    49,    33,   -29,     1,    13,     4,     8,   -14,   -41,    -4,    25,    49,    29,     1,   -10,    30,    19,    20,    47,   -35,   -10,    -1,    -7,   -61,     1,    19,    22,    42,    29,    43,    56,    25,    20,   -17,     1,   -40,   -24,   -20,     0,    42,    37,    40,    -1,   -26,   -26,    -2,    37,   -32,     8,     0,   -14,   -81,    -7,    11,    30,    36,    34,    25,    59,     7,    12,     3,    -1,   -32,   -15,    15,    56,    45,    39,    31,    24,   -22,   -38,   -37,   -26,     3,     9,   -11,   -20,    -8,    17,    29,    -3,    13,    31,    49,    56,    -6,    -5,     3,    29,     7,    -2,    22,    33,    47,    26,    24,    14,     1,     8,   -40,   -25,   -52,    -2,   -15,   -37,    -5,    19,    71,    18,    12,    30,    32,    29,   -34,     6,    11,     6,    22,   -25,     7,     2,     7,    40,    72,    33,     2,   -18,   -41,   -30,   -63,    -7,    -4,   -30,    16,    26,    68,    46,    40,    50,    45,   -15,   -19,   -33,     1,    34,   -25,     6,    -8,    -7,    -4,    30,    19,    35,     8,    -9,   -43,   -70,   -73,    -2,     2,   -44,     7,    12,    60,    45,    35,    55,    43,    -4,   -41,   -67,    18,    22,     2,    -4,   -18,   -23,   -32,   -10,     2,    -5,    18,    19,   -30,   -83,   -46,    10,   -10,    33,     4,    14,    30,    32,    62,    42,    -3,   -23,   -24,   -36,    21,     1,     9,   -22,     7,   -11,     6,     7,    -5,    -4,    29,    11,   -32,   -90,   -38,     9,    -6,    22,    19,    16,    12,    33,    42,    53,     1,   -21,   -32,     7,     4,   -21,   -14,   -10,     5,    28,    28,   -13,    14,    17,    34,   -36,    -8,   -62,    -3,     1,     1,     7,     6,    10,    29,    36,    49,    46,    36,     1,    21,    12,     9,    -1,   -11,    -2,    -4,    13,    31,    37,     4,    12,     8,   -40,    -2,   -38,    -9,    -6,    -4,   -44,    -5,    17,     9,    34,    23,    51,    29,    13,    49,    23,     6,     5,     6,   -18,   -23,   -18,     7,    12,   -24,   -16,   -22,   -54,     5,    35,    -7,     1,    -2,    11,     0,   -24,    -4,    22,    38,    25,    14,    -2,    23,    21,    21,    15,   -15,   -58,   -42,   -23,   -22,   -11,   -41,   -25,   -40,   -13,    17,    28,     5,   -10,    -7,   -12,     1,   -32,   -15,    28,    13,    11,    26,    29,    21,    10,   -15,    10,    -1,   -36,   -29,   -12,   -31,   -35,   -28,   -21,   -18,    11,   -65,   -22,     2,     7,    -2,     6,    33,   -59,   -48,    -5,    15,   -22,   -36,    35,    18,    20,    10,     0,    16,    23,    40,    30,    -8,    23,    12,    44,    13,     3,    -2,    -5,     0,    -5,    -8,     0,   -30,   -46,   -62,   -71,   -12,    -3,   -17,   -13,    36,    -8,    11,    33,    19,    21,     6,   -16,    -8,   -32,   -24,     8,   -37,     0,     0,     8,    -5,    -5,    -9,    -8,    -6,   -16,   -13,    -5,    -1,    -7,    -2,     8,     1,   -16,    -9,   -15,    -8,    -3,     6,    -6,   -24,   -14,   -50,   -37,   -14,    -5,     7,     6,    -5),
		    76 => (    5,    -3,     7,    -3,     1,    -5,   -10,     3,     6,     8,    -3,     3,     3,     5,    -5,    -7,     4,     3,     4,    -2,     8,    -5,     3,    -2,    -9,     3,    -6,    -2,    -5,    -8,    -4,    -2,    -4,     8,    12,    18,    30,    16,    11,    19,    18,    11,   -10,   -14,   -24,     6,    -3,    -4,    54,    22,     9,    16,     6,     3,     1,     3,     4,    -4,    12,    10,    45,    16,    -1,    32,    41,     5,   -14,     1,    -2,    10,   -23,   -12,   -14,    16,    -2,    13,    18,    67,    82,    66,    61,    28,    -7,    -4,     4,     1,   -21,   -21,    -4,     1,     3,    -7,    -6,    -5,   -14,    -9,   -61,   -59,   -59,   -31,   -39,   -50,    14,    62,    62,    40,    17,    58,    60,     5,   -48,    -7,     8,     7,   -16,     3,    21,    11,   -19,   -28,   -33,    -5,   -17,   -28,   -54,   -72,   -80,   -62,   -26,   -34,   -25,     6,     8,    49,     5,    56,    18,   -16,    30,    37,   -10,    -5,   -24,   -29,    20,     9,   -12,   -17,   -12,    -6,   -35,   -46,   -50,   -47,   -36,   -16,   -25,   -10,     0,     4,   -15,    16,    32,    50,    58,    51,    65,    38,    -8,    -6,     2,    -7,     9,    12,   -14,    -8,   -30,    -8,   -32,   -31,   -22,   -34,   -62,   -68,   -55,   -13,   -12,    14,     2,   -15,     8,    43,    57,    32,    25,    56,     6,    -5,     3,    -4,    27,    13,   -31,    -6,    -3,    21,   -46,   -47,   -42,   -75,   -51,   -76,   -25,     3,    13,   -21,   -22,     8,   -25,   -23,    16,    32,    22,    61,    -2,    -1,    -3,   -14,    34,     3,   -53,   -24,   -15,    -7,   -61,   -64,   -75,   -71,   -61,   -43,    11,     6,    19,     4,     0,   -15,   -19,   -10,   -55,   -29,    48,   -31,     6,    -9,     1,   -26,    45,    -5,   -48,    -7,    13,    -9,   -55,   -65,   -70,   -71,   -39,    18,    21,    11,    -6,     9,   -12,   -22,   -19,   -39,   -50,   -33,   -25,   -17,    -5,    -9,    -2,   -16,    33,   -12,   -31,    -9,    -8,   -50,  -105,   -79,   -57,   -11,    -4,    22,   -19,   -26,   -52,   -66,   -13,   -17,   -36,   -41,   -34,   -28,   -24,   -31,     3,    -6,    10,   -24,    13,     8,   -53,   -48,   -43,  -101,   -60,   -57,   -26,     2,    23,     0,   -25,   -81,  -102,   -64,   -64,   -38,   -28,   -36,   -52,    -7,   -11,   -18,   -10,    -5,   -10,   -39,     9,   -14,   -40,   -52,   -61,   -61,   -67,     4,   -21,    19,    -6,   -16,   -26,   -54,   -89,   -65,   -51,   -31,   -15,   -21,    -3,   -13,   -32,   -13,     9,     7,    -6,   -23,    -8,   -10,   -33,   -38,    -2,   -19,   -20,   -13,    17,    23,   -17,     7,     4,    -1,   -15,   -19,   -11,   -63,   -36,    -7,    -5,    -2,   -34,   -11,     2,     0,     4,   -20,   -25,   -27,   -21,     6,    31,   -25,     9,   -15,    23,     5,     8,   -29,    15,    -1,    -9,     3,     5,   -40,   -73,   -61,    -6,     3,   -14,   -18,     2,     1,   -20,   -11,   -27,   -36,    21,    16,   -15,    10,   -19,    18,    35,    -3,   -11,   -17,    -5,    18,     6,   -26,   -46,   -48,   -64,   -27,   -18,   -11,   -10,   -28,     5,     5,   -18,   -23,     8,   -33,   -14,    -7,     9,     5,    -1,     6,    21,    13,     2,    11,    -9,   -24,    11,     6,   -39,   -59,   -34,   -15,   -24,     6,   -19,   -14,    -7,    -6,   -23,   -41,   -11,   -42,   -32,     4,    12,    -6,    46,   -23,   -17,   -44,   -29,   -22,   -29,   -40,    38,    25,     5,   -34,   -10,   -20,   -27,   -18,   -24,   -48,     7,    -7,    -8,    -6,    30,   -16,   -36,   -19,    -2,     7,    -2,   -17,   -39,   -29,     0,    16,    -1,    -1,    44,    65,    44,    -1,   -17,   -27,   -15,    -3,   -47,    -7,    -2,    -7,     5,   -24,    22,   -21,   -27,     4,   -35,    17,   -10,   -38,   -13,   -52,     0,    30,    11,    20,    53,    39,    35,     5,   -39,   -28,    -6,     2,    -5,   -18,    -6,    -5,   -13,   -26,    27,     2,    39,    19,   -14,    -7,     2,   -17,   -18,    -1,    52,    10,   -18,   -23,    -1,     9,     0,   -20,   -33,   -31,     3,    -4,    -7,     1,     6,    -7,   -28,   -23,    12,    -3,     2,     3,    31,   -30,    18,    41,    36,    24,    18,     2,    -7,   -27,   -26,   -36,   -50,   -43,   -32,   -12,    -3,    -7,     2,    -7,    -1,     0,   -12,     4,   -11,   -19,   -70,   -20,    33,   -14,     3,    35,    54,    22,   -37,   -41,   -20,   -46,   -35,   -39,   -39,   -10,   -10,   -29,   -20,   -29,     4,     7,    -9,    -9,     3,   -23,   -31,   -14,   -39,    23,    19,     8,    21,    33,    30,     7,    -8,   -22,   -10,   -59,   -47,   -36,    -3,   -10,    -2,     5,   -21,   -23,    -7,     5,     5,     7,    -5,    -4,   -14,   -18,   -10,   -11,   -27,   -24,   -11,   -21,   -11,   -25,    -9,    -9,    13,     1,    -3,   -28,   -10,   -14,   -11,     6,     2,   -12,     2,    -3,    -8,     9,    -7,    -7,     1,   -34,   -42,   -44,   -24,   -14,    -7,     2,     2,    -8,    -9,     4,   -12,    -3,    -9,   -10,   -31,   -11,    -9,   -17,     1,    -5,     3,    -7,     7,   -10,     0,    -4,    -6,   -17,   -15,   -12,   -10,     1,   -20,   -16,    -9,    -2,    -2,    -2,    -7,     3,     1,     5,   -21,    -8,   -15,    -1,     2,     7,    -7,     7,    -8,     4,     9,     6,     6,     8,    -8,    10,     9,     7,     6,     3,    -4,    -3,   -11,    -1,    -5,   -12,     4,    -3,   -10,   -15,     5,    -3,     1,    -8,     1,    -9),
		    77 => (    2,    -3,    -6,     4,     5,     1,   -10,     9,    -1,     2,    -6,     9,    -5,     9,     5,     3,     3,    -2,     1,    -7,    -7,   -10,     8,     6,     2,    -1,     8,     0,     6,     3,    -3,    -2,    -2,    -4,     1,     8,     5,    -2,   -13,    -2,    -4,    -7,   -11,   -35,   -44,   -28,     8,     8,    10,     1,    -1,     0,     5,     0,    -1,    10,     5,     8,     1,    -6,     1,     7,    -2,   -10,    -3,     0,   -26,   -16,    -3,    -6,    -7,    -9,    -1,     2,   -10,    -1,     0,    -4,     0,    -8,    -5,    -2,    -4,     7,    -3,     2,    -9,    -8,    -9,    -6,    -5,     6,   -24,   -24,   -22,   -29,   -15,   -22,     6,   -30,   -36,   -70,   -21,   -36,   -21,   -18,   -37,    -8,   -15,    -8,    -7,     8,     4,    -1,     5,    -6,   -27,   -13,   -23,   -67,   -54,   -46,   -64,   -98,  -112,   -84,   -59,  -110,   -81,   -93,   -86,   -51,   -55,   -21,   -74,   -43,   -26,   -20,    -8,    -8,    -9,    10,   -10,   -41,    -7,    53,    44,    31,    71,    68,     1,    28,    10,    23,   -16,    -2,   -10,   -38,    -2,   -22,   -40,   -82,   -84,   -61,   -80,   -68,   -20,    -8,     7,     0,    -6,   -23,   -15,    29,    38,    53,    57,    -1,    10,    33,    49,    50,    63,    15,    54,    40,    28,    32,    37,     9,    25,    -5,   -10,   -24,     1,   -19,     0,     7,   -13,    -7,   -23,   -18,   -26,    40,   -11,    10,    -6,    37,    60,    58,    23,    36,    23,    55,     6,    20,    30,    -3,     3,    -7,     9,   -10,   -14,   -10,   -26,    16,    -1,   -14,   -16,   -44,   -39,   -33,   -55,   -49,   -55,    -3,     6,   -16,     6,    12,    -6,    22,   -13,     2,   -36,   -20,   -44,   -42,   -41,   -16,   -28,   -32,     0,    -5,   -13,    10,     3,   -33,   -57,   -44,   -92,   -29,   -55,   -37,   -30,   -44,   -24,   -39,     4,   -45,     2,   -10,   -34,   -24,   -26,   -36,   -30,   -11,   -33,    19,    -5,   -16,   -37,   -33,    -2,   -39,     0,   -25,   -43,   -26,   -52,   -29,   -82,   -97,  -100,   -26,   -19,     8,   -15,   -23,    -5,   -69,   -18,   -56,   -38,   -18,   -39,    17,    -5,    -8,   -33,    -4,   -29,   -31,   -34,   -60,   -79,   -67,  -103,   -69,  -113,   -68,   -51,   -18,    -1,   -15,   -26,   -26,   -21,   -20,    28,    35,   -27,   -62,   -33,    28,    -1,     2,   -18,     9,    -2,   -28,   -43,   -82,   -68,   -94,   -65,   -81,   -63,   -41,   -34,   -12,    -3,   -47,   -58,   -22,   -30,     7,    10,   -12,    -3,    -3,   -20,    27,     8,    -4,    14,     0,   -13,   -31,   -20,     5,   -35,    -6,   -27,   -15,   -17,     0,    -6,     7,    21,   -25,     3,   -12,    33,    35,   -13,   -38,   -31,    -2,   -37,   -32,    -8,    -3,     0,   -14,    25,    -1,    17,    36,     0,     4,    11,    21,    31,    21,    21,    19,    21,     3,    19,    67,     1,     7,    18,   -69,   -42,   -25,   -25,     8,     2,     0,   -16,     6,    34,    27,    24,    39,    38,   -10,    17,    -3,   -17,     5,     1,    17,    44,    27,    -6,   -13,   -33,     7,   -25,   -80,   -82,   -52,    -9,   -19,     9,    -7,   -19,   -23,     7,     3,    -7,   -50,    -1,    -4,    -6,   -33,    -3,    10,     7,    37,    16,     0,    -4,   -12,     7,   -15,   -46,   -62,   -73,   -46,   -32,   -26,    -6,    -6,   -24,   -22,   -35,   -18,    28,   -36,   -15,    -6,   -15,    23,     2,   -20,    15,   -13,   -31,   -30,    -3,    -4,    24,    -9,     9,   -13,    13,    20,    38,   -52,     3,     3,    -9,   -24,     1,   -24,   -27,   -14,     0,   -45,   -28,    28,    13,   -18,   -11,   -11,   -79,   -53,   -10,     4,   -27,   -35,   -45,   -37,   -12,    27,    53,   -48,    -6,     5,     8,   -13,    22,   -33,    -6,   -59,   -63,   -14,   -28,     3,   -29,   -23,   -11,   -40,  -107,   -45,    -4,   -13,   -85,  -106,   -53,   -61,   -27,    35,   -26,   -16,     8,    12,    11,    -8,   -28,   -11,   -21,   -42,   -33,   -18,    -1,    23,   -28,   -25,   -20,   -46,   -62,   -31,   -85,   -81,   -32,   -44,   -51,   -25,   -59,   -68,   -15,    -8,    -4,     2,    -5,    -1,   -22,    22,     1,     7,   -17,     4,     5,    -3,    33,    14,   -23,   -12,   -32,   -14,   -48,   -35,   -68,   -45,   -21,   -14,   -31,   -33,   -11,     3,     4,    -4,   -14,   -13,    38,    -1,   -15,    13,    22,    -4,    -2,     4,    -2,    20,   -49,    -3,    23,    -3,   -22,   -61,   -79,   -50,   -12,    -2,   -49,   -15,   -23,     4,     5,    -6,   -14,   -66,    -6,   -45,     7,    -6,    -1,   -26,   -14,    -9,     2,    32,   -20,   -20,   -55,   -60,   -38,   -35,   -71,   -33,   -36,    -1,    -5,    -3,   -27,    -5,     0,    -2,   -15,   -43,   -19,   -33,    -3,    32,    19,     7,   -44,     5,    19,    26,    -8,    36,   -58,   -62,   -13,   -12,   -61,   -64,   -48,    10,    -9,   -34,   -16,     8,     7,    -9,    11,    17,    20,    10,   -46,    13,    25,   -52,    -8,    24,    30,   -22,   -13,   -42,   -72,   -37,   -21,   -26,   -41,   -29,   -15,    -2,     3,   -11,    -3,     2,    -2,     6,     2,   -35,   -11,   -28,    -4,    43,    44,    29,     2,     4,    34,    33,    40,     1,    -2,     3,     6,     9,     5,    -1,     2,    -2,     3,    -8,     8,    -6,     2,     0,    -6,     9,    12,     2,     3,    -6,    15,    -5,   -19,    -3,    11,    13,    10,     1,    -1,    -1,    13,     9,    -5,     0,     6,    15,     8,     7,     0,    -4),
		    78 => (   -9,    -7,     1,     8,     5,     9,    -3,    -2,     2,    -1,    -5,     9,     3,    -5,     8,     3,    -4,     6,     3,     3,    -7,     0,     8,    -7,    -9,     5,     6,     9,     5,     9,    -7,    -6,    -9,    -9,     0,    -1,     9,     5,    -2,    -7,     5,     3,    -5,   -27,   -49,   -36,    -3,     3,    -2,     0,     3,     8,    -5,    -9,    -6,     0,     7,    -8,    -1,     6,     9,     1,    -4,     3,   -14,   -25,   -57,   -41,   -14,    -8,   -11,    -1,     2,   -15,   -20,   -11,   -12,   -25,   -38,   -17,   -19,   -15,    -3,     4,     0,     1,   -16,    -3,    -4,   -33,   -21,   -50,    28,    16,   -11,   -17,    -3,   -17,   -32,   -18,   -10,   -25,    -5,   -13,   -16,   -14,     3,    10,    -1,   -13,   -26,     7,    -1,     5,     3,    -1,   -30,   -50,    -5,     1,   -13,   -48,   -46,   -58,   -17,   -17,    -5,   -41,   -17,    35,    36,   -20,   -15,   -23,   -32,   -26,    -5,   -19,    10,   -13,     8,    -9,    -6,    -5,   -29,   -39,    11,     8,   -28,   -53,   -40,   -30,   -35,    -9,   -15,    -2,     3,     7,    24,    13,     4,     0,   -17,    -8,    -5,   -11,    -8,   -28,     2,     8,   -25,   -47,    -9,   -39,     1,     8,    -3,    -4,   -30,   -27,     6,     8,    -3,    18,    -9,    -5,     4,     1,     6,     0,     7,    -3,    -2,    -3,    -7,     5,     2,   -41,   -19,    -3,   -25,   -17,    13,    -1,     8,     9,    20,    -2,     4,   -28,    -4,    35,     8,    -8,    29,   -25,    -6,    -4,   -11,   -20,   -14,   -17,   -10,   -10,   -17,   -21,   -19,     1,   -24,   -16,    20,     1,    -6,    -3,     9,    -4,   -14,   -17,    -3,    34,    18,   -38,     8,   -10,   -37,   -14,   -10,     4,    -6,    14,    -3,     4,     0,   -15,   -39,     1,    -9,   -50,    10,   -12,    11,    -4,    -4,   -34,   -24,   -13,    -7,    29,    12,   -37,    12,     1,    -8,    -2,    -2,   -16,   -31,    -6,   -22,   -49,     3,   -12,   -36,     9,   -10,   -45,   -42,     5,    -5,   -30,     7,     2,   -10,   -33,   -42,    14,   -25,    11,     4,     1,    -8,   -22,   -23,   -39,   -30,   -10,    29,   -35,     2,     5,   -18,    -2,   -23,   -43,   -39,    13,   -12,   -37,   -13,   -24,   -37,   -48,   -15,    24,    -3,     1,    22,    11,   -13,   -46,   -28,    18,    -2,    -1,    40,   -40,    -8,     6,   -25,   -22,   -33,   -23,   -28,    -2,    -2,   -26,   -26,   -24,   -19,   -42,   -41,    25,    20,    10,    20,    10,    -2,     7,    14,   -25,   -15,   -21,   -15,   -59,    -6,     0,   -35,   -22,   -39,   -36,   -28,    -8,   -16,     2,   -52,   -35,   -53,   -57,   -25,    -2,   -12,     5,    31,    11,     4,    13,   -15,   -21,   -26,   -33,   -32,     1,     3,    -3,     4,   -21,    -5,   -21,   -47,   -19,   -12,     1,    -3,   -16,    -7,   -71,   -19,   -25,   -49,   -29,   -17,     3,    -2,   -11,   -33,   -32,   -28,    -9,   -92,   -12,     0,     8,    -1,   -15,     1,    -3,   -25,   -27,   -21,     7,    -2,   -28,    -6,   -52,    -3,     3,   -19,    -3,   -14,   -19,   -15,   -11,   -19,   -26,   -12,    -6,   -81,   -30,    -2,    -4,    -6,   -12,     5,   -14,   -16,    -2,   -11,   -26,   -14,   -16,   -30,   -13,    15,     0,   -17,     4,   -16,   -20,   -21,   -10,   -25,   -18,   -11,     1,   -45,   -31,     6,    -1,    -6,   -11,    -3,   -15,   -20,   -10,   -19,   -45,   -44,   -32,   -50,     7,    25,    16,   -14,   -31,    -8,    -5,    -3,   -13,   -21,   -11,    -1,    -7,     0,   -31,     2,     4,     0,   -21,    -1,   -16,   -12,     0,   -24,   -35,   -10,   -38,    -3,    18,     9,    -4,     9,   -33,     2,    -9,   -16,   -31,    -6,   -13,     8,    -5,     1,   -17,     2,    -8,   -29,   -29,     5,   -13,    -9,   -28,   -45,     0,   -12,   -19,    15,    15,     0,    26,    30,   -12,    -6,   -15,   -25,   -13,   -13,    -5,    -4,     0,   -46,   -39,     1,     4,   -10,    -5,     4,   -29,   -21,   -17,   -22,    15,    -4,   -16,    -8,   -15,   -33,     2,    -8,    19,     4,   -11,   -43,   -27,   -26,   -12,     3,    -9,   -36,     9,   -35,   -15,   -13,    -2,   -20,   -37,   -27,   -48,    -2,    31,    -2,   -38,     7,   -16,   -33,   -43,     0,    38,     7,     8,   -22,    -7,   -18,   -15,   -15,     2,   -43,    -1,   -18,   -18,    -5,   -16,    -5,   -32,   -14,   -21,   -12,    21,    17,     9,     7,   -16,   -32,   -34,    25,    23,     2,    -6,   -13,   -38,   -31,   -16,   -16,    -8,   -29,     6,     2,     4,   -14,    -3,   -14,   -27,   -24,   -18,   -27,    -1,    20,    18,    53,    16,     6,     0,    49,     1,   -12,   -48,   -22,   -16,   -23,   -10,   -12,    -3,   -50,     5,     3,    -6,    -7,   -13,    -2,   -13,   -31,   -22,   -27,   -15,   -22,   -24,     6,    -2,     8,    10,    23,   -48,   -46,   -40,   -36,   -15,    -4,   -10,   -34,    -9,    -8,     3,    -3,     8,   -26,   -21,    -7,     1,   -15,   -31,   -29,   -28,   -28,   -69,    -9,    11,     5,    29,   -47,   -67,   -46,   -30,    -5,   -13,     1,     4,    -2,   -18,   -17,     4,    -2,     4,     9,    -8,     6,   -23,   -22,   -16,    -1,   -26,   -38,   -47,   -40,   -54,   -73,   -35,   -16,    -2,    -5,   -14,   -55,   -32,   -28,    -8,     2,     9,    -1,     4,     7,    -8,    -3,    -4,    -8,    -2,   -16,     2,   -12,    -6,   -13,     1,     6,   -22,    -2,    -5,   -27,   -33,     0,     4,   -10,    -6,    -6,   -10,     1,    -5,     7,     7),
		    79 => (    1,     0,     8,    -1,    -3,    10,    -9,     2,     3,    -8,    -5,     2,     9,     5,     5,     5,     6,    -9,    -1,     0,     2,     0,     4,    -3,     0,     9,     4,    -4,     5,     6,    -1,     0,     7,     5,    10,     7,    10,     8,     1,   -15,   -18,   -15,     5,     4,     4,    -4,    -4,     3,   -10,     0,     5,     7,    -7,     1,     8,    -7,    -2,    -5,     5,    -6,     9,     0,    -7,    -2,    -3,   -14,   -10,   -11,    -4,    -9,   -20,    -8,    -9,    -7,    -7,    -6,    -1,     5,     6,     6,     0,     0,    -1,     4,     1,    -2,    -6,     3,     8,    -7,    -7,   -10,   -18,   -11,   -25,   -44,    -9,   -26,   -36,   -29,   -35,    -5,    18,    30,   -19,   -11,   -22,   -11,    -3,     0,     9,     2,     1,     7,     5,     2,     1,    -8,   -39,   -11,   -11,   -30,   -34,    35,    24,    26,     2,   -29,   -33,   -51,   -65,   -58,   -68,   -31,   -25,     7,     3,   -36,   -21,    -8,    -8,     4,     1,    -9,     0,     1,    -7,   -17,   -64,   -80,   -52,    52,    -1,     6,   -14,    22,    70,   -23,   -10,   -12,    24,   -35,   -38,   -17,   -25,   -34,   -38,    -5,     0,   -29,   -11,    -1,   -10,   -43,    -5,   -65,   -25,   -35,   -21,   -29,    20,    21,    37,    21,    10,    18,   -21,   -49,   -58,   -11,   -27,   -18,    -9,   -18,   -23,   -16,    10,    -8,   -16,     5,    -8,   -64,   -61,  -120,    44,   -74,    16,    45,    24,    19,    18,   -23,   -20,   -60,  -113,   -54,   -31,   -27,   -25,   -25,   -14,   -15,   -21,   -20,   -17,   -51,   -19,   -12,   -19,   -39,   -80,   -89,    56,   -17,    40,    48,    42,   -27,   -71,   -13,   -50,   -15,   -39,    23,   -13,   -32,   -17,   -34,   -36,   -25,   -63,     0,     0,   -34,   -18,   -10,   -49,   -46,  -113,   -19,    48,     1,    27,     4,   -58,   -53,   -40,     3,   -11,    21,   -42,    17,    -7,   -40,     9,   -25,   -17,   -44,   -27,   -13,     3,   -12,     3,     6,   -25,   -21,   -48,    30,    53,    35,   -24,    11,   -39,    21,    75,    47,     0,    35,    52,    29,   -35,   -80,   -34,   -51,   -22,   -33,    -4,   -32,   -10,   -21,     1,    -8,   -22,   -28,   -14,    -1,    33,     9,     5,     4,    41,    52,    69,    25,    44,    56,    14,     2,   -32,   -38,   -51,   -44,    -9,   -38,     2,   -28,    10,    -4,   -15,     2,   -11,   -27,   -48,   -25,   -13,   -16,   -13,    12,     0,    37,     1,     5,    15,    19,     1,    10,   -20,   -25,    -2,   -75,   -72,   -28,   -39,   -11,     5,   -13,   -12,   -42,   -26,   -25,   -47,   -10,   -19,    11,   -43,   -15,    -8,    25,    -3,    49,    39,     1,   -79,   -31,   -39,   -53,   -13,   -29,   -37,   -24,   -38,     1,    -3,   -10,   -25,   -32,   -23,   -24,   -49,   -20,   -64,    -9,   -42,   -26,    -6,    25,   -27,   -13,    15,    10,   -33,   -55,   -36,   -10,    29,   -12,    -3,   -33,   -14,    -9,     6,     8,    -9,   -26,    -5,   -18,   -14,  -100,   -85,     3,    22,    37,    34,    -9,    -7,   -40,    19,    18,   -68,   -55,   -69,    10,    24,   -17,     8,   -20,   -16,   -22,    -5,    -7,   -19,   -13,    -2,   -20,   -21,   -51,  -117,  -102,   -59,    -1,   -13,   -63,   -42,   -37,    -4,   -36,   -32,   -89,   -57,   -15,    16,    -3,    11,   -26,     4,   -10,    -1,    -5,   -27,     2,     3,    22,    17,   -25,   -39,   -76,   -97,  -149,   -79,   -47,   -19,   -30,   -20,   -28,   -38,   -80,   -46,   -16,   -40,   -39,    22,   -10,   -15,   -11,    33,     7,   -23,   -15,   -16,   -34,   -25,   -29,   -40,   -46,   -65,  -125,   -52,   -28,   -19,   -46,   -20,   -11,   -44,   -69,   -95,   -40,   -44,   -62,   -30,    -4,    -9,   -19,     9,   -17,    -6,    -1,   -10,   -53,   -64,    39,   -36,   -49,   -58,   -81,   -24,   -24,   -13,   -24,   -31,   -52,   -24,     1,   -72,    12,    -4,   -12,   -19,   -15,   -20,    10,    -1,   -18,   -12,   -10,   -13,    12,   -44,    14,    16,   -21,     3,   -27,   -15,   -17,   -30,   -46,   -30,   -39,    -4,   -20,   -63,     1,    22,    -4,    40,    11,    -6,     2,    -1,     7,   -26,   -15,    21,    31,   -59,     2,    33,    64,    17,    -6,   -13,   -13,   -54,   -42,   -51,    -8,    -4,     2,   -18,   -30,    -8,    38,    25,    27,   -32,     1,     6,    -9,   -56,   -32,     0,   -18,   -63,   -41,    32,    42,     2,    33,     4,    -2,    -8,   -28,    -4,   -11,    20,     8,    -6,   -25,   -21,    18,    52,   -43,    -9,    -8,     7,     9,    -3,   -25,    -5,   -35,   -36,   -50,     2,    33,    28,    46,    21,    21,    27,    19,    -4,   -10,    21,    -6,    14,   -45,    17,    12,    39,   -13,    -7,     5,    -5,     1,    -4,   -52,     1,     1,   -12,    -1,    17,    -4,    20,    -7,   -38,   -24,    -2,   -14,    12,    -2,   -40,   -52,    27,    -2,     2,    10,    -4,    -8,   -10,    -6,     0,    -4,    16,   -20,     2,    -1,    27,    45,    -2,    13,   -29,   -35,   -36,   -39,   -15,     2,     8,    40,   -44,   -57,    31,     8,    26,    26,    -2,    -6,     4,    -3,     2,    10,    -3,    23,     9,    -4,   -16,     7,   -77,    -5,    41,    17,    -7,    -6,    60,   -19,   -62,   -48,   -28,   -36,    -7,     4,   -12,    14,    16,    -5,    -9,    -5,    -1,     9,     9,    -8,   -16,   -13,     6,     9,   -17,   -22,    -9,    27,     4,   -17,     1,    28,    53,   -33,     4,     0,     4,   -12,    -7,     3,    -8,     7,     6,    -5),
		    80 => (    1,    10,   -10,    10,    -5,     4,     2,    -7,    -7,    -8,    -2,     5,    -7,     8,     5,    10,    -9,    -9,    10,     8,     0,    10,    -4,     0,    -3,    -8,    -9,     5,    -5,     9,     6,    -4,    10,     9,    -3,    10,    -3,    -8,    -9,     6,     5,    11,   -16,    -6,     6,     3,   -12,    -3,     1,     2,     0,     1,    -2,    -6,    -7,    -1,    -7,     2,   -10,    61,    55,     0,     7,    12,   -10,   -16,    -6,   -44,   -37,   -62,   -67,   -61,   -38,   -45,   -35,   -44,   -33,   -36,   -41,   -26,   -35,   -17,    -3,    -6,    -6,    -2,     9,    73,    44,    23,   -12,   -18,   -31,   -26,   -28,   -16,   -22,    28,     8,   -20,     7,   -12,   -16,    -4,    10,   -67,   -48,   -41,    -1,   -11,   -33,    -8,    -1,     3,    -6,    -3,   -16,   -21,   -30,   -33,   -31,   -18,   -20,   -27,   -46,   -21,   -12,    10,   -26,     6,    35,    13,    36,    22,    68,   -20,    -2,   -24,   -40,    -5,     1,     5,   -13,    12,     7,     4,    13,   -57,   -70,   -58,   -63,   -90,   -51,     0,   -10,   -10,   -19,    20,    21,    18,    47,    29,    73,   -12,    -5,   -28,   -36,   -17,    -9,     5,   -14,   -11,    10,    48,     7,     7,   -50,   -91,   -77,   -81,   -13,    39,    -1,    11,   -55,   -21,     2,     6,    -9,    54,    38,   -38,   -66,   -81,   -45,     0,    -7,    -4,    -7,   -17,    27,    55,    10,   -18,   -31,   -21,   -30,    10,     1,     5,   -34,    -8,   -17,   -14,    -3,    29,    16,   -32,    25,    19,   -13,   -17,   -58,    18,    23,   -19,    23,   -19,     6,    34,    24,   -24,   -28,   -42,   -65,   -59,   -23,   -21,    36,   -29,    15,   -10,    18,    11,     9,    35,    33,    21,   -42,   -56,   -60,   -11,    -3,    -6,    28,    -7,   -25,    32,   -21,   -33,   -16,   -80,   -26,   -52,   -19,   -11,    35,    19,   -37,    -7,    14,    -1,    18,    -9,    16,    41,    35,    11,   -42,     5,     4,    -2,    15,    -3,   -40,   -16,   -66,   -25,   -31,    10,   -29,   -11,    31,    -5,     7,    23,     2,   -35,   -60,   -23,    50,    33,    43,    39,    36,    15,   -74,    -8,    -7,    28,   -23,   -20,   -47,   -47,   -35,    31,     9,    -9,   -20,     6,     6,   -25,   -12,   -33,   -75,   -92,   -88,    -1,    15,    18,     1,    -3,   -11,    -2,   -41,    -5,     9,    25,    -9,   -13,   -20,   -35,   -34,    -5,    -8,   -11,    27,    31,    29,    34,    17,   -17,  -132,  -120,   -29,    24,   -39,   -11,    17,    65,    -7,   -15,   -34,     0,     9,    21,    17,   -33,   -25,   -22,     1,    10,    12,    23,     6,    29,    19,    23,     3,   -36,  -159,   -59,    31,    -4,   -34,   -43,     5,   125,    37,    28,   -32,    -8,     2,    -3,    -1,   -84,   -22,   -11,    15,    41,     1,    14,   -36,    -2,   -10,   -17,  -133,  -111,  -120,   -50,   -27,   -24,   -23,    12,     9,    55,    18,   -15,   -58,    -2,     2,     5,   -19,   -90,    13,   -30,     4,    47,    14,    17,   -53,   -21,    29,    -4,   -94,   -62,   -19,    -2,   -32,   -20,   -65,     9,    12,    35,    58,   -38,   -66,   -17,    10,     7,    -1,   -65,    17,    -2,    -2,    42,    28,   -25,   -25,     4,   -38,   -63,   -25,    -8,     3,   -17,    12,   -35,   -15,   -35,   -15,     4,    34,   -52,   -28,     5,    -1,   -10,   -28,   -31,    11,    39,    17,    44,   -21,    14,    -1,   -29,   -86,   -61,   -37,   -10,   -29,    -1,    -5,    17,    17,   -44,   -31,    11,    30,   -57,   -30,     5,   -10,     5,   -20,    -5,    19,     6,    13,    39,    54,    25,   -46,   -86,   -67,   -28,     2,     7,   -10,    -2,    16,   -32,    -5,   -13,    16,     8,     6,   -27,   -17,   -13,    10,    12,   -54,   -17,    63,    -3,     4,    29,    13,    26,   -41,   -79,   -34,   -43,    -2,    12,   -33,     9,   -25,   -17,   -49,   -13,    17,    -1,    23,   -37,    -7,     8,     3,    14,   -75,    18,    53,    11,    27,    -7,    20,    17,    -9,    15,   -16,   -21,   -10,   -54,   -12,   -14,   -14,   -52,   -59,   -20,     7,    -7,     7,   -32,    10,    10,     4,     9,   -74,    20,    11,     9,    30,    44,    11,    21,     2,    -2,   -27,   -18,     3,    23,     1,    -7,   -40,   -50,   -70,   -73,   -44,   -12,    38,   -20,     9,    14,     4,    -8,   -83,     0,    -2,    37,    47,    19,    17,    14,    18,   -24,   -29,     7,    31,     2,   -70,   -55,   -24,   -29,   -84,   -50,    -9,    -6,    32,     4,     1,    11,     8,     0,   -13,   -59,   -67,    10,     7,     1,     9,    28,    33,    29,     3,    23,    24,   -43,   -66,   -42,   -61,   -56,   -80,   -37,    14,     2,   -47,     0,    -5,    -7,     0,    -4,   -18,   -13,    58,    75,    -4,   -17,     6,    40,    67,    43,    60,   -63,   -55,   -57,  -115,   -98,   -55,   -59,   -29,     7,    -8,    -2,    24,     6,    -4,    -9,     6,    -9,     1,    -1,   -39,   -76,   -70,   -71,   -60,   -38,   -50,   -61,   -82,   -60,   -24,   -67,   -70,   -64,   -78,   -56,    -4,   -15,   -13,   -12,    -2,    -1,    -8,     4,     9,     5,    -6,    -9,    -8,   -56,   -76,   -18,    -1,   -19,   -32,   -37,   -20,   -28,   -22,   -41,   -43,   -72,   -77,   -17,   -47,   -20,   -20,   -11,     0,     5,    -8,     5,    -8,   -10,     9,     8,     1,     5,     7,    -9,    -3,    -1,     2,     7,     7,    -4,     1,    -1,    -4,     4,    -1,   -13,    -8,   -13,   -13,   -10,     1,     0,     8,    -7),
		    81 => (   -8,     4,     9,     9,    -6,    -6,     1,    -8,    -9,     5,    -4,     9,     2,    -3,     9,    -2,     4,    -1,     6,    -1,     6,    -2,     8,    -2,    -9,     7,    -7,     8,    -4,     3,     6,     0,     1,    -9,     1,    -2,     2,     9,    -1,    -6,    -2,   -15,    10,    13,    -5,   -14,     1,    -8,    -3,    -1,    -5,     5,     5,    -3,     5,    -6,    -6,     5,    -7,     9,    -2,     7,    -1,   -10,   -12,   -11,   -11,    -8,     0,     2,    51,    62,   132,    98,    49,   -32,     8,   -44,   -33,   -25,    -4,     7,     8,    -5,    -3,     0,    23,    18,   -10,   -34,   -69,   -23,    44,    14,   -28,   -50,   -42,   -10,    21,    73,    82,    16,     3,   -35,     2,    45,   -10,    -2,   -34,    -1,     5,    -4,     6,     9,    25,    22,    47,    21,   -14,   -18,    69,    53,    32,    -6,    -5,   -29,    -7,    19,    24,    13,   -16,   -16,    35,    46,    21,    34,    -6,   -25,   -23,   -32,    -2,    -9,    -5,    -7,    54,   105,    45,    39,    27,    11,     8,   -52,   -53,    10,    33,     8,   -17,     9,     3,    18,    34,    36,    31,    11,     6,   -12,   -29,   -29,     7,     4,   -67,     5,     9,    22,    45,    15,   -31,   -39,    21,   -11,    -1,    -9,    -6,   -11,   -39,    28,    14,    49,    28,    -8,    13,    -5,    -4,    -6,   -15,    -7,   -10,     7,   -75,   -66,   -65,    -4,    25,    31,   -50,    10,    35,   -29,    -6,   -43,    -9,    28,    -9,    10,    27,    54,     9,    -5,    18,   -15,   -17,     1,   -31,   -17,    -3,    -6,   -84,   -51,   -62,   -11,    12,     2,   -14,    24,    13,    10,    22,   -41,   -43,     9,    30,     4,    31,   -43,   -26,   -21,    11,   -27,    -3,    -3,   -32,    -6,     4,    -4,   -82,   -33,   -41,   -44,     1,    22,    36,     5,     8,    62,    49,   -30,   -55,   -16,   -29,   -30,   -31,   -22,   -18,   -22,   -31,     0,   -11,     6,     5,   -11,     2,    -3,   -64,   -11,   -72,   -36,   -65,     7,    27,    42,    18,    67,    17,   -17,   -28,   -18,   -42,   -33,   -13,   -60,   -38,   -44,    -3,    -6,   -12,    -9,    12,     2,    -2,    13,   -14,    -6,   -60,   -33,   -57,     1,   -28,    19,     5,    36,    14,   -14,    -8,   -41,     5,   -44,   -40,   -53,   -34,   -26,     7,     1,    -9,    -7,    -6,    10,    -5,    -4,    -9,   -22,   -42,   -43,    19,    37,     8,     3,   -19,     6,    -4,   -33,   -43,   -11,   -13,   -47,   -18,   -54,   -79,   -35,   -19,   -18,   -10,   -13,     6,    17,     0,    -2,   -11,    -9,   -56,    22,    37,    38,    52,   -21,   -29,    -2,   -11,   -45,   -19,    27,   -14,   -33,   -37,  -115,   -53,   -45,   -38,   -33,   -29,    -3,    -4,    -2,    -5,     0,     6,    -2,   -48,    42,    35,    -9,   -16,   -66,   -86,   -49,   -31,   -27,    13,    18,    -2,   -29,   -47,   -76,   -68,   -79,   -52,   -34,   -20,   -31,     3,     6,    -9,     6,    -3,    15,    -9,   -39,   -24,   -24,   -45,   -58,   -73,   -76,   -88,    -7,    38,     8,   -11,   -32,   -45,  -101,   -57,   -60,   -48,   -50,  -116,   -17,    -5,   -13,     5,    -3,    13,   -24,   -21,   -22,   -35,   -34,   -77,   -42,   -46,   -81,   -70,    -7,    50,    37,   -12,   -44,   -36,   -78,   -68,   -83,   -29,   -57,   -39,   -15,   -10,   -16,    -5,    -4,    -4,   -42,   -11,   -19,   -33,   -59,   -59,   -57,   -64,  -138,   -77,   -62,    23,   -22,   -20,   -24,     3,   -30,   -40,   -30,     0,   -33,   -61,   -65,    -5,   -23,   -12,     5,     6,   -11,   -11,   -50,   -97,   -56,   -97,   -64,   -70,  -176,  -153,   -86,     0,   -30,   -13,    12,   -15,   -13,    34,    22,    51,   -23,  -115,   -26,   -26,   -21,    -3,     0,   -11,   -22,   -34,   -89,   -51,   -12,    -4,   -35,   -48,   -84,   -54,   -42,   -29,    21,    42,     6,   -37,    -3,    17,     0,    -5,    22,    -6,    -4,   -39,   -12,     6,    -9,   -25,    33,    -3,   -67,   -28,    11,    13,    29,    58,     8,   -14,     5,    21,    19,    55,    33,    79,    59,    49,    -3,    19,    24,    13,     7,   -30,     7,    21,    10,   -34,    35,    43,    16,    46,    40,    50,    49,    27,    28,    -3,    19,    19,    44,    12,    46,    75,    23,    28,    -6,   -37,   -20,    16,    33,   -38,     8,    22,     5,   -95,   -58,    29,    69,    23,     5,    12,    20,    21,    16,    11,    18,    -6,    15,   -17,    18,    10,    41,    44,    22,   -74,   -47,    10,    -7,    -4,     2,     9,     5,    -9,   -27,    14,   -14,    23,   -11,    -5,   -18,   -26,     4,     4,    30,   -35,   -55,   -75,   -61,   -20,    12,    35,    41,   -17,   -41,   -41,   -51,    25,     6,     1,     0,    -8,     1,   -17,   -28,   -39,    -8,    12,    23,   -12,    -8,   -70,   -46,   -91,   -75,   -69,   -42,   -27,    -8,    10,    17,   -23,   -31,   -44,    -7,     1,     8,     0,    -4,     9,   -11,    -4,    -6,   -19,    -7,    -6,   -44,   -20,   -28,   -40,   -47,   -31,   -60,   -45,   -52,   -62,   -52,   -62,   -51,   -40,   -18,     0,     5,     2,    -7,    -8,     9,    -6,     2,   -15,   -17,   -20,   -16,   -12,   -43,     2,    -7,   -21,   -33,   -23,   -41,   -11,   -43,   -25,   -36,   -26,   -21,   -14,     4,    -8,    -5,     7,    -4,     5,    -5,    -3,    -8,     0,     9,     2,    -3,    -2,    -5,   -15,   -15,    -2,   -12,   -10,   -12,   -12,    -9,    -8,    -2,     1,     1,    -4,    -1,     4,     6,    -4,    10),
		    82 => (    2,     2,    -7,    -6,     0,    -4,     4,    -9,    10,     0,    -1,     2,    -9,    -1,    12,     9,    -3,     2,    -6,     5,    -4,   -10,     7,    -3,   -10,     4,    -2,    -2,     1,     9,     9,    -2,    -8,     9,     6,   -23,   -38,   -15,   -35,   -32,   -38,   -68,   -29,     4,    33,     5,   -39,   -74,   -49,   -26,   -37,   -12,    -3,    -6,    -3,     3,     6,     9,    -1,   -53,   -55,     8,    -3,    -9,     0,    62,    53,    24,    14,    17,     8,    25,    -1,    -6,   -29,   -48,   -29,   -22,   -17,    -2,     9,    11,    -1,     1,    -2,    -5,    -3,   -59,   -75,    -9,    -2,    20,   -22,    25,    11,     9,   -17,    20,    43,    23,    23,     5,   -26,   -32,   -21,     8,   -39,   -95,    10,    13,     5,     1,    -1,     6,   -15,    16,    15,   -25,     7,   -10,   -50,    24,    50,     7,     7,    29,    38,    13,    22,    12,    51,     6,    -2,   -17,   -45,   -22,   -30,   -10,   -21,    -1,     0,    -9,    14,    -4,    -5,    13,    14,   -47,    -5,    13,   -32,   -22,    12,     0,     0,    -9,    34,   -14,     9,   -24,   -15,   -14,   -29,   -16,   -65,    -2,   -26,   -21,    -4,     3,     5,   -23,   -25,     4,     2,    37,   -33,   -28,    11,   -19,   -43,    40,    -3,    11,    46,     7,    14,   -38,   -21,    -4,   -24,   -34,   -79,    32,   -16,   -11,    -8,     5,    -8,   -22,   -24,   -10,    23,     0,   -33,   -28,    28,     7,    -2,   -31,     2,    22,    -2,     7,   -54,   -12,    23,    36,    -7,   -79,   -30,    10,   -39,   -18,   -16,    15,   -16,   -34,   -20,   -49,   -29,     2,    20,    16,    39,    22,   -46,   -28,   -56,    -4,    -1,    10,    18,    38,     3,     7,     3,   -37,   -66,   -80,   -30,   -12,    -2,   -16,    -8,   -28,   -18,   -66,   -56,   -71,   -86,   -23,     3,   -45,   -68,    -4,    -8,   -41,   -10,    15,    28,   -29,   -12,    44,    -2,   -36,   -35,   -42,   -28,   -24,    -8,     4,    -8,   -45,   -46,   -64,   -72,  -138,  -196,  -177,  -143,  -115,   -35,   -43,    -8,   -46,     4,   -19,    19,     3,    -4,   -15,    -4,   -18,   -60,   -48,   -22,   -10,    -2,   -27,   -26,   -53,   -53,   -66,   -98,  -119,  -157,  -134,  -113,   -62,   -47,   -65,   -15,   -44,   -31,   -71,   -69,     2,    -2,     5,    22,   -19,   -59,    -7,   -24,   -18,    10,   -31,   -66,   -50,   -83,   -61,   -56,   -73,   -20,   -18,   -11,    13,    -9,   -12,     9,   -29,   -52,   -62,   -45,   -24,   -13,    19,    44,   -49,   -49,    57,     7,   -13,    -9,   -29,     4,   -18,   -40,   -29,     9,    75,    32,    -8,   -19,    15,    72,    49,    20,    11,    -2,     2,   -27,   -34,    -5,    27,    58,    -4,   -11,    25,    -4,    -1,    -1,   -30,   -41,    50,    32,    -7,    50,    76,    63,    44,    62,    48,    40,    64,    57,    -7,    31,   -53,   -28,   -10,    23,    -4,    11,    11,   -11,    35,    30,    28,     1,   -18,    10,   116,    50,    62,    37,    35,    30,    32,    54,    19,    30,    16,   -27,    20,   -10,     9,   -23,    -2,   -29,   -18,   -12,    33,    -7,    48,    89,    55,    -2,     3,    10,    47,   -17,    61,    93,    43,    19,    29,    36,     5,   -34,    20,    21,    17,    13,    17,    -5,     2,   -29,   -35,   -19,   -14,   -40,    67,    89,    36,     7,   -14,     6,   -26,    26,    18,    61,   -17,    28,   -23,   -31,    14,     1,   -11,    44,    30,    30,     5,    -2,   -29,    -6,   -68,   -48,   -56,   -73,    10,    20,    59,     6,    -7,   -36,    12,    -4,    45,    47,     0,    -1,   -21,   -31,   -17,    -2,    12,   -11,    -2,    32,     9,    29,    41,    22,   -19,   -32,   -28,    11,    45,    25,    56,     4,   -34,   -34,   -14,    28,    27,    33,    28,    16,     8,   -27,     7,     2,   -11,   -29,    -7,     9,    -2,    35,    41,     6,    33,    35,    15,    53,    50,    41,    29,    -6,   -39,     3,    -5,    20,    63,    21,     3,   -10,   -36,   -21,   -41,   -53,   -46,   -47,    -9,    -1,   -38,   -26,    -7,   -12,    -1,   -15,    12,    61,    -9,    17,    -3,   -10,    26,     0,    15,    26,    19,    16,    16,    25,   -32,   -38,   -10,   -12,   -48,   -34,   -31,   -36,   -12,   -32,    -2,    24,    40,    17,    34,    18,   -33,   -22,    -5,    -9,    -6,    -4,    13,    30,   -30,   -27,   -12,    -9,   -30,   -10,     8,   -18,   -43,   -57,   -21,   -36,   -42,   -55,    -9,     4,     9,   -13,   -19,   -23,   -58,   -63,    -7,    -7,   -10,    15,    51,    46,     8,   -51,   -11,   -33,   -60,   -18,   -37,    -5,   -74,   -40,   -67,   -25,   -34,   -45,   -77,   -37,    -2,    30,   -48,   -45,   -34,   -42,     7,     4,     7,   -27,   -19,   -19,    -8,   -18,   -39,   -47,   -79,   -93,   -69,   -55,   -89,   -68,   -57,   -56,   -24,   -35,   -77,   -94,   -54,   -86,   -53,    14,    26,    26,     2,     1,     3,   -13,     2,   -19,   -16,   -12,   -27,   -54,   -71,   -25,   -16,   -23,   -64,   -50,   -32,   -48,   -60,   -38,   -80,   -60,   -36,   -47,   -17,   -19,    16,    34,     0,     4,     7,    -4,     4,   -18,   -27,   -24,   -18,   -21,    -9,    -7,    -6,     0,    -2,   -26,   -13,   -64,   -49,   -40,   -27,   -15,   -13,    -8,   -20,     9,     0,    -4,     0,     8,    10,    -1,    -2,    -6,     0,     2,    -8,     3,     8,   -19,    -8,    -8,   -18,    -3,    -6,    -5,     0,   -13,   -14,   -23,   -29,   -18,    -7,    -1,    -2,    -6,    -7),
		    83 => (    9,     2,     5,     6,    -4,    -4,    -8,    -9,    -7,    -1,    -4,    -7,    -3,    -1,   -15,   -13,    -4,    -4,     5,     1,     8,    -1,     6,     9,     3,    -8,     6,     9,     0,     5,     2,    -6,     6,    -8,     2,    -8,   -10,    -2,   -17,   -12,   -14,   -44,   -33,   -32,   -17,   -49,   -24,   -26,   -14,   -11,   -11,    -3,    10,     5,    -8,    -9,    -3,     3,    -2,    -1,   -22,   -19,   -24,   -26,   -49,   -63,    24,    -3,   -22,   -39,   -52,   -51,   -35,    -5,     7,   -44,   -60,   -79,   -72,   -60,   -11,    10,    -8,     3,    -6,     7,   -11,   -13,   -11,    23,    42,   114,   108,    42,    47,    45,    34,    14,    -8,    55,    71,    47,    41,    93,   165,    16,  -103,  -107,   -54,   -30,     2,     3,     9,    -5,   -65,     3,    22,    33,    13,    69,    88,    -1,    49,    23,    26,    -8,    19,     1,    31,    49,    40,    42,    17,   -55,   -56,  -211,  -163,   -61,   -43,     5,     3,     9,    -9,    -5,    -7,    35,    79,    98,    10,    23,    37,   -17,   -32,     5,   -19,    -5,    45,   -25,   -10,    28,     8,   -12,   -16,    14,    17,   -79,   -36,     4,     5,    12,    22,    -4,   -10,    69,   106,    88,    42,    44,    20,     3,   -27,    15,    -4,    30,    25,    10,    11,    -6,     4,   -13,    -2,    10,    34,   -93,   -44,   -15,    -3,     6,     2,    19,    -9,    15,    99,   127,    66,     4,     9,    59,     9,   -34,    10,    -2,    24,   -17,   -32,    18,   -16,   -18,   -27,   -12,    28,   -83,   -52,   -24,   -29,   -10,   -39,    -3,    17,    71,    12,    34,     9,   -15,   -12,   -46,   -56,   -33,   -14,    53,    26,    33,   -41,    28,     8,   -36,    24,     4,   -25,   -55,   -51,    -3,    -1,   -21,   -97,   -21,   102,    98,    43,    44,    51,   -24,    20,   -32,   -26,   -16,   -26,   -24,     5,    56,    27,    -9,    18,   -22,    59,    47,  -113,   -48,   -35,     6,   -10,    -4,  -107,     6,    22,    50,    61,    77,     0,   -21,   -50,   -59,   -32,   -51,   -16,   -27,    -4,    34,    41,    16,   -44,   -35,    19,    73,   -51,   -54,   -42,     1,    -9,   -38,   -49,    56,    87,    82,    50,    20,    37,   -21,    -9,   -46,   -47,   -15,    -3,   -43,     7,    10,    22,   -39,   -53,   -26,     4,   -22,  -136,   -95,   -45,   -10,   -10,   -12,   -50,    22,    57,    82,    58,    30,     9,   -34,    16,   -21,   -28,   -30,   -34,     8,    10,    -4,     9,    18,   -28,   -61,   -26,     4,   -86,   -59,   -20,    -6,     9,   -14,   -43,     3,    88,    61,    38,    29,    68,    -6,    26,   -21,   -29,   -10,   -19,    37,   -93,   -26,    43,    36,   -31,   -34,   -43,    26,   -15,   -94,   -23,    -8,    -2,    23,   -10,    20,    39,    65,    64,    -7,    28,     2,   -20,   -12,    -1,   -25,    18,   -43,   -45,   -12,    25,    28,    19,    12,   -18,    26,   -15,  -130,   -57,     7,   -12,    27,   -23,    12,    30,    81,    49,   -46,   -24,   -51,    -5,   -35,   -15,   -37,   -30,   -16,   -44,   -48,   -16,    52,     6,    16,    30,    58,    66,  -133,    24,   -27,     7,     3,    12,    86,    80,    68,    11,    27,   -60,     3,     6,   -49,   -79,   -13,     7,   -21,   -48,   -36,    41,    64,    11,   -26,    30,     7,    44,  -150,   -63,   -34,     1,    14,   -17,    42,    53,    14,   -18,    10,   -23,   -15,   -36,   -36,     1,     0,   -48,   -31,    14,    14,    30,    59,    -9,     6,   -30,   -23,   -31,  -120,   -36,   -18,   -20,    13,    -6,    27,    68,    47,     0,    -3,   -19,   -47,    -1,   -16,   -38,    38,     0,    37,    -3,    25,    61,   -31,    19,   -24,   -16,   -75,   -22,  -119,    -7,   -31,    -7,   -19,    20,    14,    26,    45,   -24,   -33,   -42,   -73,   -37,   -42,    -9,    12,    45,    40,     3,    38,    32,   -16,    19,    -9,   -19,   -28,    18,   -60,   -48,   -36,    -5,    17,   -49,    11,    25,    31,     0,   -13,   -43,    -2,   -35,   -31,   -15,     1,    40,    27,    77,    53,   -10,   -14,    33,    27,    32,    35,    -5,   -84,   -37,    -3,   -10,   -11,    20,    -5,     9,   -43,    32,    56,    -1,   -16,   -28,     0,    17,    37,    57,    62,    42,    19,    27,    56,    -5,    29,    46,   -14,   -67,   -82,   -44,    -8,   -10,     0,    43,    32,   -45,    26,    56,    65,   -12,    11,    32,    16,   -21,    13,    36,    19,   -28,    22,   -14,    43,     6,    38,    86,    18,   -51,   -57,   -34,    -8,     7,     8,    19,     5,   -25,   -13,    24,    57,    21,    17,    11,    29,    -3,   -19,   -16,    27,    21,    -6,   -21,   -37,     3,    87,    83,    40,    72,    29,   -45,     8,     3,     2,    48,    81,    71,    -1,    55,    50,    36,    62,    21,   -19,   -17,     8,    21,   -18,    -3,     7,   -36,    19,   112,    71,    40,    46,   -73,   -43,   -14,    -3,     8,     0,    12,   -24,     1,    67,    53,   -10,    22,    24,   -31,   -13,    23,    69,     5,   -10,   -10,    13,    31,    36,   -31,   -86,   -99,   -97,   -76,   -23,   -16,    -9,    -1,     7,    -1,   -12,   -97,    44,    22,     6,    29,   -23,   -18,   -44,   -44,   -25,   -34,     2,    87,    93,    86,    16,   -19,   -37,  -104,   -50,    -5,    -6,     3,     8,    -1,    -7,     7,     4,   -16,   -30,   -28,   -13,   -22,   -62,   -54,   -45,   -36,   -59,   -52,   -33,    -4,   -13,    -5,   -45,   -56,   -17,   -18,   -12,     8,     6,     6,     4),
		    84 => (    1,    -2,     9,     6,     5,     1,     4,     3,     8,     0,     1,     0,   -33,   -18,   -12,   -17,     0,     3,     5,    -7,     6,     1,     4,    -2,    -3,     6,    -1,    -6,     5,    -7,     3,    -4,    -6,   -20,   -32,   -44,   -25,   -42,   -38,   -37,   -46,   -51,   -11,   -46,   -42,    -8,   -24,   -23,   -43,   -28,   -18,   -38,     1,     4,     6,    -8,     8,     5,   -21,   -36,   -50,   -61,   -54,   -56,   -91,   -78,  -111,  -120,    11,    24,    -3,   -60,   -55,   -70,  -104,   -57,  -117,   -54,   -56,   -37,   -20,   -26,     9,     5,     7,    -2,    -6,  -107,   -69,   -75,   -43,   -64,   -50,   -97,   -85,   -89,   -54,  -119,   -14,    -8,   -59,   -35,   -33,    -6,    42,    -1,   -54,   -63,   -35,   -23,   -11,     0,     4,    10,   -46,  -103,   -10,    -1,    21,     2,   -50,     3,   -14,   -72,    -7,   -15,   -34,   -45,   -21,    -5,   -13,     6,    -1,   -32,    12,    17,    24,   -18,   -69,   -11,   -10,    -9,   -53,    -7,     3,   -14,    -5,   -12,    26,   -15,    38,     1,    43,   -34,   -20,   -49,   -33,    27,    -9,     6,   -45,   -19,     8,    -5,   -24,    25,   -28,    -3,    -4,     6,   -28,   -43,    21,    53,    34,   -47,   -16,   -53,    -6,    16,    -3,   -34,   -79,   -83,   -64,   -47,   -66,   -37,   -82,    -3,    -6,    -6,   -19,    -8,    -1,   -35,     8,   -95,   -35,     1,    23,    40,   -40,   -50,   -73,   -34,   -16,    -6,   -54,   -43,   -58,   -73,   -62,   -19,   -36,   -46,   -41,   -30,   -33,   -24,    12,    48,    43,   -60,   -32,   -81,    55,    15,    42,    17,   -70,   -75,   -82,   -35,   -70,   -47,   -34,    -9,   -98,   -56,   -56,   -14,   -23,   -12,   -39,   -45,   -30,    -8,    38,    43,     0,   -20,    -1,   -65,    46,    12,   -36,    -2,   -50,   -32,   -42,   -43,   -65,   -18,     1,   -25,   -57,   -22,   -34,   -14,     3,    25,    19,    46,    24,    31,    49,   -36,   -61,   -20,    10,   -40,    32,     8,   -27,    30,   -20,   -49,   -24,    -5,    -3,     2,    37,   -14,   -27,    39,    32,    64,   -15,     3,    27,    19,    16,    -5,    -7,    10,   -32,   -13,    -6,   -48,    -7,     1,     2,    58,     0,     4,    18,    63,    49,    30,    61,   -17,     6,    41,    64,    13,   -26,   -12,    -1,    10,    28,    26,   -10,   -13,   -68,   -60,    -2,    -4,    29,    32,   -10,    43,    35,    26,    38,    48,    46,    44,    55,    23,   -18,    -5,     6,   -10,   -33,    -6,   -11,    25,    45,    25,    69,    40,    33,   -69,     7,   -11,    -5,    57,    26,    51,    20,    37,     2,    26,    29,    73,    65,    38,     1,   -20,    32,    22,   -40,     8,    10,    47,    34,    44,    35,    92,    84,   -41,     7,    13,   -89,    25,    83,    59,    29,    24,    50,    35,    28,    23,    45,    -1,   -14,   -26,    36,    61,   -33,    51,   -23,    59,    29,   -25,    -2,    53,    53,   -10,    -5,    15,    89,    42,    -2,    48,    17,   -21,    11,    23,    30,    23,    14,    10,   -11,    35,    54,    10,    -2,    45,    -6,    -3,    54,    31,   -22,    36,   102,   -14,     1,     5,   -20,    57,    19,    43,    56,    42,    30,    12,    -5,   -15,    19,     1,   -12,    62,    21,    28,    58,    77,    22,    11,    -1,     2,    -6,    31,    64,   -24,    -7,   -15,    25,   -22,    71,    52,    23,    33,     4,     9,     3,    -2,     4,    21,    19,    19,    30,     9,     5,    36,   -28,     0,    13,    14,    14,     9,    41,    -3,   -55,     1,    53,    23,    55,    -1,   -12,   -13,    18,    36,     3,    27,     9,    41,    45,     6,     7,    12,    23,   -20,   -16,     3,   -10,   -30,   -16,   -59,   -18,   -21,     3,   -38,   -28,    73,    -4,    56,     9,   -47,    24,     7,   -28,     7,     3,   -17,    35,     4,   -21,   -25,   -33,   -62,   -44,   -37,   -66,   -72,   -19,   -44,   -22,   -20,    -3,   -10,   -51,    49,    28,    -1,     5,     2,    11,   -41,   -93,   -52,   -68,   -32,   -14,   -41,   -20,   -51,   -62,   -52,   -93,   -70,   -52,   -65,   -22,  -103,   -18,     0,    -3,   -16,   -79,    24,    32,    12,   -44,   -73,   -24,   -43,   -64,   -38,   -54,   -40,   -64,   -29,    -2,   -25,   -40,   -65,   -23,   -54,   -28,   -44,    12,   -61,   -67,    -4,   -11,     1,     0,   -59,   -92,   -16,     0,   -72,   -79,   -70,   -13,   -21,   -49,   -55,   -31,   -18,   -37,   -45,   -36,   -15,   -49,    11,     7,    30,   -31,   -23,   -11,   -18,    -7,    -3,    -3,   -79,   -37,   -93,     0,    25,     6,   -56,    27,   -27,   -20,   -24,   -30,   -20,   -25,     3,   -29,   -10,   -29,    12,   -19,   -50,   -67,     6,    -4,     8,    -3,     3,     0,   -10,   -73,    -6,    21,    31,    28,    19,   -36,   -12,   -65,    22,    33,   -32,    -2,   -36,   -80,   -51,    -9,    23,   -12,   -39,  -114,   -18,   -28,     4,     2,    -7,   -22,   -13,    15,   -55,    13,     1,   -24,   -52,   -19,   -21,   -68,   -56,   -26,   -84,   -13,   -29,   -40,   -64,   -18,    -4,    27,   -10,   -72,   -34,   -24,    -3,     4,     7,    -1,   -60,   -28,   -16,   -61,   -69,   -30,   -33,  -100,   -71,   -50,  -104,   -93,   -67,   -91,   -36,   -22,   -99,  -136,  -130,  -116,   -32,   -30,    -9,    -7,    -6,     8,     1,     7,    -7,    -5,   -13,   -11,   -14,   -22,   -24,   -79,   -87,   -47,   -64,   -82,   -27,   -43,   -89,   -55,   -63,   -77,   -57,   -52,   -14,     6,    -6,     4,    -8),
		    85 => (    3,    -2,     8,   -10,     0,     1,     2,   -10,    -2,    -8,    -9,    -7,    -6,   -14,    -2,     6,     5,    -6,     4,     0,    -6,    -9,     1,     4,    10,    -2,    -7,    -7,    -5,     9,    -2,    -6,   -10,    -5,    -9,     8,     3,     7,   -16,   -37,   -35,   -41,   -31,   -29,   -42,   -39,   -49,   -61,   -34,   -32,   -15,    -7,   -10,     3,    -4,    -2,     2,     9,   -18,   -18,   -13,   -12,   -27,   -19,   -96,   -75,  -113,   -99,   -78,   -81,   -81,   -14,   -10,    16,    20,   -19,    23,    10,    -9,    22,   -36,   -19,     6,     5,     2,     7,   -30,    33,    47,   -31,  -106,   -85,   -16,     9,    33,   -56,   -67,   -12,   -37,    56,    41,    20,    78,    60,    67,   128,   101,    72,   -30,    32,    24,     1,    -4,    -3,   -36,    36,  -110,   -97,   -54,   -33,  -106,   -29,    34,   -28,   -26,   -49,    14,    49,    47,    79,   147,    68,    74,    88,   154,    71,   -50,    10,   -35,   -27,     3,     8,   -49,    50,  -119,   -39,   -35,   -31,    -1,    35,    44,     6,   -31,   -53,    20,    20,    51,    71,    87,    92,   114,    22,    71,    23,   -29,   -35,   -52,   -57,     3,     4,   -11,  -112,   -17,    57,    57,    24,    49,    23,    22,     0,     1,   -49,    -6,     4,    13,    -3,    64,   102,    63,     1,    55,    47,    76,    75,    12,    15,    -3,   -17,    -8,  -124,   -69,   -27,    27,    11,     6,     0,     1,    45,   -38,   -21,   -24,   -76,   -18,   -26,    45,    79,    26,    36,   119,    99,    90,    22,    40,    71,   -32,   -38,   -53,  -132,   -41,   -47,    20,    32,    -9,    -3,   -43,    19,    30,    -2,   -29,   -57,   -76,   -12,   -24,    74,    53,    55,   101,    87,    57,    10,    31,    45,     6,     0,   -53,   -71,   -34,   -29,   -17,    20,    12,   -29,    11,     6,    -8,    -4,   -45,   -78,   -77,   -58,   -13,    64,     7,    17,    53,    71,    72,    37,     5,    -2,    -5,   -12,   -36,  -112,    22,    -2,   -46,   -50,     2,    27,   -45,    36,    32,   -28,   -45,   -34,   -88,   -71,    22,    10,    12,    55,    50,    79,    93,    17,   -26,   -28,    -5,    -9,     2,   -80,    18,   -38,     3,   -38,    12,   -15,   -22,    -3,    11,   -24,   -60,   -32,    34,    18,    -2,     9,   -43,   -15,    39,    67,    85,    57,   -30,   -22,     3,    -1,   -15,   -59,    70,   -12,   -14,    30,    25,    38,    77,     6,    57,   -16,   -15,   -49,   -11,   -22,   -12,   -46,   -50,   -40,     2,    17,    23,    67,   100,   -33,     8,    -6,    -7,   -71,     7,    11,   -14,    48,     1,    -2,    25,    34,    44,   -15,   -36,   -10,   -16,   -38,   -57,    15,   -17,    38,   -43,   -63,   -65,   -43,    71,   -31,     2,     3,   -23,   -76,    42,    21,    63,    -8,     0,    38,    37,    34,   -20,     6,    13,    -6,    -3,   -25,    12,    -4,    38,   -11,    30,    -1,   -13,   -77,   -78,   -32,    17,    -3,   -47,   -14,    54,    74,     6,    33,   -14,    17,    31,    -9,   -13,     4,   -14,   -74,   -25,    10,   -13,   -11,   -20,   -11,     6,    23,    18,   -34,   -61,   -18,    -1,   -11,   -54,   -18,    20,    66,    85,    30,    10,    14,   -22,   -27,   -40,     2,   -19,   -40,   -64,     4,    39,     9,   -29,    31,    47,    -5,   -49,   -99,   -88,   -25,     3,   -15,   -68,   -13,    46,    86,    32,   106,    58,     2,    -7,   -18,   -76,   -14,    13,   -39,   -21,   -32,    11,     9,    34,     8,    39,     2,   -32,  -101,  -152,   -93,   -19,   -11,   -70,    -3,    12,    25,    91,    74,    68,    31,   -48,   -17,   -66,   -73,    25,    13,   -15,   -52,   -18,   -16,    40,   -10,    -7,     6,   -44,  -100,   -86,   -76,     8,   -25,    38,    56,     5,    52,    81,    37,     1,    10,    11,    13,   -32,   -53,    13,    33,    16,    14,   -23,    -1,   -40,    22,    -4,    29,    35,   -19,  -101,   -58,    -4,   -18,    65,    48,    59,   111,    46,     3,    21,    48,     8,    23,   -19,    20,     4,    53,    14,    13,    12,    14,   -19,    -1,    -3,    35,   -43,    19,  -124,     5,    -3,   -12,   -55,    -7,    36,    70,   108,    24,   -21,     7,   -17,   -27,    10,     5,   -10,   -27,    -2,    -2,    20,    -6,     9,    21,    19,     7,   -27,    18,    15,     0,     4,    -5,   -99,   -52,   -10,    10,   -12,    45,     2,    15,    -9,    25,   -18,   -20,    39,    21,    24,    42,    -9,    45,    22,    -9,   -33,     8,    10,    33,    75,    -5,    -4,    -4,    30,   -14,    13,     3,    25,    17,   -18,   -14,    55,    26,    32,    49,    33,    32,    24,    15,   -84,   -30,     9,   -19,   -45,    -8,    47,    40,    90,    -9,    -2,   -10,   -54,   -35,   -68,    -8,     1,    -1,    33,    42,    14,    19,    35,    52,    46,    33,    48,    19,    22,     2,   -17,   -14,   -20,   -56,    15,   -92,   -41,    -5,    -3,    -8,   -12,    46,   -99,   -94,    -2,   -19,     5,   -19,    -6,    -8,    -2,    17,   -33,    50,    56,    48,    16,    53,    49,    49,    92,    82,    62,   -24,    -4,   -10,    -3,    10,     4,   -34,   -56,   -70,   -90,  -124,   -60,   -24,   -16,    25,    51,   124,    65,    88,    24,     6,   -26,    23,     3,     4,    -1,   -68,   -26,    -3,    -1,     3,    -7,    -7,   -10,    -3,     9,    16,   -12,   -14,   -21,   -18,     6,    -2,    11,    -9,  -100,   -48,   -15,   -10,   -30,   -25,   -63,   -81,   -57,   -46,   -10,     6,    -6,    10),
		    86 => (    1,     2,   -10,     7,     9,     0,     4,    -6,     0,     1,     6,     6,    34,    25,    -6,    -1,     3,    -4,    -6,     1,     4,    -5,     1,    -7,     6,    -5,    -9,     0,    -9,    -4,    -7,   -10,     3,     1,    30,    38,    34,    39,    41,    15,    47,    33,   -52,     3,    -7,    30,    25,    37,    49,    16,    11,    -5,    -9,     7,     3,    -4,    -2,    -9,    17,    -5,    23,     7,    37,    26,    42,    54,    31,    23,    45,    25,    18,     3,    31,    31,    46,    52,    85,    72,    53,    24,     9,    26,   -10,    -9,    -9,    -5,   -33,    -5,     8,    36,    67,    77,    70,    70,    82,    65,    39,    59,    41,   -14,     6,    53,    49,    -1,    18,    66,    76,    70,    51,   -18,    -3,    -4,     1,     7,   -69,   -33,    30,    68,    84,    57,    20,    49,    76,    41,    58,    -7,    17,   -25,    30,    41,    11,    26,    61,   -26,     2,    33,    30,    33,   -11,    22,    -5,    -2,   -44,   -40,    36,    45,    33,    42,    51,    59,    69,    23,    36,    -4,    10,    -3,    38,    19,   -36,   -27,     7,   -17,    31,    35,    37,    61,    22,    14,    -6,     2,     0,   -15,    38,    11,    50,    18,     9,    58,    76,    21,   -21,   -23,   -22,   -15,     7,   -13,    18,    12,    12,    50,    16,    25,    26,    24,    -5,   -18,     2,     6,    -4,   -30,    18,    19,     7,    56,    38,    67,    32,     7,    -1,   -29,    -5,   -26,     0,    16,    63,    13,    43,    18,   -13,   -32,    19,    -5,   -25,   -46,    -4,    -5,   -31,   -46,    45,    16,   -14,    18,    31,    32,    31,     0,    15,   -29,    16,   -20,   -36,    63,   -31,    18,    34,    63,   -49,   -62,   -66,   -92,   -58,   -78,     4,    -8,   -47,   -51,    17,    -8,   -19,     5,    24,    -3,     2,    20,    12,   -11,    -1,   -25,   -41,   -67,   -42,    25,    29,   -19,   -59,   -49,   -16,   -79,   -29,   -69,     3,     2,   -38,   -59,    12,   -27,   -25,   -24,   -17,     6,     8,   -25,    18,     5,     8,   -49,   -60,   -69,   -40,    23,     0,   -33,   -67,   -64,   -66,   -22,   -32,   -99,    -1,    -3,   -36,   -76,    -7,    -5,    -2,   -37,   -61,   -25,   -11,    18,    25,   -15,   -39,   -32,   -24,   -21,    23,    24,    -1,   -27,   -46,   -28,   -39,   -23,   -74,   -28,    -4,     1,    -8,   -49,   -12,     7,   -17,   -43,   -96,    -7,    -4,     9,    -1,   -12,   -20,    -2,    27,    75,    62,    17,   -23,    13,   -35,    57,    20,   -26,   -75,   -27,    -4,     0,   -12,   -49,   -10,   -25,   -30,   -94,  -118,   -43,   -14,   -10,   -23,    12,   -23,    12,    40,   -20,    -9,    21,   -21,    19,    -3,    75,   -36,   -42,   -62,    -5,    -9,     1,   -10,   -54,   -48,   -21,   -61,   -57,   -73,   -40,    -5,     0,    -2,   -10,     2,    20,     6,   -25,   -46,   -25,   -26,    -1,    25,    54,    -7,    -8,    -9,     1,     7,    -9,   -16,   -50,   -71,   -42,   -41,   -16,  -106,   -90,   -38,     1,   -10,   -17,   -27,    24,    17,   -40,   -34,    10,   -13,     3,     8,    -3,     0,    23,   -52,   -78,     8,   -10,   -25,   -91,   -15,    24,   -39,   -10,   -77,   -37,   -17,    -7,   -26,   -48,   -24,     4,    14,    -2,    14,    -7,   -10,    11,     7,     7,    18,    15,   -51,   -69,    -1,     0,   -23,   -78,    16,   -25,    -2,    13,    -7,     8,    19,    32,   -26,   -59,   -36,   -18,     9,    -8,    23,     5,    -7,   -19,    -3,    40,    48,    34,   -36,   -88,     2,    -8,   -15,   -98,   -14,   -31,   -10,     7,     9,    44,    63,    53,    30,   -16,    -9,    14,    15,    41,    42,    16,    33,    32,   -15,    24,    35,    52,   -37,   -41,     7,   -27,   -81,   -74,     0,   -24,    30,    38,    46,     8,    90,    81,    60,    14,    26,    -2,    -1,   -12,    -6,    17,    17,     2,    -5,    -9,     4,     0,   -28,   -17,     6,   -23,   -22,   -59,   -22,   -28,   -31,    78,    65,    67,   104,    84,    85,    46,    65,    67,    -4,   -36,    -9,   -43,     9,    -5,   -17,   -24,   -58,   -12,   -61,    -2,    10,    -1,   -55,   -27,   -29,   -54,   -31,    50,   147,    88,    69,    33,    49,    48,    58,    15,   -12,   -18,   -20,    31,    19,    -9,   -12,   -15,   -93,   -76,   -53,   -10,    -7,    -7,   -13,   -36,   -61,   -89,   -63,     6,    40,    68,    51,    42,    31,     5,     7,    -9,   -32,   -23,   -21,    -1,    25,    23,   -10,   -31,  -121,   -71,   -43,    -3,    10,     0,    -3,   -51,   -33,   -45,   -49,   -49,   -52,    -3,    -5,    -9,     2,    -9,    -9,    20,    19,   -52,   -17,    48,    31,   -15,   -51,   -82,   -97,   -33,   -35,   -10,    -2,     7,     4,     1,   -24,   -20,   -10,   -54,   -99,  -100,   -99,  -126,   -64,   -87,   -59,     1,    50,    65,    44,   -36,   -21,   -82,   -45,   -46,   -28,   -11,     4,     7,     6,     5,    -4,     6,   -10,   -30,   -41,   -70,   -50,   -37,   -43,     1,    32,    13,   -26,   -35,   -41,   -37,   -37,   -16,   -72,   -37,   -43,   -59,   -18,     2,    10,    -4,   -10,    -5,    -3,     0,   -18,   -24,    -4,     3,     0,     6,   -17,   -24,    -6,    10,   -14,   -18,    -1,     8,    -3,    -1,   -23,   -11,   -13,   -17,    -7,    -2,    -7,     1,    -4,    -6,    -1,     8,    -6,    -5,     4,     3,    -7,    -2,    -9,    11,    -6,     2,     1,     1,    -3,     7,   -12,    -2,    -7,   -12,    -4,     7,     6,    -6,    -5,     5),
		    87 => (    5,    -4,     6,     2,     5,    -5,    -8,     1,     7,    -8,     6,     2,     8,     1,    -2,     2,     7,     7,    -5,     5,     4,     4,     2,     6,    10,    -6,     3,    -9,     7,     0,    -4,     7,     1,     3,    -8,    -7,     4,    -1,    -1,   -22,   -34,   -25,    -2,   -43,   -81,   -71,    -3,    -5,    -3,     6,    -2,   -11,     2,     8,    -7,    -4,     0,    -6,     5,     4,   -13,    -2,     5,    -7,    -9,   -14,   -49,   -87,   -13,   -10,    -1,   -63,   -23,   -29,   -23,   -13,    -1,    -7,    -3,    -3,    -2,     6,     7,     8,     4,    -1,     7,   -15,   -10,   -19,   -43,   -76,   -55,   -48,   -27,   -37,   -56,   -47,   -34,   -45,   -46,   -35,   -25,   -56,   -19,   -21,   -28,    -5,    -4,   -11,     2,     6,     6,     7,     1,     4,   -55,   -36,   -24,   -96,   -95,   -84,  -171,   -63,   -32,    -6,   -12,   -27,   -76,   -58,   -56,   -59,   -61,    51,     4,   -52,   -64,   -34,   -13,    -6,     8,    -9,     5,   -80,   -33,    75,    10,    47,    24,    36,   -34,   -90,   -99,    -2,   -37,   -62,   -33,   -61,   -77,   -40,   -31,   -24,   -37,   -91,   -38,   -56,    -5,     1,     8,    -4,    41,    56,    46,    73,    50,    52,    30,    37,    81,    -7,     6,   -50,   -47,   -53,   -25,   -11,   -41,     3,    -4,     2,    26,   -75,   -14,   -52,   -26,   -20,    -1,    14,    56,     1,    88,    81,    96,   115,    17,   102,    94,    42,    38,    25,    15,   -17,   -29,    -3,    14,     4,    11,    -3,    85,    19,   -14,   -55,   -14,   -28,   -34,   -13,     2,     9,    10,    38,    17,    76,    15,    50,    49,    41,    67,    15,    27,    25,     3,    -8,   -15,     8,    -6,    -7,    65,    -1,   -45,   -80,   -49,   -37,    -9,     2,    72,    33,    27,     5,     2,    26,    25,     3,     4,    16,    76,    42,    64,    30,     8,     2,   -11,     3,    18,     1,    40,    19,   -81,    11,    61,   120,    -6,   -33,    29,    -9,   -31,   -23,   -17,   -28,    18,     2,   -17,   -40,   -40,     6,   -11,    -6,     6,    37,    27,   -18,    22,   -31,   -25,   -25,   -30,    44,    60,   112,     7,   -21,    23,   -25,   -31,   -56,   -30,   -24,   -27,   -15,   -63,   -14,   -57,   -81,   -25,    -4,   -13,    -9,   -34,   -19,     8,   -47,     3,    18,   -61,   -79,   -58,    15,     2,    22,   -36,   -44,   -34,   -62,   -59,   -67,   -80,  -104,  -122,   -49,   -64,   -47,   -34,    17,    21,    -2,    11,    13,     9,   -14,   -33,   -39,  -140,   -18,   -69,    12,     2,     0,    19,   -53,   -96,   -37,   -34,   -51,   -57,   -44,   -56,   -42,   -21,   -41,   -17,    48,   -13,    19,    21,    -2,   -58,    33,   -26,    -5,   -71,   -44,   -56,   -30,   -12,     8,    -9,   -19,   -29,   -20,     0,     0,   -33,   -28,    17,     8,    24,    15,    26,    20,   -33,    52,    25,    48,    -5,    33,    -6,    22,     6,   -47,   -40,    -5,     6,    -5,   -10,     1,    -9,     1,    -3,   -15,   -47,    -8,   -29,   -16,    -2,    14,     6,    14,   -36,    30,    38,     2,   -50,    64,    -1,    28,    -9,   -43,   -13,   -35,    10,   -15,    -2,   -32,   -10,   -10,   -19,   -10,   -23,     1,    30,   -16,    22,    39,     0,    -8,    -7,    -7,    17,     6,    19,     6,   -17,   -34,    10,   -95,   -71,   -11,    -2,     9,   -58,   -55,   -61,   -40,    33,    38,     7,    40,    46,    14,    24,     1,    -1,   -14,    21,   -12,   -46,   -20,    18,     3,     8,   -10,     6,   -39,    17,   -44,    10,     4,    -8,   -32,   -42,    -6,   -31,    41,     6,     7,     9,    -4,     0,    -6,   -25,   -30,   -37,   -17,   -44,   -21,    -8,   -51,   -17,   -15,   -24,   -46,    36,   -42,    -2,     8,   -10,    -7,   -38,   -63,   -18,     7,     7,    -8,   -38,     8,    -7,    11,     6,   -20,   -45,   -30,   -81,   -45,   -56,   -85,   -36,   -10,    51,   -10,   -53,   -23,    -9,    37,   -12,   -31,  -102,   -87,   -45,    -1,    11,   -10,   -36,    14,    -9,     2,   -13,   -34,   -21,   -89,  -102,   -65,   -60,   -66,   -87,     5,     9,   -68,   -57,    -8,    -7,    -9,   -23,   -68,   -40,   -46,   -53,   -89,   -66,   -54,   -22,   -24,     3,     7,   -24,   -27,   -34,   -64,   -79,   -58,   -71,   -50,   -70,     1,    -9,   -31,   -12,     4,   -14,    -7,   -15,   -89,     5,   -19,   -28,   -14,   -72,   -59,   -13,    -9,   -10,   -24,   -43,     4,   -13,     4,   -34,   -26,   -49,  -145,  -116,   -77,   -41,   -10,   -57,    -9,    -7,    -4,   -31,  -109,   -13,    -4,    15,    22,   -73,   -29,    -1,    -7,     6,    -2,    -2,     6,   -21,    -8,   -68,   -23,   -44,   -59,  -108,   -47,   -44,   -23,   -56,     6,    -1,     2,    21,   -10,    30,    31,   -12,   -17,   -13,   -29,   -51,     0,   -11,     6,    -5,   -17,   -35,    40,   -46,   -19,    18,    23,   -60,   -46,   -40,   -15,   -12,     2,     5,     6,   -29,    28,   -26,   -35,   -29,    68,    31,   -21,   -44,   -29,   -20,   -12,    -7,   -42,     1,    -4,   -15,     3,   -31,   -14,   -17,   -17,   -59,   -12,   -20,    10,     7,     7,    -9,   -36,  -128,   -96,  -111,   -31,    -3,   -26,   -39,   -66,   -47,   -17,     4,    53,     0,   -26,    -2,   -54,     7,    -9,   -20,   -37,    -7,     3,     1,     6,    -7,     7,     7,     1,     4,     9,    -1,   -22,    16,    50,    63,    43,   -13,   -25,   -35,    41,    48,    67,    57,   -13,    -7,    -6,   -27,     2,    -4,    -7,     1,    -8),
		    88 => (   -4,    -4,     3,    -4,    -7,     2,   -10,     9,    -5,    -3,     9,     7,     7,     6,     5,     6,    -7,     3,     6,     4,    -8,     9,    -4,    -1,     7,     9,    -1,    -3,    -5,    -3,   -10,    -3,    -5,    -1,    -8,     2,    -7,    -9,    -8,   -17,   -27,   -25,   -41,  -101,  -109,   -90,   -18,   -16,   -19,   -12,   -18,    -4,     3,     5,   -10,    -8,     1,     9,    -2,    -1,     2,     0,   -19,    -6,   -40,   -38,   -53,   -62,   -41,   -22,    -3,   -51,   -66,    21,    30,    -2,   -42,   -61,   -66,    -7,   -12,   -16,    -6,    -2,     2,     5,    -8,   -22,   -19,   -81,   -67,   -85,   -55,   -30,    20,    27,    34,     7,   -10,   -49,   -71,   -98,   -46,   -16,    16,    39,     4,    22,    24,   -25,   -11,     7,    -8,     5,    13,    -4,   -42,   -88,   -62,   -63,    34,    19,    71,    70,    12,   -67,    -2,   -32,   -30,     9,    -3,   -41,   -33,     9,   -40,    13,    26,    24,    16,   -18,     1,    -6,   -30,   -26,   -80,   -69,   -74,     5,   -25,    23,    52,    42,    12,    34,     7,    39,    42,    55,    23,     1,    -3,   -20,   -60,   -51,    30,    12,   -27,   -37,     7,     9,   -63,   -60,    16,   -54,   -72,   -44,    -6,   -11,    19,    12,   -19,    -3,    26,    40,    37,    14,    23,   -35,   -16,    -1,    23,    19,     7,    28,    -3,   -11,     3,   -60,   -34,    15,    33,   -27,   -42,    -5,    15,    23,     6,    -2,   -14,    -9,     2,    59,    59,    20,    -7,   -24,    20,    20,    46,    58,    23,    13,     7,   -41,   -32,   -42,   -33,    81,    43,     3,    20,    22,   -45,    10,    23,     0,    -9,    10,    12,    28,    26,    16,    18,   -12,   -12,   -26,    -2,    31,   -17,    19,    31,     8,     7,   -29,   -46,    46,    88,     0,     5,   -27,   -18,    10,     7,   -33,   -17,   -21,     5,    25,    -9,   -31,    -8,    12,     3,    -4,   -25,     6,    -8,    59,    84,   -62,   -10,   -29,   -62,   -39,    44,    -5,   -12,    -1,   -35,   -45,   -42,   -48,   -25,    32,    36,   -16,   -73,   -52,   -41,   -31,    -6,   -30,    18,    20,    29,    22,    60,   -52,     9,   -16,   -45,   -22,    31,    -4,    28,   -17,   -26,   -18,   -63,   -31,    -6,    29,     0,   -87,   -81,   -49,   -35,   -11,   -19,   -14,   -19,    48,    16,   -40,    34,   -47,     3,    -6,    -9,    11,   -44,    -4,   -57,   -71,   -40,   -44,   -13,    32,    34,    22,    24,     2,   -31,   -47,   -19,   -25,    11,     4,    22,    -1,   -35,  -105,  -116,   -65,    -7,    -3,     2,   -24,   -53,   -29,   -49,   -41,   -24,    57,    57,    48,    70,    36,     1,    19,    -3,   -23,     8,   -19,    21,    49,    28,     8,   -69,   -93,   -88,     6,   -16,    -8,   -15,   -37,   -49,    -4,    19,   -23,    25,    66,    68,    81,    62,    41,     7,    22,    -6,   -17,     0,    36,    42,    40,   -14,   -42,   -37,     7,   -48,   -22,   -12,    -3,   -24,   -10,   -59,   -10,    49,    49,    54,    86,   100,    52,    43,    58,    22,    10,    14,     3,    29,    28,    37,    18,    19,   -48,   -42,    69,   -78,   -25,    -8,     0,   -30,   -29,   -44,   -29,   -14,    40,    19,    66,    79,    70,    24,    -6,    -6,    -3,    36,    74,    67,    15,    45,    29,     1,    -4,     0,    33,  -101,   -36,    -8,   -12,   -48,   -27,     8,   -48,   -56,     0,     7,     7,    28,     9,   -18,   -31,   -13,    43,     3,    12,    26,    23,     9,   -11,   -13,    16,    21,   -25,   -11,   -45,    -9,   -18,   -50,   -76,   -37,   -51,   -19,   -35,   -30,    -4,   -19,   -38,   -37,   -11,    34,    -8,     0,   -37,     8,   -20,   -63,   -55,   -19,    31,   -15,   -60,    -6,   -18,     4,     4,   -26,   -91,   -45,   -77,   -66,   -68,   -61,   -53,   -32,   -37,     6,    37,    44,    16,    36,   -19,   -19,   -41,   -35,    -4,    24,    10,   -31,   -75,   -44,   -30,    -9,    -1,   -41,   -85,   -48,   -43,   -40,   -10,     3,   -48,   -26,   -27,    32,    40,    67,    45,    22,    11,   -31,     3,    19,    12,     5,    -2,   -68,   -59,   -56,    -4,   -21,   -22,   -52,   -16,   -39,     0,     7,    -7,    -1,    -4,   -27,    46,   109,    45,    33,    61,    40,    35,    -6,     2,    15,   -38,   -24,    -2,   -38,   -30,   -58,    -9,   -20,   -17,   -25,     2,    42,    20,    -8,   -25,   -30,     5,     9,    53,    29,    18,    82,    67,    22,    -9,    -8,   -34,    20,   -25,    18,    27,   -25,   -56,   -55,   -15,    -8,    -4,   -15,    -5,    22,    10,   -23,   -46,   -27,    41,    50,     5,    35,    81,    58,    43,    24,   -31,   -10,    -1,    35,     6,    27,    36,   -79,   -66,   -36,    -1,     1,     6,   -28,   -23,   -16,   -33,   -36,   -50,   -35,     6,    -8,    17,    68,    90,    60,     6,   -15,   -35,    12,    76,    60,    14,   -55,   -28,   -92,   -46,   -22,    -2,    -4,     0,   -28,    -5,  -100,   -69,    -4,   -29,   -64,   -65,    -9,    45,    40,    56,    20,    12,   -62,   -24,     6,    13,   -34,   -91,   -87,   -55,   -48,   -19,   -35,    -7,     7,    -1,     5,   -41,   -35,   -39,   -65,   -48,    51,    31,   -36,   -18,   -12,    22,    -8,   -82,   -40,   -27,   -55,   -56,  -108,   -85,   -44,   -32,   -10,    -2,     3,    -6,     1,    -4,     3,     2,     0,   -16,   -12,    -1,   -53,   -73,   -40,   -12,   -13,   -45,   -86,   -61,   -64,   -53,   -31,   -18,    -7,    -3,   -16,    -6,     8,     8,    -1,    -6),
		    89 => (    1,    -9,     6,     7,    -7,     2,     8,    -5,     4,     0,     2,     2,    -7,     4,     5,    -8,     9,    -9,     0,     2,    -1,     0,     1,     7,     3,     9,     4,    -4,     6,     5,    10,     7,     6,    -3,     1,    -5,    -1,     6,    -2,   -25,   -49,   -32,    -2,    -4,   -14,    -5,   -36,   -29,     3,   -15,   -12,     0,     9,     0,     6,     4,     6,     4,    -7,   -41,   -19,     0,    -3,   -17,   -13,    -2,   -12,   -37,    -2,   -12,   -55,   -23,   -17,   -13,   -21,   -21,   -28,   -14,   -15,    -3,   -12,     0,     0,    -9,    -1,    10,     9,   -23,   -39,   -46,   -39,   -48,   -12,   -19,    -5,   -30,   -27,   -41,   -56,   -47,   -40,   -42,   -66,   -42,   -27,   -26,   -24,    -7,    -7,   -10,     2,     8,    -3,     9,    -6,    -8,   -26,   -10,   -53,     9,   -32,   -16,   -19,   -46,   -77,   -60,   -38,   -34,   -16,   -16,   -37,   -64,   -74,   -36,   -20,   -18,    -5,   -49,    -9,     8,    -5,     3,     5,   -22,     2,    -6,   -13,   -21,   -22,   -31,   -71,   -26,   -27,   -26,    -2,    -8,     5,   -28,   -16,   -34,    -4,   -12,   -40,   -26,    -5,   -19,   -22,    -6,     3,    -1,   -10,   -29,    -1,   -12,   -42,   -40,   -92,   -43,   -32,   -37,   -20,    22,    67,    39,    21,    28,     0,     5,    21,    -1,   -31,   -36,   -19,   -33,   -14,   -20,     3,    -1,   -22,    -1,   -28,   -55,   -71,   -66,   -96,    -5,   -19,    25,    27,    -2,   -19,    29,    -4,    -1,   -20,    -5,    -7,   -11,   -34,   -29,   -54,   -23,    -3,   -16,   -30,   -25,   -11,   -33,   -10,   -61,   -47,   -97,   -33,   -42,    22,    -1,   -26,    -2,    -1,   -82,   -32,    -4,   -10,   -10,     7,   -34,   -25,   -52,   -78,   -21,   -14,     0,     4,    -4,   -15,   -26,   -61,   -73,   -46,   -70,     2,    19,    -5,    25,   -14,   -16,    12,   -40,   -40,   -15,    45,    17,    13,   -40,   -31,   -16,   -31,   -74,    -6,   -32,     8,   -19,   -33,     2,   -10,   -23,   -37,    20,    18,     8,   -46,   -31,   -72,   -56,   -30,   -38,   -69,   -44,    43,     4,   -11,   -56,   -22,     3,   -36,    -8,   -11,   -25,     2,   -67,    -7,    29,    -6,   -27,   -26,    -6,    17,   -14,   -33,   -87,   -52,    -9,   -21,   -34,   -39,     1,   -26,     0,    -4,   -21,   -12,    29,   -44,   -19,    -9,   -29,    -9,   -12,     8,    23,    13,    13,     9,    -6,    35,   -20,   -35,   -73,   -19,   -47,   -76,   -47,   -28,   -21,   -55,    -9,     2,    26,    -3,    10,   -86,   -35,    -9,   -13,    -8,   -42,   -33,    44,    40,    18,     9,     2,   -11,   -59,   -34,   -40,   -67,   -53,   -21,   -13,    17,   -51,   -53,    -8,    -8,    29,     1,   -28,   -61,   -37,   -14,    -6,   -10,   -33,   -48,    -5,    24,    15,    14,    10,    43,   -56,   -26,   -86,   -62,   -40,   -28,    18,     7,   -30,    26,    25,     2,     6,    15,   -68,   -42,   -24,    13,    -7,    -1,    -6,   -43,   -13,     4,     3,    30,    21,    23,   -45,   -20,   -82,   -71,   -67,   -36,   -30,   -34,   -53,    20,    18,    42,    16,     8,  -101,   -72,   -19,     8,    -4,     9,    -4,   -47,   -35,    23,   -29,    46,    -3,     6,   -20,    25,   -18,     1,   -18,   -37,   -50,   -59,   -30,    50,    19,    28,   -22,   -14,   -79,   -33,   -36,    -5,     4,     4,    -5,   -36,   -33,    33,   -34,    -1,    39,   -36,    -1,    -9,    -9,   -12,   -50,   -20,    -3,     3,     0,    19,    14,    21,   -23,   -15,   -46,   -11,   -15,   -31,   -12,     1,     7,   -38,   -20,    34,    28,    24,    -6,   -25,    -7,    51,    20,    32,     7,    16,   -20,   -28,    24,    33,    11,   -19,    12,    22,   -35,   -72,    -1,   -38,   -29,    -6,    -2,   -24,   -14,    15,    66,    50,    79,   -23,     7,    47,    99,    23,   -11,   -30,    -6,    -7,     5,    43,   -30,   -10,   -20,   -10,   -39,   -25,    18,   -40,    -6,     5,   -11,   -15,   -18,    -4,    28,    15,   -10,    10,    18,    -6,    -1,    -6,   -30,   -67,   -31,   -22,    18,    49,   -23,   -16,     4,   -11,   -15,    54,    21,   -38,     0,     5,     7,   -38,   -24,   -56,   -16,     9,    35,    21,     5,    -3,   -11,   -28,   -26,   -23,    -1,     7,    -4,    24,     8,    14,   -37,     1,     4,    65,   -14,   -76,    10,    -6,     6,   -14,   -20,   -34,   -32,   -40,   -41,    -3,    -7,   -26,   -42,   -17,   -48,    29,    11,   -13,   -10,    -2,     6,    13,    -7,    23,   -12,    52,    13,   -59,     2,    -3,    -3,    -9,    12,   -34,   -39,   -35,   -49,   -49,   -85,   -91,   -82,   -68,   -14,    17,    42,   -33,   -14,   -36,    29,     8,    22,    67,    -6,    58,    20,   -36,    -3,     4,     1,   -18,     5,    -4,    -8,   -19,   -12,   -30,   -40,   -78,   -71,   -16,    55,   -12,    -2,    -1,   -19,     9,    24,    39,    47,    64,    44,    48,    18,    -3,     6,    -4,    -7,    34,   -24,   -22,    10,    -8,   -27,   -25,   -39,    -1,    13,    38,    53,    -5,   -32,   -40,   -51,   -14,    62,    76,    49,    78,    36,    30,   -15,   -18,     5,     2,     5,     5,    12,    22,     4,    -1,     7,    -3,    -5,    -3,    -6,   -18,   -38,   -21,   -69,   -87,   -46,    -9,     8,    57,    34,    24,    29,    -5,    -1,     8,    10,    -2,    -6,    -1,     9,   -17,    -5,    -2,     2,     2,     3,     8,     8,    -6,    -3,   -26,   -11,   -34,   -56,   -39,   -39,   -24,   -33,     4,   -13,     4,     0,     1,     5),
		    90 => (   -9,     3,    -6,     4,     4,    -4,    -7,     3,    -1,    -4,     6,     4,     1,     8,     2,    -7,    -6,     8,   -10,     8,     1,    -2,     3,     1,    -8,     8,     3,    -9,    -8,     0,    -5,     9,    -1,     4,    -7,    -5,    -6,     1,    -8,    -8,     9,     8,   -13,    -8,    -1,     5,     2,     6,    -2,     1,   -10,    -1,    10,     3,    -1,    -5,     6,    -8,     1,    10,    -2,     3,   -21,   -11,   -15,   -22,   -21,   -12,   -18,   -26,   -18,    -9,    -4,     6,    -3,   -10,    -4,     0,    -5,   -14,   -11,     4,     1,     0,     0,    -8,     1,     9,   -12,     2,   -12,    -1,     6,    -9,   -13,   -21,   -36,   -16,   -11,   -11,     9,    21,    20,     1,     0,     2,   -10,   -17,    10,     7,    -2,    -1,     8,    -3,     8,   -15,   -13,   -36,   -25,    15,     7,     3,    -4,   -29,   -19,   -19,   -14,   -12,    26,    34,    15,    31,    29,     1,    -6,   -11,    -2,    -9,   -11,     6,    10,     5,    -8,     7,    -3,    -9,     9,   -32,   -12,   -18,   -19,    -9,     4,     6,   -14,   -13,     2,   -13,     3,    40,    39,     4,   -11,   -11,   -10,   -10,    -8,   -28,    10,    -3,   -16,   -15,    -9,   -24,     9,    15,     5,   -19,   -16,    -6,   -12,   -21,   -11,   -18,    21,     8,     2,    17,    28,    19,   -12,   -12,   -15,   -42,    -9,     2,     4,   -12,   -20,   -22,    -4,    12,    32,     6,   -17,    16,    13,     7,    15,     9,     1,    37,    10,    23,    46,    13,     2,    10,    29,    -1,    -7,    -1,   -24,     3,     2,    -8,    22,   -19,    16,    18,    12,    26,    12,   -25,   -17,     6,    23,   -19,    -6,   -16,     2,    17,     7,    15,    36,    32,    19,    20,   -14,   -11,   -21,   -15,    -9,     1,    11,    -4,    46,     7,   -12,    -2,    14,    16,   -13,   -48,   -53,   -41,   -38,   -41,   -19,    -9,    -4,     0,     3,    42,    24,    -9,    12,   -15,    -2,    -7,     6,     5,     5,     1,    -3,    38,    35,    31,    26,     4,   -47,   -39,   -45,   -31,   -22,     3,   -44,   -29,   -29,   -16,   -20,   -23,    30,     7,    -9,   -15,   -22,    -2,     8,    30,     5,   -10,    24,    40,    17,   -22,     5,   -41,   -48,   -66,   -51,     3,    11,    13,   -24,   -28,   -43,   -63,   -52,   -31,     2,     5,    34,     1,    -4,    -5,    -5,    -3,     7,   -10,    28,    19,    11,   -16,    -6,   -34,   -56,   -66,   -42,     2,    -8,   -16,   -62,   -71,   -44,   -46,   -47,   -19,    -2,   -11,    20,    16,    -8,     9,     9,    -6,     3,     5,    46,     7,    41,   -21,   -24,   -50,   -74,   -76,   -37,   -20,    -8,   -25,   -56,   -45,   -55,   -52,   -51,   -25,     4,    22,    22,     7,     1,   -15,     5,    -2,    -3,   -31,    52,    33,   -12,   -39,   -55,   -63,   -55,   -47,   -46,   -37,   -22,   -52,   -46,   -40,   -44,   -47,   -45,   -23,   -31,   -11,   -24,    15,   -15,    -6,    -7,     7,    -2,     5,    46,    21,    -8,   -28,   -36,   -55,   -44,   -47,   -26,   -25,   -26,    -9,   -21,   -39,   -34,   -40,   -44,   -21,     5,    -3,   -16,     4,   -13,     0,     7,     4,   -18,    -3,    26,    36,    25,    -6,   -18,   -26,   -31,   -28,   -34,   -27,    23,   -21,   -20,   -61,   -59,   -57,   -23,   -41,   -10,    40,     1,    16,   -24,    11,     5,    -6,   -18,    22,    40,    30,    32,    32,   -21,   -27,     7,    -2,   -20,   -24,   -17,   -32,   -61,   -60,   -60,   -53,   -34,     2,    24,    -5,    -8,    15,   -55,     9,     4,    -3,    -9,    -5,    59,    18,    17,    30,    -8,    -8,    -2,   -22,   -10,   -18,   -49,   -22,   -48,   -50,   -70,   -41,   -20,    20,     3,    12,     4,    -9,   -12,    -6,     9,     2,     9,    -2,    38,     3,     9,    17,    -8,     3,    11,    -9,     1,   -15,   -16,   -25,   -36,   -14,   -15,    -5,    23,    -1,     3,   -18,     5,   -33,   -17,     4,    -9,     1,     8,     0,    29,   -14,    29,    16,     6,   -25,   -16,     9,   -18,     3,    11,    -3,    20,    24,   -29,    -7,     6,    -6,    16,   -13,    -4,   -25,    -5,     0,     4,     2,   -12,     0,     2,   -32,     3,    39,     3,     3,    -8,    18,   -17,     1,    -5,    -2,   -19,     7,     4,    19,    13,     7,   -22,    -1,   -19,    -2,     9,    11,     9,    -4,    -5,   -16,   -21,   -13,   -28,    30,    11,   -11,     6,    14,   -15,     4,   -10,   -21,    20,    23,    -4,     9,     8,   -17,   -10,   -15,   -24,     2,    11,    12,    10,    -3,    -3,   -19,   -12,   -15,    13,    26,    -9,   -19,    -6,     0,     9,   -22,    -9,    -4,   -23,    -4,   -16,     9,    -2,     1,    -1,   -23,   -33,   -25,   -24,    -5,    -5,    -6,   -10,    -9,   -16,    -8,    36,    27,    19,   -21,    -3,    -6,   -19,    10,    22,    17,     5,    12,    17,   -15,   -18,     1,    -6,   -12,    -1,     1,    -5,     7,    -7,     3,     4,     0,   -11,    -8,    22,    41,    41,    10,     2,    -1,   -17,   -15,   -28,     3,    -1,   -17,   -44,   -59,   -51,   -36,   -33,   -22,    -5,    -7,    -4,    -3,     6,     9,     6,    -1,    -3,   -23,   -34,    -1,   -10,    -1,   -11,    -3,     4,   -22,   -21,   -16,   -26,   -77,   -43,   -42,   -43,   -29,   -12,   -31,    -1,    -8,     6,    -6,     8,     1,    -7,    -1,     4,    -3,    -1,    -4,     2,    -8,     0,    -4,     9,   -14,   -12,    -4,    -3,    -2,     0,   -10,     4,   -20,   -27,   -24,    -1,    -3,     0,   -10),
		    91 => (   -4,    -1,     6,    -4,     6,    -4,    -7,    -3,     6,     3,    -2,     4,     9,    -5,    -3,     9,    10,     7,     9,    -4,    -7,    -3,     5,     7,     4,     7,     9,    -6,    -3,     4,    -1,     5,    -3,    10,    -2,     0,     5,    -2,    -3,    -5,    -4,   -18,    52,    26,    30,   -33,    -9,    -1,    -6,    -5,    -7,     0,    -6,     3,     0,     6,    -5,     9,    -6,     5,     8,    -9,     4,     9,   -32,   -34,   -25,   -28,    -9,    18,    18,    36,    84,    51,    45,    16,    26,   -55,   -41,   -51,    -5,     0,   -10,    -1,    -1,    -6,    63,    31,    -6,   -32,   -58,    35,    10,     9,   -44,   -72,   -32,    -2,    -7,     4,    16,     2,     7,   -44,   -14,   -33,   -28,   -33,   -27,    -5,    -1,    -5,     6,    -3,    61,    57,    50,     3,   -17,    21,    41,    36,    20,     6,   -47,    10,   -16,    18,    -9,    -3,    -4,   -46,   -49,   -23,    45,    36,    32,   -22,   -17,   -25,    -3,    -9,    24,    17,    68,    57,     9,    11,    39,     6,   -10,    -8,   -20,   -22,   -46,   -12,   -12,   -15,   -23,   -17,   -54,    18,    46,    60,    48,   -40,   -22,   -33,    -9,    -7,   -29,     2,    69,    27,    21,    -5,   -42,   -33,   -11,   -15,    19,   -23,   -14,   -33,   -43,   -30,   -22,   -78,   -24,    29,    53,    47,    15,    -3,   -14,   -14,     7,    -3,   -35,   -39,   -35,   -28,   -41,    24,   -76,   -17,    71,    52,    44,   -11,    12,   -28,   -62,   -31,   -15,   -52,   -15,    37,    52,    58,    12,   -28,   -38,   -14,    -9,     1,   -44,   -30,   -36,   -37,   -34,    47,   -63,   -17,    64,    -5,    42,    -2,   -17,   -23,   -30,   -51,   -45,   -46,    25,    28,    27,     9,     9,   -20,   -43,   -17,     1,    -2,   -40,     1,   -30,   -39,   -24,    57,   -20,    10,    28,    -3,   -33,   -42,   -33,   -25,   -44,   -80,   -47,   -66,     8,     4,    25,    20,     6,   -10,   -38,   -20,    -6,    -6,   -28,    -2,   -28,   -19,   -39,    21,    15,   -26,    43,     6,     4,    -2,   -11,   -27,   -65,   -58,   -14,   -16,     0,     4,    25,    37,   -24,    -4,     9,    19,    -9,     5,    -4,     0,     1,   -29,   -55,    24,   -39,   -15,    -4,   -24,   -11,   -26,    28,     2,   -52,   -18,   -13,   -17,   -14,   -27,    34,    19,   -23,     5,     0,    47,   -10,     7,   -29,    -1,     8,   -19,   -23,   -27,   -52,   -43,     3,     0,   -15,   -30,    14,   -16,   -17,   -12,    -8,   -17,   -19,   -30,     2,    12,   -38,    14,    28,    54,     5,    -5,   -22,    -2,   -11,   -22,    -5,    -8,     3,   -12,   -16,   -24,    10,   -22,     2,     5,   -28,   -18,   -45,   -20,   -31,   -40,   -35,   -79,   -39,    36,    10,     8,    -2,     9,    11,    12,   -16,   -33,    10,   -16,   -21,   -34,   -68,   -92,   -32,    28,    20,    21,     2,   -10,   -14,   -62,   -47,   -54,   -61,   -34,   -22,   -43,    -3,     3,     7,     4,    -4,    -3,   -21,   -68,   -34,   -34,   -46,   -70,  -105,   -89,   -31,    18,    38,   -31,   -41,    15,     5,   -50,   -58,   -28,   -57,   -31,   -73,   -63,   -53,   -13,     4,    -8,     0,    -4,   -22,   -15,   -32,   -35,   -47,    -9,   -41,   -28,   -45,   -14,    48,    11,   -22,    14,    10,   -17,   -15,    -6,     0,   -26,    46,   -66,   -50,   -13,    10,    -2,    -5,   -13,    -7,    -7,   -14,   -22,     8,     2,    24,     9,   -34,   -13,    31,    -7,    23,   -21,    17,     8,    32,    28,    25,    -8,     1,   -49,   -35,   -34,     6,   -10,    -6,   -35,   -22,     4,   -41,    -2,    27,    52,    30,   -45,   -54,   -37,    16,     8,     9,    35,     8,    13,   -31,   -12,    15,     2,    12,    -3,   -32,     2,    -9,     1,    21,   -35,   -21,    -6,    58,    65,    81,    75,    59,     9,   -60,    -3,    -9,    26,    41,     5,    13,   -27,    -4,     3,    38,    86,    28,    25,   -33,   -13,     9,     2,    -4,   -19,    21,    40,    59,    68,    44,    40,    33,    -2,   -23,    -7,    21,     0,    25,     3,     6,    12,    53,    49,    60,    34,    20,     2,   -23,    -6,    16,    19,    -9,    -6,   -20,   -43,   -24,    -2,    -6,   -21,   -23,   -46,   -13,     8,   -32,     3,   -40,   -25,     4,    22,    21,    -8,    29,    11,    -3,    31,   -16,    -2,    29,    13,   -26,   -18,   -18,    34,    -6,   -20,   -54,   -46,   -42,   -54,     9,     7,    -3,    17,   -41,   -16,    -7,    -4,     5,    -1,   -45,   -31,   -10,    -1,    10,    -8,    -9,    -8,    -9,   -21,     9,    42,    52,    22,    -5,    -7,    11,     3,    43,    11,   -34,   -33,   -33,    23,   -19,   -15,    38,     5,   -21,   -29,   -26,   -36,    46,     0,    10,     3,     7,   -12,     1,    -1,     0,   -17,   -17,   -18,    10,    10,   -12,     3,   -32,   -68,   -30,   -37,   -22,   -58,    -5,   -53,   -21,   -21,   -47,    31,    42,     5,    -8,    -1,    -1,   -19,   -15,   -23,    -6,   -21,   -28,   -17,   -30,   -10,    -1,    35,    37,   -24,   -54,   -37,   -37,   -39,   -71,   -48,   -22,   -16,     6,     2,    -4,     1,    -6,    -3,     3,   -16,   -16,   -44,   -41,   -29,   -16,   -14,   -10,    -1,   -12,   -30,   -40,   -29,   -25,   -38,    -6,    -8,   -15,   -17,   -10,    -7,     7,     7,     4,     4,     3,    -8,     2,     6,    -8,     3,    -8,     0,    -5,     8,   -17,   -31,     8,    -7,    -9,     3,    -5,     6,    -6,    -8,    -1,     0,    -1,    -2,    -1,     3,     3,    -4),
		    92 => (    7,    10,    10,     7,     3,    -1,    -6,    -7,    -3,    -7,    10,    -9,   -10,   -12,    19,    17,    10,    -6,    -8,    -4,     1,     0,    -8,    -5,     4,     1,    -6,     3,    -6,     6,    -3,     4,    -4,     8,   -10,    12,   -15,   -32,   -45,   -64,   -13,   -18,    -7,    27,    36,     3,   -28,   -79,   -50,   -54,   -37,    -8,    10,    -8,     0,     7,     5,    -7,    -5,   -24,   -26,     2,    10,     4,     5,    66,    64,    74,     6,    21,    56,    91,    76,    33,   -34,   -71,   -38,   -16,   -37,   -11,    -4,     1,     9,     8,    -7,    -2,     4,   -51,   -63,    28,    39,    52,    -1,   -45,   -68,   -89,  -114,     1,   -13,     1,     6,   -35,   -86,   -56,   -49,   -11,     3,   -55,   -60,    -5,   -10,     1,    -5,    -3,   -15,   -42,    -1,    22,    93,    74,    55,    91,    26,   -22,   -32,   -33,   -23,    13,   -27,    -9,    12,   -18,   -14,   -43,     5,   -43,   -72,    -6,   -48,   -15,     3,    -6,   -39,   -23,     0,   -40,   -33,     8,    56,    17,    43,     1,    14,    14,    22,     8,    -4,     8,    24,    31,    16,    50,   -18,   -30,   -63,    20,   -85,   -22,    -4,    -5,     7,     2,    20,   -10,    -8,   -12,    40,    -6,    11,   -42,    10,   -34,     2,    -1,    25,    15,    36,    15,    -4,    18,    -9,   -26,  -107,   -13,   -78,   -19,    -9,    -7,    30,     1,    38,    86,    25,    11,    26,    -8,   -58,   -30,    -4,    13,   -18,    13,    31,   -27,     9,   -13,    10,    49,    42,   -76,    16,    46,   -50,   -34,   -45,    52,    33,    12,    -7,    71,    27,   -16,    22,    16,   -18,    17,    16,     4,    -5,   -41,   -26,   -10,   -35,     9,     4,   -32,     2,    44,   -13,   -28,   -83,   -25,     6,   -35,     9,    39,   -50,     5,     4,   -24,     3,   -21,     0,    25,    30,    26,   -19,     0,   -17,    -7,     0,   -18,    -4,   -14,    41,    -7,   -37,  -110,   -14,   -18,    10,     4,   -21,    21,   -24,    50,    79,    11,    10,   -27,    46,   -17,     3,     4,   -14,     3,   -21,    52,   -28,   -32,    -8,    12,   -22,   -72,   -41,   -33,   -27,   -33,    -4,   -40,     7,     5,   -16,    22,    38,    28,    11,    24,    29,    -9,   -38,   -52,   -12,   -41,    -9,   -31,    -2,    15,    17,    -6,   -52,   -41,    19,    21,   -25,   -47,    -4,   -23,   -76,    -1,   -27,     6,    71,    35,    -1,    48,   -10,   -51,   -29,   -23,   -54,   -41,   -43,   -25,    30,    57,   -20,    47,    42,   -42,    50,    13,    -1,   -12,    -7,   -43,   -27,    -9,   -10,    32,   116,    37,   -18,     5,   -13,    -7,   -14,    12,   -45,   -33,   -41,   -13,    21,    37,    -9,    12,    42,    88,    67,    72,    76,   -11,     6,    -4,   -16,     8,    34,    41,    73,    79,   -43,    27,     7,   -65,   -30,   -43,   -32,   -20,   -16,    -4,    -6,    31,   -58,    26,    75,   132,   109,    56,    49,    23,    -1,   -30,    58,    65,    -3,    17,    36,    31,    47,    10,   -21,   -13,   -16,   -36,   -10,    -1,   -13,   -33,   -11,   -28,    17,    43,    41,    38,    -8,    42,    89,    71,    -4,    -4,    74,    68,   -43,   -33,     8,    70,    31,    71,    31,     6,    28,    -6,   -20,   -16,   -10,   -31,   -20,    15,   -18,   140,   114,    71,    15,    79,    96,    53,     0,   -13,    68,    47,   -14,   -25,    15,   -11,   -12,   -11,     8,     2,     5,    -3,    21,   -12,   -22,    -4,    -8,   -11,    41,   147,    81,    32,    24,    37,    38,    35,    -5,     1,    11,    26,   -17,   -12,     6,   -30,    16,   -18,   -27,     4,    12,    -4,   -46,   -25,   -35,   -47,    -6,    35,   128,   111,    86,    62,    48,    42,   -12,    19,     5,   -39,    15,   -18,    -3,    -4,   -24,     0,    22,    16,    25,    35,   -20,   -24,     8,    29,   -21,   -54,    22,    71,    80,   108,    75,    31,    -2,   -24,    15,    53,   -10,   -23,    67,   -34,   -12,    -3,    -4,     1,    -1,    29,    46,    52,     2,     0,   -39,     6,   -43,   -13,    26,    85,   106,   131,    53,    41,    19,    10,     8,    -8,    -6,    -4,    64,   -25,    41,   -11,    12,     0,    46,    74,    42,     1,    21,    21,   -43,    -1,   -10,   -42,    92,   147,   109,    95,   122,    17,   -19,    12,   -14,    -7,    -1,     1,   -21,   -46,   -15,    18,   -34,    -2,    40,    37,    15,    21,   -28,    -2,   -28,   -17,     5,    32,   124,   124,   113,    87,    84,    35,   -47,    20,    -8,    -5,    -9,     7,     2,   -60,    -4,    19,    31,    12,    16,    70,    32,    19,    13,    11,   -25,   -20,    80,   149,   120,    87,   119,   108,    79,    49,   -41,     3,     3,    -8,     6,    -1,   -50,   -20,   -39,   -69,    29,   -27,    -2,    35,    39,    17,   -62,   -98,   -15,    12,    93,   128,   170,   120,    70,    95,    70,   -19,    23,     7,    23,    -1,     9,    -2,   -20,   -10,   -57,  -109,    39,   -31,   -31,   -42,   -61,   -57,   -76,   -75,    11,    18,    14,    65,   107,    29,     6,    17,   -43,   -40,   -22,     0,    18,    -8,     9,     8,     7,    -9,   -15,   -30,   -69,  -102,   -49,  -113,  -133,  -101,   -92,  -135,  -134,  -106,  -107,  -100,   -81,  -129,   -39,   -23,   -48,     5,     3,     0,     4,     2,     4,     8,    -9,     8,   -16,   -13,   -19,   -16,   -12,   -13,   -50,   -60,   -44,   -52,   -58,   -27,   -30,   -26,   -17,   -21,   -15,   -17,   -21,     3,    -9,     4,     6,     8),
		    93 => (   -2,    -1,    -5,     5,    -6,    -9,     4,     4,     6,    -5,     4,    -3,    -5,   -12,     3,    -5,     6,    -5,    -9,     8,     8,     9,     2,    -6,     5,    -8,    -2,     6,     9,   -10,    -1,    -2,     8,     3,    -2,    -5,     8,   -10,   -10,    -3,    -7,   -11,   -16,   -15,   -20,   -24,    -6,    -2,    -9,     1,     2,   -10,     5,     7,    -9,     4,     0,   -10,     0,    -1,    -4,    -9,    -2,     0,   -41,   -50,    59,    14,   -19,   -38,   -63,   -37,   -38,   -27,   -34,   -22,   -68,   -53,   -64,   -39,    -5,    -1,     4,    -9,    -3,    -2,    -5,    -6,     1,   -16,     9,    26,   -36,   -59,   -78,   -63,   -74,   -94,  -119,   -62,   -49,   -59,   -78,   -53,   -49,   -36,   -20,   -49,   -17,   -13,     4,     2,    -8,     3,     6,     1,    20,    57,    65,   -26,   -16,   -79,   -13,   -19,   -22,   -58,   -94,   -89,   -88,   -80,   -76,   -80,   -60,   -19,   -29,   -24,   -18,   -39,    -1,    10,     8,    -6,     2,    12,    27,    55,     4,   -21,    -8,    24,    48,    37,    36,   -19,   -29,   -17,   -28,   -24,   -58,   -82,   -53,   -48,   -50,   -20,   -12,   -51,   -17,    10,     3,    -2,     4,    35,    19,   -33,    16,    43,     1,    34,   -17,    25,    12,   -26,   -36,   -44,   -58,   -51,   -37,   -72,   -59,   -46,   -48,   -47,   -36,    -5,   -31,     3,    -3,    19,    -6,    31,     7,    -8,    43,    15,    28,    -8,   -10,   -44,    -3,     6,   -14,    25,   -42,   -61,   -85,   -95,   -59,   -56,   -41,   -47,   -34,    -7,   -24,   -11,     7,     7,   -32,    18,     0,    -4,   -14,   -41,   -11,    -9,   -48,     0,    54,    57,    63,    42,   -12,   -83,   -98,  -102,   -77,   -34,   -42,   -48,   -32,   -17,   -18,     6,    -6,   -27,   -26,     5,   -13,    19,   -32,   -22,   -41,   -14,   -20,    39,    51,    56,    67,     5,   -42,  -115,  -106,  -105,   -70,   -39,   -30,   -14,   -24,   -32,   -26,    -8,    -2,   -44,   -18,    53,     6,    28,    -1,   -23,   -38,     2,     5,    25,    41,    34,     9,   -37,   -56,  -118,  -128,  -100,   -81,   -74,   -40,    -2,   -18,   -22,   -12,    -1,    -5,   -65,    -3,    69,    40,     8,   -11,    -2,   -14,    20,    30,    17,    31,    -2,   -33,   -39,   -43,   -56,   -47,   -67,   -51,   -70,   -55,   -20,    -5,   -47,   -29,     0,     3,   -49,   -59,    47,   -15,    -4,   -47,   -31,    24,    17,    52,    43,    38,     8,     6,     5,   -41,   -41,    15,     1,    -4,    28,    54,    37,   -38,   -30,   -19,    -8,     2,   -19,   -45,    53,    32,    10,    -4,   -20,    23,    37,    38,    32,    32,    27,    11,   -23,    -6,    -7,    16,    -4,   -14,    16,    30,    48,    45,   -40,   -26,     2,   -11,    20,    -5,    25,   -45,   -30,   -29,   -21,    11,    35,    18,    -8,    -9,     3,   -24,    -9,    13,   -25,    -5,    43,    -5,     7,     6,    86,    31,   -51,   -19,   -12,    -3,    24,     4,    13,   -50,   -42,   -32,    -5,    22,     5,   -19,   -38,   -32,   -32,    -7,   -34,     4,     4,    -2,    30,    56,    37,    34,    32,     8,   -42,    -7,    -2,     8,     8,    -1,     3,   -51,   -78,   -32,   -52,    11,    44,   -35,   -41,   -40,   -71,   -87,   -27,   -36,   -35,    -1,    16,    47,    49,    47,     4,    -7,   -34,   -32,   -16,     9,     1,   -10,    37,   -16,   -37,   -30,   -62,   -26,   -30,   -74,   -41,   -41,   -44,   -80,   -79,   -41,   -42,   -63,    27,    23,    70,    35,    24,    -6,   -28,   -14,    -6,    -8,    -5,     9,     4,     4,   -22,   -50,   -33,    -1,   -23,   -81,   -34,   -16,   -40,   -34,   -64,   -32,    -4,   -13,     3,    24,    34,    24,     3,    13,   -25,   -15,   -31,     9,     1,   -15,   -21,   -27,   -19,   -22,    19,    -5,   -15,   -36,   -22,     9,    22,     8,   -16,     9,    31,   -14,     0,     7,    18,     9,   -21,    16,    -7,   -42,   -22,    10,     1,   -20,   -41,   -30,   -36,   -48,    -1,    17,    21,   -16,    12,    14,    24,    34,    37,    47,    -3,   -21,   -14,    28,    29,     9,    -5,    22,   -17,   -13,    -8,    -9,    -4,     1,     4,    24,    -8,   -62,   -45,   -26,   -17,   -30,   -26,   -39,   -17,     9,     3,     5,   -17,   -34,    -4,    -1,   -41,   -15,    13,   -21,    -2,   -20,    -5,     3,    -3,     1,    -3,     2,    -9,   -56,   -53,   -54,   -48,   -31,   -42,     0,    -4,   -40,   -14,   -41,   -40,   -16,   -15,   -14,   -17,    -9,    16,   -27,   -21,     4,     7,     7,     4,    14,   -28,    -8,   -13,    -9,    -1,   -23,   -22,   -30,     1,    19,   -14,   -29,   -12,   -32,   -23,   -51,   -21,   -27,   -25,   -20,   -42,   -11,   -18,     0,    -1,     6,     3,    20,   -14,   -28,   -22,    22,    32,    18,     0,     1,    71,    13,   -28,    -8,   -14,   -37,   -52,   -31,   -11,   -34,     4,   -11,   -54,   -26,   -18,     4,     2,     9,     1,     5,   -40,    -3,   -16,     6,    19,     8,    -2,   -16,   -20,   -12,    26,    16,   -18,   -33,   -28,     3,   -10,   -71,   -46,   -43,   -63,    -2,    -3,     4,     8,     2,     8,    -2,   -20,   -19,   -24,   -22,   -26,   -51,   -46,   -18,   -42,   -31,     1,   -54,   -23,     4,     2,   -29,   -25,   -26,   -10,   -46,    -6,     8,     2,    -2,     7,     1,    -4,    -4,    -5,     3,    -6,    -7,    -2,    -7,   -22,   -14,   -24,   -23,   -36,   -25,   -48,    -6,     5,     2,   -36,   -19,   -23,   -13,     7,     1,    -2,     9,     4),
		    94 => (   -4,   -10,     4,    -4,     4,     8,     1,    -3,     4,     6,    10,    -7,   -17,    -6,   -17,   -13,    -3,    -6,    -5,    -9,     6,     4,     0,     8,    -7,     3,    -1,   -10,     8,     9,     0,     6,     2,     0,   -18,   -38,    -8,   -36,   -36,   -40,   -41,   -35,    -9,   -50,   -47,   -25,     2,     0,   -42,   -12,   -17,    -5,   -10,    -3,    -1,     2,     4,    -4,     3,   -52,   -78,   -18,   -39,   -55,   -29,   -40,   -70,  -111,   -74,   -48,   -70,   -30,    -8,   -25,   -49,   -47,   -50,    -8,   -37,   -33,   -49,   -24,   -10,     0,    -3,    -7,    -2,   -58,   -97,   -21,   -71,   -69,   -36,   -54,   -65,   -30,   -39,   -84,   -55,   -39,    28,   -37,   -57,    -1,   -12,     7,    11,    19,   -52,   -35,     5,     9,     8,     5,   -26,   -47,     7,   -28,   -59,     5,     6,   -19,   -59,    -7,    28,   -32,   -29,   -80,   -28,   -44,   -44,    46,    33,    26,    -4,   -30,   -55,    12,   -17,    -2,    -3,     1,   -26,   -54,   -55,   -29,   -40,    -5,    19,    12,    58,   -19,   -16,   -34,   -60,   -77,   -30,    12,    94,    19,     6,    16,   -32,   -34,   -55,    22,   -36,     6,     4,     0,   -10,   -10,   -31,   -29,    -9,     5,   -14,   -11,   -68,   -30,   -33,    -9,   -88,  -141,   -25,     7,    40,    54,    84,    82,   -39,   -24,   -40,   -32,   -10,   -29,    10,   -20,   -39,     0,   -34,    -6,   -12,    51,   -12,   -36,   -54,    11,    37,   -24,  -110,   -98,   -14,    21,    38,    30,    25,    24,   -28,   -30,   -58,   -48,   -18,   -29,   -39,   -45,    37,    -4,   -21,    -1,    18,    27,   -33,   -51,   -40,    20,     3,   -44,   -67,   -51,   -51,    80,    10,    29,     1,   -47,   -49,   -67,   -55,   -23,   -46,   -22,    -2,   -42,    27,   -20,   -27,   -36,     6,    -8,   -23,   -15,   -61,    -5,   -18,   -14,   -41,   -71,    -5,    49,    23,   -13,     2,    38,    12,   -52,   -49,   -14,   -13,   -20,    -1,   -31,    34,    47,    -6,   -33,   -48,     4,     9,   -32,    22,     1,   -15,    -9,   -49,  -100,   -25,    34,     9,   -13,   -25,    33,   -38,   -82,   -73,   -12,    -2,   -18,     6,   -64,   -20,    37,   -43,     0,   -12,   -19,    26,    -2,    19,    30,    14,   -24,   -96,   -74,     5,    37,     4,    -6,   -34,   -71,   -67,   -67,  -106,   -43,   -11,   -45,     7,   -32,    15,    -5,   -37,     0,    44,    14,     2,    -8,    46,    18,    25,   -70,   -74,   -71,     2,     7,    12,   -12,   -43,   -60,   -62,     7,    23,    14,   -29,   -43,     2,   -32,   -11,   -11,   -16,     4,    48,    11,     2,    14,    29,    28,   -14,   -67,   -77,   -61,   -23,    20,    25,   -30,   -47,    11,    37,    33,   -32,   -21,   -49,     8,     5,     2,   -58,   -14,    64,    38,     1,    22,   -14,    51,    62,    46,    -8,   -20,   -21,   -45,    -4,     6,    15,    12,    13,    38,    -4,     8,   -17,   -45,   -39,    -3,     3,    -6,    86,    -3,    51,    15,   -12,   -13,     6,    11,    43,    29,    29,     6,   -32,   -50,   -17,    -6,   -11,    28,    -7,    27,    72,   -21,   -64,   -73,   -29,     8,    -1,    -8,     4,   -48,   -26,   -44,    16,     2,   -22,    -7,   -10,   -69,   -39,   -25,   -41,   -16,   -11,     6,    18,   -16,    38,    12,    -5,   -76,   -20,   -38,   -49,   -22,    -7,     9,    21,   -70,     2,   -10,     2,    25,    31,   -11,    -1,   -10,   -73,   -10,     3,    27,    -8,    15,    21,   -20,     9,    28,   -37,   -26,   -52,    29,    -8,   -31,   -22,     7,    22,   -40,    14,    29,    21,    40,    -1,   -11,   -22,   -28,   -73,   -13,    19,    48,    -7,    19,    11,    19,    42,     6,   -59,   -12,   -49,   -39,   -16,    -6,     5,    -8,   -42,     4,   -12,    10,    46,     1,     8,     9,    -6,   -82,   -81,   -24,   -13,    52,     7,   -32,    37,    23,    25,    38,   -38,   -27,   -47,   -63,    -1,    -8,    -4,     5,   -22,   -11,    10,   -26,     3,    17,    -2,   -32,   -58,   -15,    -8,    -1,     4,     9,     3,    24,    32,    32,    29,    41,   -44,   -13,    -4,   -22,    -4,    -2,    -7,     4,   -51,   -10,     8,   -13,    11,    19,    17,   -46,   -44,   -46,   -10,    -1,    -1,    12,   -22,    29,    21,     8,    30,    37,    32,   -25,    35,    -8,   -30,    -6,     8,     9,    -4,   -52,   -76,    29,    12,   -12,   -51,   -76,  -115,   -54,   -37,     1,    -9,   -16,   -21,   -34,    14,    29,    38,    47,    13,   -15,    -7,    62,    18,    -5,     0,     1,    -5,   -33,   -53,   -41,    -8,   -21,   -10,   -76,  -100,   -53,   -44,   -33,    -8,    -2,    26,   -42,     1,    27,    46,    73,   -42,   -29,     5,    18,    14,    -5,     8,     7,    -6,   -11,   -24,    -7,     0,    -9,   -30,   -48,   -59,   -53,   -29,    -9,   -48,   -27,     4,   -18,     2,   -17,     9,   -11,   -54,    -6,   -45,   -30,   -20,     3,    -5,     8,   -26,    -8,   -28,    -4,   -12,     3,   -21,   -50,   -70,   -27,     2,   -29,   -87,    -3,    12,   -13,   -50,   -91,   -45,   -63,   -77,   -37,   -53,   -38,   -25,     6,     0,    -6,    -1,   -10,   -39,     3,    -6,   -12,   -15,   -47,   -86,    -9,   -28,   -56,   -88,   -55,   -92,   -70,   -69,   -63,   -97,   -72,   -80,   -11,    -8,     7,    -5,     6,     8,    -8,     8,     6,   -10,     5,   -10,   -24,   -16,   -29,   -50,   -42,   -40,   -23,   -37,     6,   -54,   -71,   -47,   -37,   -41,   -27,   -45,   -17,     7,     1,     4,    -7),
		    95 => (   -4,     5,     5,    -2,    -5,     4,     7,     1,     7,     9,    -4,    -7,     6,    -5,    -2,     1,    -3,    -7,     0,     4,    -5,    -9,    -6,     3,    -8,     7,     3,    -8,    10,    -1,    -6,     4,    -4,     9,    -1,     6,    -4,     8,   -10,    -7,    -1,     3,    -8,   -13,   -18,   -24,    -6,    -4,    -4,    -4,     8,     6,    -4,   -10,     1,     7,    -2,    -2,    -6,     7,     7,    -8,   -13,   -21,   -25,   -39,   -35,   -32,   -42,   -27,   -18,    21,    -7,    -7,    -6,    20,    29,    14,    12,    40,   -11,    -7,     0,    -6,     0,     1,   -18,    10,    -4,   -10,   -40,   -56,   -15,     2,    38,    10,    39,    56,    75,    26,   -20,   -41,    57,   -15,   -14,    17,   -21,   -27,   -30,     8,    15,    -4,     6,    -6,   -24,     1,   -30,   -32,    30,    -2,   -54,    44,     1,    34,    37,   -37,   -41,   -15,    12,   -23,    13,    45,   -35,    11,    39,    48,    87,    81,    25,   -22,     5,     8,   -17,     5,     0,     8,   -23,   -45,     6,    61,    58,     3,   -46,   -51,   -34,   -15,    26,     4,    18,     6,    15,    39,    41,    39,    61,    52,    49,   -19,    -4,   -11,   -11,   -13,    23,    15,   -36,   -14,    54,    10,    18,   -51,   -44,    -8,    19,    57,    23,    50,    36,   -15,    14,    29,    55,   -11,    31,    29,    50,     2,     1,    -1,    -2,   -33,    -4,    -7,   -24,    30,    34,    44,    37,    -4,   -51,   -23,    52,    47,    76,    57,    20,    15,    17,    13,   -18,   -35,   -26,    36,    36,    14,    -1,    -7,   -56,   -43,   -48,   -24,    -1,    15,    67,    48,    45,   -33,   -22,   -47,    -9,    14,   -18,     8,    16,   -31,   -12,   -51,   -28,   -29,   -26,   -36,    58,    11,    -5,   -13,   -55,   -52,   -29,   -15,     4,     8,    34,    37,    22,    35,   -70,   -88,  -104,  -125,  -137,  -178,   -98,  -132,  -127,  -120,   -79,   -59,   -57,   -36,    58,    30,     7,    -6,   -18,   -41,   -17,    -7,   -23,     5,    28,    27,    13,   -17,   -66,   -86,  -102,   -74,   -72,  -150,  -163,  -143,  -173,  -165,  -151,   -69,   -39,   -21,    18,    35,    -6,    -4,    -5,    -8,    -5,   -21,    -2,   -10,    21,    14,   -33,   -14,   -22,   -30,    -1,    21,    26,     2,   -41,   -47,   -84,   -94,  -111,   -90,   -70,   -17,     3,    11,    -1,    -4,     1,    30,     3,    28,    34,    12,    46,     7,    37,     6,   -19,   -24,   -25,    18,    20,    17,    19,   -18,     5,    10,   -42,   -25,   -45,   -35,    -3,     4,    -5,     6,     2,    15,    36,    16,   -26,   -23,   -10,    19,     2,    23,   -23,   -27,   -39,   -43,    -3,    -4,    11,     7,     3,     3,     8,    31,   -12,   -22,   -28,   -46,     3,   -17,   -13,     3,    51,    20,    44,     1,   -11,    31,    -1,   -16,   -17,   -44,   -33,     7,    -9,   -34,   -20,   -40,    -5,   -13,    29,    13,    80,   -39,   -53,   -28,     2,    18,   -11,   -65,   -42,   -57,    22,   -46,    -1,   -14,    31,    29,   -18,   -23,   -27,   -34,   -16,   -70,   -38,     2,     9,   -21,    -6,    -8,    68,    -1,   -42,   -45,   -10,    -9,    -6,   -36,   -70,   -55,   -33,   -16,   -26,    10,    23,     0,   -14,   -38,    -8,   -11,   -10,   -30,   -70,   -31,   -14,    10,    15,     9,    -3,   -37,   -76,   -68,    -5,   -15,   -28,    37,     1,   -37,    17,     8,   -29,   -12,     6,     5,    -3,   -26,   -48,   -65,   -31,   -38,   -16,    25,    15,    16,    20,     6,     5,    -7,   -74,   -71,    -6,     2,    31,    51,   -23,    14,   -13,    -2,    -7,   -47,     3,   -17,   -35,   -56,  -103,   -56,   -46,   -45,   -11,     3,     0,    40,   -32,   -35,    -8,    -3,   -80,   -68,     7,     2,    57,    51,    23,     3,   -26,   -55,   -86,   -47,   -27,   -63,   -30,  -104,   -53,   -71,   -59,    13,    17,    30,    44,    21,     7,   -28,    51,     2,   -15,   -48,    -4,    -6,    30,    39,    37,   -11,   -36,   -32,   -27,    -7,   -19,   -19,   -21,    11,   -18,    26,    10,    36,    24,    21,     0,     9,     1,   -12,   -24,    -9,   -53,     6,    -9,    -6,   -16,    19,    35,    -5,     9,     2,   -35,   -63,     2,   -18,   -12,    -2,   -36,    42,    17,    53,    11,   -15,     1,    25,    32,    50,    17,    54,    -9,     2,    -7,     4,   -37,    17,   -14,    16,     1,   -11,   -16,   -33,   -41,   -14,   -19,   -17,   -31,    37,    38,     9,     9,    -7,     8,     3,    12,    84,    18,    82,    76,    -2,     1,    -9,    28,    28,    -2,     5,    -9,   -22,    32,     7,   -19,    -4,   -12,    -3,    10,   -23,   -22,   -21,   -23,   -33,    41,    11,    42,    39,    23,    58,    94,   -10,    -5,    -5,     2,    38,    53,    26,    41,   -23,   -14,    32,   -14,   -37,    -5,    28,    18,    47,   -40,    -7,    -5,     8,     9,    20,   -17,   -56,   -11,   -21,   -10,     3,    -9,     3,     9,    49,   -43,   -25,    61,    33,    56,    65,    45,   -10,    63,    44,    46,    36,   -33,    -1,    35,    54,    49,    39,    75,    45,    32,    -9,     6,     1,    -8,    -9,    -5,    -5,    -9,   -15,   -14,    -9,     2,     5,    -1,    12,     5,    54,    29,     9,   -81,   -36,   -18,    10,   -47,   -30,    11,   -23,   -15,     6,     9,    -5,     4,    -4,     3,     5,     6,    -7,     0,     2,    -9,     9,     3,    -4,    -4,     4,   -20,   -14,    -8,    -1,    -3,   -17,   -39,   -49,   -42,     0,     2,     5,    -4,    -6),
		    96 => (   -5,     6,    -7,     3,    -7,    -3,    -7,    -8,     7,     4,    -6,   -10,    40,    42,   -10,    -1,     8,    -9,     0,     7,     3,     1,     4,     4,     3,     7,     6,    -7,     2,     9,    -1,     3,     6,    20,    20,    39,    59,    37,    30,    19,    57,    87,   -27,    17,    39,    53,    50,    14,    44,    22,    22,    14,     6,     4,     6,    -8,    -2,     5,     3,    -4,    57,    63,    42,    43,    24,    27,    46,    65,   102,    72,    37,    35,    44,    49,    16,     3,    12,   -13,   -11,   -13,    16,    12,     8,     2,    -5,     5,    -8,    80,     2,    10,    70,    84,    45,    30,    49,     9,    23,    77,    51,    30,   -13,   -45,   -32,    -6,    20,   -32,   -14,   -14,    -7,   -13,     0,     8,    -5,     1,   -15,    94,     6,    72,    55,    -1,    -5,    13,    14,    12,    39,     8,    -2,   -26,   -39,   -10,   -18,   -26,   -80,   -44,   -60,   -61,   -60,   -45,    -5,    14,     1,     2,   -13,   -18,    28,    22,    -4,   -25,   -34,     9,    17,     3,    47,     5,   -63,    -4,   -68,   -21,   -24,   -52,   -88,   -90,  -105,   -72,   -41,   -28,    17,    16,     6,   -10,    -8,   -49,    23,   -14,   -30,   -63,   -55,    50,    21,    36,    29,     5,   -23,   -70,   -51,   -57,  -117,  -118,   -79,  -118,  -108,  -101,   -50,   -15,     8,   -35,    -5,     0,    -7,   -60,    27,    13,   -51,   -69,    -4,    -4,    27,    25,    11,     3,   -40,   -78,  -108,  -112,  -139,   -95,   -66,   -18,  -112,  -112,   -81,   -32,    16,   -45,    -6,     3,     5,   -53,    38,     1,   -23,   -20,    34,    23,     6,    -3,   -18,     0,   -98,  -161,  -117,   -66,   -70,     1,     5,    24,   -34,   -59,   -79,   -71,     6,   -51,     0,   -12,     0,   -15,    42,    -9,   -40,   -12,    25,    -8,   -10,    14,     0,  -107,   -70,   -53,   -17,    -5,    -8,    56,    64,    52,    30,    16,    -3,   -60,   -46,   -23,    -5,   -13,    -4,   -18,    19,    18,   -26,    -2,    25,   -28,    12,   -12,   -16,  -120,   -75,     4,    16,    53,    45,    24,    29,    20,   -10,    -7,    19,   -24,   -62,   -72,     6,    10,   -11,   -32,    36,    31,   -40,    13,     8,   -19,   -23,   -29,   -50,  -104,   -53,    -1,    32,    26,    26,    28,    34,    -2,    -1,   -12,     8,     5,   -29,   -37,    -4,     1,   -19,   -56,    12,    -6,   -12,    -1,    14,   -13,   -23,   -23,   -56,   -29,    33,   -31,    37,   -16,    26,    36,    37,    19,    40,    40,    46,    22,   -46,   -44,    -3,    -2,   -19,   -53,   -17,    34,    18,   -24,    -1,   -12,    11,   -51,   -73,   -20,    -6,    -2,    26,    -2,   -47,    28,     4,    27,    29,    63,    50,    16,   -38,     8,     5,    -3,   -13,   -46,   -33,    15,    47,   -17,    35,   -10,    16,     6,   -36,    -2,     6,    25,     9,     2,    41,   -30,    19,    12,    42,    53,    11,    90,   -10,     1,    -7,     3,   -18,   -31,   -40,   -13,    40,    -6,     3,     7,     0,    -5,   -11,    31,    30,    10,   -12,   -16,    11,   -26,    17,    27,    -9,    -7,    19,    64,    -1,   -58,     3,    -2,   -21,   -45,   -20,     7,    33,     6,   -16,     4,    26,    44,   -25,    -8,    26,    -1,    10,    -5,   -51,    14,   -23,    -7,   -27,    10,    43,    63,    -1,   -35,    -8,     4,     7,   -40,   -27,   -21,    -2,   -10,    29,   -27,     0,   -26,   -15,    12,    39,    27,   -18,   -36,   -31,     1,   -55,   -12,   -23,     3,    68,    61,    -6,   -33,    10,     8,    -3,   -41,    24,   -23,   -52,    24,    -1,   -26,   -74,   -44,   -31,    -2,    19,   -13,   -12,     5,    -9,   -15,    -9,   -18,    10,    37,    37,    10,   -23,   -20,     2,   -10,    -3,   -16,    41,   -35,   -27,    13,    19,     2,    -2,   -52,   -50,   -24,    44,    36,    31,   -15,   -54,   -22,     1,   -14,   -17,    -1,     2,    33,   -27,     4,     5,    -9,     2,   -27,    39,     1,   -56,   -15,   -48,   -13,     9,   -36,   -51,   -22,    22,    82,    43,    17,    41,   -26,    29,   -23,   -39,   -43,   -23,    26,     6,    -1,     6,    -5,    -8,   -17,    11,    -8,    -4,    18,   -36,   -18,   -23,   -39,   -49,    12,    32,    26,    10,    24,   -30,   -53,     9,   -35,   -19,   -43,   -50,    -6,    12,     6,     9,     2,   -11,   -15,   -17,    -3,    17,   -52,   -90,   -59,   -43,   -74,   -38,     7,    -7,   -30,   -43,   -21,   -36,   -54,   -28,   -76,   -83,   -86,   -90,   -22,    18,     1,     0,    -8,     1,   -12,   -23,    -6,   -10,   -28,   -38,   -74,  -102,   -78,   -58,   -13,   -13,   -69,  -127,  -133,  -112,   -68,   -17,   -62,   -67,   -44,   -77,    -3,    -6,    -7,     6,    -7,    -4,    -1,   -10,    -2,     1,   -15,   -15,    -4,    -3,    17,     3,   -34,   -57,   -56,   -80,   -40,   -65,   -79,   -23,   -19,   -20,     0,    -6,    -7,    -2,     1,     8,     9,   -10,    -4,     5,     1,   -12,   -19,   -18,   -14,   -10,     2,    -7,     1,    -4,   -10,     1,    -5,    -8,   -22,   -56,   -24,   -38,   -31,    -9,     9,    -4,     6,     5,    10,     0,    -6,    -6,     1,     7,   -12,   -10,    -9,   -10,   -27,   -13,    -5,   -21,   -14,    -9,   -10,   -12,     4,   -15,    -4,     4,    -4,     4,     2,    -2,    -7,     2,     1,     4,    -8,   -10,     2,     8,     1,    10,    -7,   -20,    -5,     8,     5,    -3,     2,    -1,    -2,     3,    -7,    -5,     4,     4,     6,    -9,    -7,     0,   -10),
		    97 => (   -2,     4,     9,    -9,     9,    -4,    10,     4,    -7,    -3,     0,    -1,    -1,     4,    -9,    -2,     6,    10,     2,     8,     3,    -3,   -10,     6,    -7,     3,    -1,    -3,     3,     6,     3,     8,    -7,    -8,   -10,     7,    -7,    -1,    -6,   -37,   -21,   -23,     7,   -18,   -45,   -65,    -2,   -15,    -2,    -6,    -3,     2,    -9,    -1,    -5,    -5,    10,    -3,    -8,   -10,   -19,    -4,    -8,   -17,   -10,   -37,   -40,   -78,   -12,    -6,   -16,   -31,   -19,     0,    -4,    -1,   -19,   -15,   -26,   -28,    -3,    -3,     1,     1,    -1,    -5,     8,   -17,    -6,   -50,   -45,  -102,   -89,   -76,   -89,  -110,   -97,  -110,   -57,   -25,   -23,   -21,     0,   -32,   -44,   -46,   -76,   -20,   -15,   -21,    -5,     3,     3,    -2,   -11,   -15,   -56,   -74,   -79,   -86,  -132,  -138,  -128,   -70,   -72,   -69,   -66,   -45,   -94,   -72,   -51,   -46,   -53,   -29,   -59,  -108,  -109,   -60,   -20,     8,     2,     2,     7,   -67,  -113,    21,   -52,   -18,    13,    22,   -36,   -25,     5,    32,    44,    -8,    42,    15,     2,   -50,   -90,   -57,   -36,  -122,   -83,  -104,   -50,    -2,    -1,    -1,    39,    40,    33,   -30,   -25,   -23,   -30,     3,   -11,     2,    19,     5,    18,    37,   -10,   -24,   -11,    12,    50,    35,    37,   -45,   -83,   -64,   -61,   -38,    -9,    47,    50,    18,    38,   -44,   -21,    10,   -12,    -2,   -17,    13,    23,    12,    18,   -23,   -22,    74,     4,   -17,     5,    -4,   -11,   -17,    -3,   -68,   -87,   -44,   -46,   100,    24,    -7,    23,    -1,   -30,    14,    21,    41,    36,    22,     3,   -17,   -27,    -2,   -13,    27,    46,    13,    31,     1,   -26,   -28,   -34,  -101,  -117,   -35,    10,    50,   -16,    10,    31,    23,    29,     8,    32,    62,    57,    10,   -46,   -21,    22,    20,     4,    30,    36,    -2,    39,    -2,    21,   -25,   -46,    -8,    -4,   103,     5,    40,    28,     0,    30,    27,    -7,    33,    55,    28,    30,   -38,   -66,   -17,    30,    67,    31,    -1,    25,    15,    46,    -1,   -14,   -38,   -38,    26,     2,    88,    -7,     8,    66,    16,   -19,    -6,    -7,    19,    32,    23,   -33,   -33,    26,    51,    89,    59,    41,     1,    33,   -22,    18,   -27,     1,    23,    14,   -73,   -41,    56,     1,    29,    63,    16,   -31,   -29,    -6,    -6,    24,     6,    17,    50,    42,    44,    88,    80,    51,    27,     5,   -46,   -15,    -1,    66,     2,    22,    46,    35,    51,     2,    15,    62,     0,   -51,   -30,    15,    -7,     3,    16,     3,    34,    43,    31,   101,    65,    43,    18,   -41,   -38,   -69,   -23,    10,   -21,     4,    45,   -14,   -39,   -11,    24,    26,   -42,   -64,    -7,   -12,   -35,    -5,     8,   -22,    15,     6,    14,    59,    12,    16,    26,   -21,   -21,   -31,   -60,   -19,    12,    40,   -42,   -51,    -2,    -5,    -1,    13,   -40,   -50,   -10,     5,   -18,   -70,   -62,   -26,   -16,   -25,     5,   -17,   -29,    -1,    24,    59,   -13,     9,     8,    55,    38,    35,    15,   -22,   -30,     2,   -14,    -4,   -32,   -15,    -5,     1,    -9,    -1,    39,    29,   -26,   -63,   -36,   -33,   -13,   -19,    69,   107,    83,    22,    68,    42,    63,    49,   -44,   -41,   -36,     4,   -14,   -12,   -21,    -1,     8,     1,   -34,    -2,    -1,    -1,   -45,   -75,   -26,     2,     2,    50,    73,    92,    17,    49,    31,    62,    51,     7,    31,   -12,   -54,    13,     5,    20,   -19,    -5,    36,    34,   -20,   -34,   -44,   -19,   -38,   -42,   -28,   -18,     7,    15,   104,    58,    31,    17,     9,    35,    13,     3,    11,     4,   -36,    -9,    20,     5,    -6,    14,    21,    21,    10,    22,   -40,   -21,   -22,   -39,   -53,   -25,   -27,    57,   107,    38,    34,     6,    18,     6,    -5,    31,   -10,   -40,   -12,     4,    25,   -10,   -25,   -66,    12,     3,    24,    21,     6,   -15,   -17,   -26,     1,     1,    19,     4,    23,    -7,    -4,    -4,    -5,   -26,   -24,    26,   -26,   -46,     5,    -1,     5,    -7,   -22,   -43,    37,    32,    36,    22,    43,    40,     6,    12,    11,   -19,    22,     7,   -33,   -51,   -39,   -22,    15,   -20,   -14,   -44,   -36,   -13,     7,    -3,    -3,   -26,   -44,   -47,    22,    62,    29,     5,     6,    20,   -11,    20,    14,   -12,   -43,    -4,   -55,   -42,   -47,   -52,   -39,   -73,   -71,   -45,     6,   -46,    -7,    -8,     9,   -19,   -79,   -40,    31,    58,    37,    21,    -3,    44,    -3,   -17,    -2,   -78,   -64,   -28,   -59,   -72,   -59,   -41,   -40,   -83,   -75,   -27,     6,   -37,     6,     0,     5,    -1,   -12,    -4,    42,    20,    36,    -1,     3,     0,    12,    -6,     1,   -45,   -55,   -36,   -29,   -83,   -76,   -64,   -18,   -70,   -78,   -44,   -39,    -6,     9,    -6,    -8,   -25,    49,    -4,    -2,     5,    13,   -34,    20,    17,   -10,   -14,    10,   -71,   -62,     3,   -46,   -61,   -84,   -53,   -13,    -4,   -54,   -21,   -10,    -6,    -3,    -8,    -4,    -5,   -53,   -36,   -51,   -28,   -26,     8,    56,    -9,   -16,    -4,    -5,     3,    10,   -13,   -50,   -13,   -12,     0,    23,    -4,    -2,    -8,    -1,     8,     5,    -1,     9,    -8,     2,    22,    27,     0,   -26,   -18,     0,    -1,   -40,   -12,   -23,   -43,    12,     4,    56,    23,   -23,     1,    29,    -3,    38,    -6,    -1,    -4,    -8),
		    98 => (    6,    -7,    -6,    -3,     6,    -4,     2,    10,     2,    -3,     4,    -5,     5,    -7,     1,   -10,    -9,    -4,     4,     5,     2,    -8,    -4,    -5,    -1,     3,     0,     1,     2,     8,     4,    10,    -7,     2,     9,     7,     4,     5,     0,     6,    -8,   -15,   -14,   -36,   -34,   -37,   -14,     9,   -12,    -8,     0,    -9,    -5,    -6,    -5,     5,     4,    10,    -9,    -2,    -1,    -2,     5,    -3,   -20,   -57,   -77,   -72,   -27,    -4,   -17,   -50,   -49,   -19,    -8,     2,   -12,   -18,   -28,   -19,    -1,    -1,     0,     2,     8,    10,   -12,    -6,   -12,   -30,   -23,   -97,    32,    46,    61,    24,    59,    67,    44,    23,     6,    21,   -18,   -45,   -36,   -58,   -35,    -4,   -12,   -16,   -10,    -5,     3,   -13,     9,   -10,   -61,   -70,   -14,    15,    21,    27,   -19,   -45,     6,   -17,   -11,   -17,    -7,     4,    -7,    19,     3,    15,   -63,   -34,   -14,    -2,     4,   -14,    -2,    -6,    -1,   -50,   -62,  -109,   -32,    20,    26,   -25,    -3,     9,   -56,   -32,    26,    -6,    13,    37,    22,     1,    30,    -3,   -25,   -39,   -32,   -12,    13,   -10,     8,    -4,   -58,   -28,   -24,   -33,     3,    84,    43,    26,    27,    12,     3,    14,    20,    35,    25,     2,   -32,    28,   -23,    -7,   -32,   -11,   -29,   -27,     3,    -4,    -9,   -37,   -22,   -48,   -16,    -4,    47,    69,   -40,   -16,    15,   -33,    -9,   -34,   -25,   -23,   -35,    -8,     1,    17,   -11,   -45,   -25,   -38,   -17,   -20,   -12,   -13,   -12,   -22,   -40,   -26,   -62,   -58,    18,    73,   -26,   -18,    39,    23,   -23,   -48,   -50,   -23,   -75,     9,     0,    10,   -15,   -19,   -10,   -50,     2,    21,    24,    -3,     6,    -5,   -16,   -12,   -76,   -57,   -10,   -22,   -25,     6,    46,    54,    24,   -27,   -35,   -20,    -8,    36,   -43,    -8,     1,    23,   -11,   -23,   -13,    11,   -64,   -60,     6,   -15,   -29,   -33,   -36,   -74,    21,   -33,   -94,   -21,    29,   101,    93,    62,    22,    -7,     6,    14,    14,   -50,    44,    24,     6,   -39,   -69,   -81,   -66,   -66,    -2,   -10,   -10,   -43,   -27,   -29,     3,    -7,   -35,    -7,   -72,     5,    49,    77,    55,    -1,   -18,   -41,   -15,   -17,   -12,   -12,   -32,   -32,   -75,   -54,   -17,   -24,     2,     5,   -18,   -10,   -17,   -38,   -20,   -53,   -79,   -81,   -96,   -95,     7,     6,    20,    62,    14,    -4,    20,    23,     6,    16,    14,    -7,   -11,   -42,   -30,   -21,    -7,    -3,   -21,    -6,   -25,   -14,    -8,   -45,   -78,  -111,   -85,   -63,   -49,    -3,    -2,    39,    15,   -15,    -7,   -26,   -53,     3,    16,   -56,   -51,   -40,   -35,   -11,    -5,    -7,     2,   -49,   -28,     9,    -3,   -30,   -40,   -58,   -10,    26,    12,    11,   -10,   -32,     1,     6,     2,   -43,   -22,    25,   -17,   -56,   -56,   -32,   -64,   -32,   -10,     8,   -30,   -35,   -45,   -23,   -29,     2,   -14,    10,    -1,    22,   -12,   -40,   -26,   -12,    30,   -21,   -40,     3,    -3,    23,   -49,   -35,   -39,   -33,   -72,   -26,    -2,   -10,   -19,   -18,   -35,    -5,    37,    28,     9,    49,     9,     2,   -39,   -10,   -63,     2,   -63,    42,   -32,    37,    37,    19,   -23,   -11,   -23,   -19,   -88,   -34,     7,    -4,   -27,   -69,    20,     9,   -20,    36,    32,     7,   -24,    -7,   -17,   -74,   -65,   -18,   -47,   -15,    15,    47,    12,    55,    44,    -1,   -37,   -30,   -17,   -41,   -10,    -6,   -14,   -23,    62,     0,    19,    44,   -10,   -39,   -26,    15,   -27,   -68,   -28,   -23,   -86,   -30,    18,    31,    28,    27,    23,    16,   -59,   -32,    -2,   -26,    -1,   -19,   -39,    42,    46,    61,    46,    21,   -46,   -26,     5,    15,   -65,   -41,   -45,   -13,   -27,    -5,   -25,     0,    17,    27,     4,   -36,   -53,   -21,   -76,   -25,    -8,    -4,   -33,     7,    41,    22,    31,    20,   -18,   -58,   -11,    11,   -47,   -11,    -9,    12,    27,   -26,   -28,   -21,    32,    26,    13,   -32,   -28,    -5,   -66,    -9,   -26,   -15,   -38,   -37,     9,    -3,     4,    -7,   -30,     2,   -24,    -4,    10,   -26,    29,   -18,   -21,   -39,   -61,    13,    29,    35,   -11,   -26,   -38,   -23,   -55,   -10,   -27,   -19,   -33,   -45,   -38,     5,    57,    41,   -34,   -22,     9,    17,    28,   -39,    -9,   -50,   -33,   -15,   -30,   -15,     8,   -20,   -58,   -21,     4,    -6,   -35,    -3,    -9,     9,   -10,   -18,   -56,    35,    11,    45,    11,   -38,   -20,   -36,     7,    -6,    -2,   -16,   -20,   -42,   -17,    -3,   -27,   -77,   -34,   -14,     3,    29,   -52,    -6,    -9,    -7,   -21,   -15,   -43,   -45,    22,    18,    12,    -2,   -36,   -31,    -6,     1,    24,    30,    48,   -29,     5,    -4,    -2,   -29,   -29,    -7,   -43,    -7,   -13,    -3,     3,     6,    -5,    -4,   -10,   -29,    -1,   -18,   -44,   -29,   -48,   -53,   -46,   -56,   -55,   -61,   -45,   -27,   -12,    -3,     0,   -24,   -10,   -11,   -11,    -3,   -10,     8,    -3,    -9,    -7,   -21,   -16,   -10,    -6,   -13,   -13,   -14,   -19,   -10,   -39,   -47,   -58,   -32,   -26,   -19,   -18,   -39,   -65,   -63,   -35,     5,    -1,    -8,    10,    -2,    -8,    -3,     8,     1,   -15,   -12,   -20,   -11,   -13,   -15,    -7,    -8,     0,   -35,   -12,    -8,   -15,   -15,   -16,   -11,     3,    -7,     8,    -6,    -4,    -6,    -8,     3),
		    99 => (    2,     5,    -2,    -1,   -10,    -8,    -7,    -8,    -8,    -8,    -1,    -3,     2,    -6,     4,     3,    -1,    -7,     8,     4,     0,     9,    -3,   -10,    -7,     3,     2,    -6,    -7,     0,   -10,     3,     3,     9,     6,     3,    -5,    -4,   -15,   -21,   -29,   -29,     6,    -8,     4,    -5,   -14,    -1,     0,    -4,   -14,    -6,    -3,    -1,     4,    -4,    -1,     6,    -6,    -7,    -6,     3,    -4,    -8,    -2,   -11,    -1,   -15,    -1,     5,   -21,     3,     4,     3,    -8,     1,   -14,   -16,   -20,    -3,     2,     2,    -9,    -3,     6,    -1,     1,   -22,   -10,   -16,   -15,   -10,   -34,   -28,   -16,    -3,     7,   -12,   -12,     3,    -5,   -14,   -15,   -18,   -34,    -8,   -29,   -17,   -33,   -22,    -4,    -9,     0,     2,    -4,   -10,   -13,   -14,   -53,    -4,     4,     2,     2,   -15,   -42,   -39,   -19,   -45,   -25,   -44,   -22,   -54,   -76,    -8,    -7,    -4,     3,   -48,   -15,    -5,     9,     7,    -8,   -20,    -7,     4,    -2,   -13,   -14,   -21,   -12,   -31,   -42,   -55,   -65,   -75,   -46,   -13,    -7,    21,   -29,   -24,   -26,   -13,    -6,   -15,   -22,     7,    -6,     7,    -4,   -22,    -5,   -22,   -31,   -28,   -48,   -14,   -29,    -2,    -7,    -5,    -3,     1,   -28,   -52,   -19,   -31,   -41,   -30,   -29,   -18,   -13,    -1,   -19,   -26,     4,    -7,   -11,   -19,   -18,   -32,   -59,   -74,   -74,   -38,   -29,     9,    -1,    23,     5,    14,    25,   -38,   -15,   -39,   -35,   -62,   -33,    21,   -23,    -7,    -8,   -18,   -35,   -30,   -13,   -20,   -40,   -50,   -58,   -80,   -52,   -41,     2,    11,    12,   -15,     7,     1,    37,   -36,   -14,    12,    -7,    -1,   -37,    -1,    -6,   -44,   -10,    -1,     0,   -37,   -28,   -36,   -47,   -29,   -53,   -15,     8,   -18,     3,    17,    23,    14,    16,    61,    16,   -20,     8,    40,     9,     0,     0,    -8,   -20,   -31,   -21,   -18,    -9,   -43,   -30,     1,   -23,   -34,   -49,   -23,     9,   -33,   -48,    23,    23,    14,    41,     6,    27,   -21,    40,    29,   -10,     5,    -9,   -37,   -34,   -34,   -14,   -27,    -2,   -80,    51,     1,   -15,   -20,   -24,    -3,    -1,   -22,   -61,     2,    12,    33,    20,    -5,   -29,   -41,    -2,     7,     7,   -13,     1,   -19,   -52,   -47,    -9,   -15,    -3,   -37,    17,    44,    37,     4,    21,     0,   -26,   -79,   -52,    -9,   -17,   -25,     3,    -3,   -14,    -2,   -10,    21,     0,    28,    -6,   -10,   -50,   -25,   -37,    -5,     7,   -39,   -14,    26,    23,    13,    24,    -6,   -28,   -94,   -26,   -12,   -66,   -62,   -37,     7,    -3,   -37,     7,     6,   -20,    36,    10,   -22,   -60,   -37,   -19,     3,    -3,   -27,   -34,    32,    28,    27,    -4,    -8,   -64,   -56,   -18,   -12,   -42,   -45,   -53,   -12,   -14,   -32,    -2,     9,    21,    24,   -16,   -44,   -50,   -28,     1,    -2,    -7,     4,   -49,    30,    45,    13,    15,     1,   -37,   -67,   -14,   -32,   -42,    -8,    -6,     3,     0,   -55,     7,    -7,   -11,    18,    19,   -49,   -57,   -31,     1,   -18,     4,   -15,   -30,    31,    58,    37,    67,    23,     9,    14,    10,   -40,     7,     1,     6,     0,   -59,   -39,   -29,   -40,     1,    -8,    39,    26,   -48,    -6,   -27,    -9,     3,   -11,   -77,    -5,    -7,    -2,    24,    38,    56,    42,    34,    47,    30,    -7,   -13,   -36,   -46,   -53,    -7,   -28,   -20,    -8,    34,   -11,   -48,   -17,   -34,   -32,    -8,     1,   -76,    22,   -21,   -37,    -8,    18,    -5,    -8,    47,    10,    -4,   -58,   -16,     0,   -18,   -16,    -4,   -51,    -9,   -21,    29,    27,   -23,    -7,   -42,   -22,    -8,   -12,   -43,    33,     1,   -43,   -38,   -26,   -55,   -48,   -18,   -18,     5,   -62,    18,     0,   -28,   -28,   -20,   -64,     1,   -39,   -11,    37,    43,    29,   -36,    -5,   -10,     0,   -16,    32,    25,    -9,   -29,   -39,   -57,   -34,   -46,   -25,   -72,   -51,    22,    19,   -29,   -54,   -20,   -30,    10,    -2,   -12,    39,    45,    80,   -41,    -7,     1,     7,   -28,    12,    14,    -7,   -24,   -26,   -31,   -53,   -35,   -13,   -10,   -33,    31,   -23,  -101,   -27,   -10,   -20,   -14,    30,   -31,     2,    19,    48,   -50,    -5,    -4,     7,   -32,   -24,   -43,   -15,   -22,   -36,   -21,   -32,   -18,   -33,    -7,    -7,    49,   -58,   -66,    -9,    -1,   -18,     1,     4,    -8,     7,   -17,   -47,   -11,    -4,     1,    -3,   -26,   -24,   -23,    -8,   -12,   -17,   -17,    -7,   -24,    -6,    -1,     3,    17,   -27,     8,    18,    -4,   -20,    39,    -2,    49,    20,    -1,   -20,   -12,    -5,     4,    -7,   -21,    -5,   -35,   -19,     2,    14,   -38,   -41,   -23,   -12,     4,   -10,    13,    16,    31,   -18,    -6,    -5,    35,    22,    30,    20,     4,   -10,   -10,     5,     0,    -8,    54,   -39,     0,    28,    11,     0,   -49,   -19,   -17,    -2,   -17,   -36,    31,    24,    14,    -9,   -17,    19,    41,    27,    31,     5,   -15,   -12,    -6,    -8,     1,     4,     8,    59,    30,    25,    27,    -4,     6,    35,   -29,   -10,   -15,   -43,     3,    15,    -5,    -7,    -5,    26,    41,    65,    34,     1,    15,     6,    10,    -3,    -2,    -4,    -9,     0,   -21,   -12,    19,    42,    34,    30,     1,     9,   -12,   -33,    -6,   -11,   -10,    -7,   -26,   -17,   -14,    -7,    19,   -22,    10,    -8,    -1,     0)
        );

 ---------------------------------INFO-
 -- COEF =86.27617

 -- MIN =-255.99998
 -- MAX =169.57208

 -- SUMMIN =-18188.84
 -- SUMMAX =13224.308
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
