----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (   -5,     1,    -2,   -11,   -12,    15,     2,     0,     9,   -12,    -4,    19,    -2,   -32,   -29,     7,   -18,    13,     8,     4,   -20,   -16,    -9,    11,    19,    20,    -4,   -17,   -13,   -14,    -1,     6,     3,   -16,    13,     7,    -2,     3,   -10,    13,    27,    18,   -28,    18,    53,    22,    -8,   -16,   -18,    14,    -4,     7,     7,    -2,     8,   -15,    13,    19,     3,    20,    53,     4,   -27,     2,   -31,   -86,    -9,   -16,    -7,   -49,   -46,   -74,   -11,   -16,   -30,   -12,   -11,   -12,   -45,   -33,   -29,   -37,     5,   -12,     8,   -19,    -6,    40,    -5,    29,    21,   -61,   -42,   -33,   -56,   -43,   -76,   -49,   -74,   -79,   -23,    52,     3,   -65,   -46,   -32,   -46,   -28,    19,    13,   -11,    12,   -13,    10,     4,    -5,   -28,   -71,    14,   -48,  -105,   -51,   -52,   -82,  -134,   -12,    -4,   -37,   -15,   -71,   -52,   -45,    -7,   -27,   -40,   -27,    10,   -21,   -37,     5,     4,    13,   -38,   -10,    -2,   -25,   -17,    -8,   -29,   -20,   -66,  -120,   -73,  -103,    15,    49,    -4,   -49,     5,   -69,   -85,     4,   -14,   -12,   -22,   -90,   -25,   -20,   -18,    19,   -41,   -27,   -27,    -2,   -22,   -19,   -40,   -41,   -36,  -129,   -92,   -37,   -11,   -43,    53,    39,     8,   -79,   -69,   -41,     9,   -87,   -37,   -83,   -23,    51,     2,   -37,   -34,   -33,    11,   -16,   -23,    14,   -30,   -36,   -83,  -132,  -129,   -47,    -4,     1,    85,    46,   -80,    -2,   -75,   -63,    25,   -46,   -75,   -29,   -80,    51,    61,  -104,    54,    36,   -12,   -18,   -24,    -3,   -15,   -71,   -45,  -126,   -27,   -24,    31,   -44,    19,    93,   -40,    16,   -82,  -101,   -22,   -56,   -29,  -102,   -36,   -25,   -24,   -18,    93,   -10,    -9,   -10,   -63,    -9,   -47,  -119,   -49,   -14,   -26,    31,   -21,   -32,    62,    15,     2,   -62,  -152,   -15,    -9,   -36,   -47,   -81,     2,    15,   -23,   -19,    23,    37,   -39,   -49,   -22,    32,    -1,   -11,   -41,   -26,   -18,    -5,   -94,  -101,   -33,   -70,    21,   -66,   -68,   -25,   -61,   -74,   -33,   -26,   -72,     8,     9,    89,   -38,    18,   -49,    -8,   -16,    -8,   -32,   -25,   -60,     6,    39,   -32,   -36,     9,   -52,    16,   119,   -86,   -69,    12,   -62,   -98,   -35,   -56,   -38,   -15,    -9,    28,    15,     1,    -5,    19,     5,    -1,   -97,    -2,    12,   -21,    45,   -19,   -39,  -101,    11,    59,   100,   -19,     4,    62,     0,  -103,   -67,   -65,   -53,    14,    -5,    44,    46,   -19,    -2,     9,    44,   -58,   -53,     7,   -20,   -74,    25,   -69,  -184,  -147,   -12,    50,    88,    26,   -13,    69,   -32,   -59,   -45,   -25,   -80,     4,    -8,    -1,     2,   -26,   -19,    36,   -44,   -60,   -49,   -12,    21,    35,    80,   -11,  -127,  -135,    -6,    16,    41,    29,   -72,     5,    -7,   -37,   -50,    14,   -64,    -5,     2,   -17,   -38,   -31,    16,   -65,    -3,  -100,   -51,   -83,   -18,    35,   109,    22,  -167,   -53,   -19,    23,    -9,   -26,   -74,    59,   -56,   -43,     6,   -41,   -49,    -7,   -16,     4,   -19,   -50,    14,     4,  -117,   -35,   -75,   -87,   -49,    49,    50,   -54,  -200,    -6,   -20,   133,   -39,   -23,   -56,   -48,    -1,   -48,   -52,   -38,  -112,    47,    -1,     8,   -68,   -34,   -89,   -26,   -59,   -55,   -64,  -157,    18,    24,    63,   -45,  -146,   -53,    -3,    66,    24,     1,    37,   -46,   -22,    25,   -46,   -60,  -109,    39,     2,     9,   -29,    22,   -30,   -51,   -23,   -12,   -50,   -82,    57,    57,   -52,   -82,  -167,   -18,    -8,     9,   -24,     4,    -1,   -15,    20,   -41,    -2,    -8,   -50,   -26,    16,    36,     7,    25,    10,   -44,   -21,   -82,   -60,    18,    45,    52,     0,   -90,   -94,    66,    20,   -54,   -41,    -1,   -77,   -33,   -34,   -30,     6,  -143,   -28,   -18,    -7,     2,   -18,   -36,    15,   -18,   -51,  -100,   -82,    25,     9,   -54,   -63,   -18,   -20,    16,    24,   -49,    -2,   -87,   -54,   -64,   -18,   -15,   -22,   -29,    15,    20,     5,    -8,   -47,   -52,   -23,   -25,     3,   -64,   -37,   -23,    18,   -21,     1,   -17,   -16,    39,   -20,   -19,   -54,   -79,   -78,   -42,    13,     7,   -74,     6,    31,    28,    -4,     9,   -38,  -117,    11,     7,    24,     5,   -38,    27,    11,    41,   -14,   -85,    67,    55,    59,  -120,   -50,   -64,   -56,   -39,    12,   -17,    -4,   -20,    28,    10,     6,     9,   -44,   -87,   -39,    16,   -32,    -9,   -39,   -87,    50,    28,    40,    55,   -61,   -55,   -67,  -143,     0,   -86,   -57,   -27,    41,    -5,   -31,   -80,   -43,   -15,    17,   -19,   -20,     4,   -50,    52,    25,    16,   -88,  -102,   -63,   -68,    12,   101,    22,    19,   -89,   -32,   -20,   -67,   -60,    33,   -37,   -48,    -3,   -13,   -19,     9,     4,    17,     6,   -14,  -143,   -56,   -53,   -51,   -23,   -52,   -86,   -98,  -147,  -137,  -168,   -69,   -43,   -50,   -54,   -39,   -72,   -28,   -48,   -37,    -4,     3,    -8,    -2,     3,    13,   -16,    -9,   -14,   -67,  -104,    11,    -6,   -65,   -37,   -19,   -54,   -42,   -49,   -49,   -25,   -74,  -110,   -46,   -79,   -48,   -21,    -1,   -19,   -12,   -15,     3,     8,   -19,    -4,   -18,    -3,    12,     6,    -6,   -10,   -20,    12,    -9,    10,   -49,    11,     1,   -30,     3,    19,     4,   -11,   -26,   -25,   -39,    -7,     2,   -20,    14),
		     1 => (   -4,   -10,    -6,    20,     3,    -7,     3,    -6,    16,   -16,     7,   -15,    -9,   -18,     9,    14,     2,     8,   -14,     8,   -20,   -10,    18,   -11,    -2,     8,   -16,    15,    19,    19,    18,    16,   -20,    19,     5,     8,   -19,   -10,    -9,   -18,   -32,   -21,    66,    49,    -2,   -32,   -20,    14,   -19,   -16,    -2,   -10,   -14,    14,   -10,    18,    12,     4,    -2,    16,     5,    -5,    16,    10,   -57,   -55,     2,   -16,   -16,   -18,   -32,   -67,   -78,   -91,  -114,    11,    37,  -100,   -30,    -5,   -17,   -28,     7,    17,    15,   -16,   122,    86,    -5,    14,    19,    98,    80,    51,    53,    29,    12,  -150,  -154,  -155,  -133,   -37,   -40,   -12,    17,   -79,    36,     6,   -54,    -5,    12,    15,    -1,    -3,    82,    71,    37,   -22,   -17,     2,    -2,   -16,   -58,  -140,  -136,  -165,    16,    68,     7,    13,    24,    34,    20,    35,   -41,  -166,   -87,  -140,   -83,   -78,     4,   -20,    82,   112,    35,     9,   -38,   -40,  -191,   -84,   -70,  -121,  -163,   -92,   -12,   115,    -8,   -12,    -4,    41,    46,   -47,   -69,  -159,  -118,   -86,   -84,   -68,    -6,    -8,    -1,    44,    39,   -34,    -4,    17,  -157,    11,    14,  -119,  -124,   -62,   -90,   -35,    -8,    37,    -5,    45,   -45,   -52,   -27,  -167,  -117,   -45,    -7,   -26,   -15,    -4,   -35,    35,    20,     3,   -33,   -63,  -173,   -38,   -90,  -140,  -105,   -19,    66,    30,    33,   -11,    77,   -17,   -63,   -43,    -1,  -105,  -113,   -46,   -49,   -36,     1,   -25,   -25,   -23,   -15,   -25,   -56,   -62,  -122,  -106,   -51,  -195,  -180,     3,    46,    36,    68,    42,    24,   -40,   -68,   -35,   -59,   -99,  -117,   -63,   -63,   -12,    14,    -4,   -25,    30,   -24,     2,   -91,   -45,   -35,   -55,  -139,  -257,   -61,   -14,   -31,     1,    81,    15,   -82,   -55,  -115,   -46,   -29,   -62,  -107,   -56,     3,   -63,     2,    24,   -11,   -27,   -10,   -11,   -80,  -104,   -69,   -92,   -14,  -131,  -102,   -51,    17,    95,    80,   -13,   -79,   -72,  -105,   -40,   -39,   -50,  -113,  -125,    -6,   132,     4,    -3,    20,    34,    37,     9,   -52,   -62,  -103,  -167,   -87,  -142,   -39,   -58,    -2,   118,     8,  -105,   -60,   -33,   -37,    18,   -32,   -68,  -123,  -113,    -7,   113,     3,     5,   -37,    90,    22,   -23,   -32,   -24,  -161,  -137,   -78,   -76,     5,   -36,    79,   -16,    46,  -164,  -176,   -60,    78,   106,   106,    73,   -31,     1,   -17,    69,     7,   -17,    -4,    26,    43,   -32,   -41,   -13,   -80,  -183,   -83,   -43,   -29,    23,    92,   -38,    32,  -151,  -174,    14,    69,     9,    -8,  -134,   -76,     5,    37,    13,   -15,    14,    42,    41,    52,   -98,   -59,   -41,   -21,  -117,   -80,    30,   -15,   -65,    92,     3,   -70,  -151,   -11,    92,   103,   129,    73,   -38,   -60,   126,   120,     2,    15,     6,    47,   116,    48,   -13,   -29,   -12,    69,     7,   -28,    70,     4,   -40,   -35,   -96,   -73,  -120,   -44,   -98,   -15,   138,    57,   -72,  -165,    41,    25,   -13,    10,    17,    15,   -50,   -39,   -10,    27,     7,    69,    44,    37,    81,    33,    37,   -65,   -30,   -26,  -142,  -120,  -128,   -14,   103,    68,   127,   158,   -40,   -28,    -8,    12,   -11,    24,   -57,    20,     9,    61,    22,    47,    17,    21,    33,   -12,    25,    27,   -34,   -62,   -48,    27,    56,    72,   122,   134,   150,    91,    -5,   -25,   -54,   -45,   -10,    -3,   -35,   -38,   -49,   -57,   -25,    21,   -65,    19,   -31,   -12,    49,   -71,  -153,  -118,    28,    78,    88,    53,    10,    10,    -3,    42,    82,    12,    58,    -9,   -17,    65,    64,   -75,    61,    77,    21,     7,   -67,   -14,    35,    32,    42,   -91,  -112,  -171,   -28,    53,   -14,   -14,   -28,   -88,     9,    84,   109,    22,    55,    -4,   -12,    66,    21,    -1,   108,    44,   -68,    -3,   -26,   -74,    28,    -4,    43,   -48,  -128,  -144,   -36,   -39,   -14,    82,   -89,   -52,     1,    42,    39,    46,    -1,    83,    54,   -25,    -6,     3,   -89,  -144,   -49,     6,   -30,     5,   -26,    41,   -60,    -2,   -32,  -123,  -130,  -109,   -37,    48,    29,    28,    39,    56,    55,    13,    11,    61,    69,    10,    -2,     7,   -76,  -171,   -31,    -6,   -45,    33,   -47,   -13,   -20,    50,   -57,   -42,  -107,    10,    76,   122,    43,    78,    56,    69,   104,   163,    19,   -16,   -16,   -19,     6,   -58,   -12,   -56,   -70,    68,   -42,   -19,    40,    -1,     9,    34,   -13,    19,    20,    36,    98,   119,     9,    -9,   -27,    51,    81,   158,   -10,     0,     7,   -15,   -22,   -50,   -89,   -27,   -78,   -47,   -78,  -136,   -40,   -64,  -154,    56,    49,   -19,    22,    17,   200,   135,    22,   -12,    20,   -35,    27,    41,    -5,    12,    14,    -2,    -6,     2,    -8,   -13,   -19,   -67,    41,  -134,   -71,  -107,   -89,   -92,  -147,   -56,   -85,   -57,   -62,   -79,   -68,   -42,   -35,   -25,     5,   -19,    16,    -9,   -15,    -8,   -14,   -34,   -68,   -86,   -43,   -52,   -66,    25,   -12,  -106,  -100,  -134,  -140,  -109,   -76,   -17,   -37,   -20,   -17,    -5,    11,   -19,     9,   -15,     4,    -8,    -4,   -20,    12,    17,     7,   -11,    -9,   -11,   -16,   -20,   -28,    13,    13,    25,    -6,   -13,    -7,   -19,   -17,    -2,     9,   -14,    16,    18,     5,    11,    14),
		     2 => (    0,   -15,     9,   -17,   -15,     8,    11,     8,    -1,    14,     5,   -19,    -2,     5,     2,     7,     3,   -20,    -7,     2,     2,    11,    -1,     8,     4,   -15,    -7,    -9,    -1,    10,     0,    -4,    16,    13,   -14,    16,   -40,   -58,   -39,   -32,   -18,   -89,   -65,   -22,    -4,    23,    -5,   -19,   -23,   -13,   -15,   -35,     7,     9,    19,    13,     7,   -15,     3,   -53,   -60,     3,    15,  -104,   -27,   -44,   -45,   -74,   -39,  -198,   -58,   -10,   -31,   -46,   -84,  -102,   -78,   -17,   -45,     8,    24,    44,    12,    15,    -8,    15,   -30,   -82,   -79,    -2,    89,   -36,   -13,    83,    86,    11,   -86,  -111,   -63,  -112,  -103,   -38,    54,   -35,  -115,   -67,   -13,   -45,   -56,    25,   -15,   -17,   -16,    19,    -6,    48,   -27,   -53,   -10,    85,    18,    -8,   -84,   -62,   -53,  -125,  -129,   -84,    33,    31,     8,   -41,    44,    63,   -15,   -97,    15,    12,   -53,   -21,     0,    15,   -28,    13,   103,    23,    -4,    -4,   -19,   -34,   -97,  -135,  -143,  -138,  -108,   -52,   -20,    11,    63,    71,    50,    84,    20,   -73,   -59,     5,   -56,   -12,    19,    19,    33,     9,    18,   -22,   -27,    50,    25,   -34,   -35,   -54,   -23,  -140,  -108,   -93,   -53,    85,    32,    58,   -23,    24,    13,  -114,   -97,    97,   -59,   -10,    11,    14,    83,     4,    -4,   -51,    -7,    57,    -6,    21,    -1,    41,    28,    61,   -51,   -52,   -42,   -34,  -106,   -27,    35,    24,    11,  -188,   -22,   136,   -69,    -9,  -106,    96,    89,   -57,   -39,    34,    -4,   -31,   -54,  -108,    10,    71,     2,    31,    44,  -128,  -162,   -58,   -69,    17,    43,   -16,    -8,    19,    23,    68,  -100,   -25,     3,   -47,   101,   -49,   -87,   -18,   -19,     2,   -69,   -49,    32,   -38,   -63,     8,    32,    20,   -49,   -43,   -16,    80,    24,    38,    31,   -19,   -17,   -95,    69,   -33,   -18,   -36,    83,  -106,   -56,    53,    50,    72,    -9,    -2,    24,     5,    46,   104,   193,    60,   -70,   -37,    11,    90,    31,    44,    15,   -88,   -48,   -70,    47,   -51,    14,   -77,   -57,   -72,    50,    14,    48,   103,    90,    51,   -52,   -39,  -109,   -36,     8,     5,     0,   -89,    -8,    55,    -3,    25,    19,   -91,    -3,   -28,    28,   -83,   -16,     5,  -163,   -45,    85,    61,    53,    54,    -4,    26,     5,  -120,  -138,   -73,   -58,   -53,   -71,   -63,   -55,    24,    41,     8,    -9,  -143,   -25,    21,   118,    -7,    -5,     6,   -10,    65,   -22,   -74,  -102,  -106,  -192,   -56,   -45,     0,   -72,  -131,   -80,  -101,   -57,    -6,   -12,   -16,   -40,   -76,   -31,   -30,    48,    68,   179,    24,   -17,    -6,   -28,     8,  -102,  -145,   -50,   -68,  -118,  -139,  -108,    35,    47,   -89,  -133,   -50,    46,    30,   -26,   -51,  -129,   -88,    19,    31,     2,    69,   135,    47,    13,   -26,    13,    26,    34,   -30,   -72,  -162,   -79,   -92,    31,    16,    75,    39,    -3,    38,   -40,    43,    42,     3,   -25,    -1,    11,    26,    36,    29,    50,    78,   -10,     7,    12,    45,    73,    30,   -45,     8,   -35,   -21,    18,    27,    46,    -1,    86,   100,    88,   138,    -8,   -97,  -173,   -97,   -43,   -27,   -39,    26,    88,    72,    15,   -28,    54,    65,     5,    52,    -5,   -57,    -8,   -30,    49,   -36,    98,    -6,     9,     4,    28,   -19,   -49,   -82,   -43,   -16,    15,   -20,    10,   -10,    77,   116,    11,     4,   -67,   129,    76,   132,    89,    -9,   -52,   -22,   -13,   -60,   -28,    41,    33,    79,    42,    -9,   -23,   -31,     3,   -31,     3,   -11,   116,    19,   104,   186,    13,   -16,   -16,   113,   148,    67,    59,    21,   -13,   -35,    94,    49,    45,   -19,   -18,    31,    55,    44,   -11,   -82,   -44,    -8,    63,    38,   129,    72,   135,   144,   -12,    17,    24,    59,    77,    79,    90,    66,    24,     5,    -7,    -1,   -60,     0,     0,    77,    49,   -34,   -24,    -6,   -45,    -2,   -36,    63,   121,    32,   134,   -20,    -5,    30,    15,   -11,    76,   111,   -22,   -38,   -25,   -24,   -39,   -67,   -66,  -151,   -72,    23,    12,    56,   127,    99,    52,   -90,    -6,    79,    89,    84,   116,     4,     0,   -17,    56,    32,    93,     1,   -76,   -89,   -63,   -54,   -77,  -102,  -123,  -162,   -68,     9,   -23,    60,    54,    23,   -54,   -22,   -17,    22,    77,   -54,   -70,     0,   -19,     2,    34,    39,    47,    14,   -11,   -34,   -19,   -77,  -103,   -94,  -142,  -111,   -86,    19,  -131,  -236,   -77,     8,   -11,    12,   -60,   -72,   -18,    37,   -22,   -12,    17,    17,   -50,    36,   -59,   -77,   -20,   -49,   -18,  -150,  -161,  -143,  -137,  -156,   -74,   -65,  -178,  -264,  -137,    41,    17,    38,   -58,   -28,    54,     3,    -7,   -17,    -4,     7,   -12,   -41,   -79,  -111,  -112,   -92,  -110,  -129,  -135,   -73,   -48,  -124,    25,   -39,  -101,   -94,  -199,  -176,   -87,    11,   -65,   -79,   -32,    13,    17,    -3,     5,   -15,    -5,     8,   -61,   -65,   -65,   -73,   -50,  -161,   -82,   -30,   -41,   -67,   -35,   -97,   -92,  -120,  -155,  -167,  -118,  -105,  -104,    -2,   -20,    14,    20,    -1,    12,    13,     6,     8,     3,   -16,     2,     1,   -14,   -12,   -70,   -51,   -11,   -57,   -44,   -48,   -43,   -29,   -33,   -43,  -121,  -131,   -45,     0,     5,    -6,    13,    -6),
		     3 => (   -3,   -18,     0,    19,     0,   -13,    13,    15,    19,     1,   -17,   -13,    -9,   -22,    -2,    -2,    19,    16,    16,     9,    -5,     0,     7,    14,    15,    19,    -9,   -13,    10,     8,    14,     5,    19,   -11,   -14,    -7,   -18,   -11,     5,   -13,   -31,    -8,   -19,   -38,   -51,   -44,    11,     7,    14,    13,     1,     0,    -1,   -17,   -17,   -13,   -10,    17,   -19,    17,   -10,    17,   -25,   -22,   -20,   -75,   -79,   -25,   -68,   -87,   -54,   -65,  -110,  -136,  -117,   -62,  -168,  -145,  -162,   -51,   -13,     2,     3,    14,    18,   -13,    12,   -21,   -18,   -48,   -25,   -58,   -58,   -58,   -88,   -64,    -7,   -19,   -75,   -78,    13,    91,    55,   -42,   -21,   -39,  -116,  -150,   -72,   -13,    -8,   -10,     5,    20,   -19,    32,    90,    39,     3,    54,    70,   110,    90,    -9,     4,    41,    75,    15,   -69,   -23,    56,     5,   -19,  -135,   -61,  -256,  -167,   -11,   -46,     9,     9,     3,     9,   -30,    31,   -46,   -57,   -81,    24,   -67,    37,    35,     7,    -9,   -15,     3,     0,    36,    64,    25,    23,    66,    27,   -37,   -60,   -46,   -45,    -3,    15,    17,    11,   -15,   -52,   -21,   -13,    -1,    48,     3,    14,   -12,    35,   124,    51,    -4,   -15,     1,     6,    75,   -79,   -46,    15,    -1,    -4,   -68,   -85,   -12,    10,    32,     0,   -75,   -39,   102,     8,    -9,    19,    -2,    46,    81,    17,   -44,    23,    53,    77,    -7,   -14,     5,    82,   -21,   -60,  -129,   -76,  -113,   -76,   -18,    14,    -8,    17,   120,    54,    30,   -57,    63,   -16,  -100,    61,    38,    88,    25,     0,   -38,   -22,    29,    -9,     8,    45,    54,   -24,  -200,  -229,   -62,   -93,   -18,   -20,   -53,   149,   122,    26,  -132,   -40,   -16,   -53,   -16,   -85,   -66,  -155,  -190,  -294,  -130,    31,    10,    29,    46,    56,    26,    14,  -144,  -294,  -121,  -131,     6,     4,   -35,   196,    85,   -73,  -146,  -168,  -237,  -198,  -215,  -197,  -351,  -288,  -260,  -108,   -33,     8,   -36,   -23,    16,    16,    69,    43,   -53,  -265,   -71,   -72,   -21,     4,   -26,   -26,   -51,  -108,  -150,  -230,  -166,  -233,  -313,  -217,  -186,   -92,    72,   105,   106,    12,    37,     1,    53,   129,    85,    60,  -147,  -133,  -116,   -49,    -1,   -16,    -6,   -74,  -107,    33,   -40,   -33,  -102,   -47,  -100,   -42,    15,   109,    99,    70,   -30,     9,   -36,    55,   -95,   -20,   -12,   -31,   -47,     6,   -18,   -25,   -18,     8,    -1,   -99,    19,   123,    76,    -4,   -52,    11,   -44,    26,    88,    48,    71,   -34,    -7,    -5,   -73,   -86,  -125,   -82,   -12,   -39,    -4,   -78,   -81,   -36,   -22,   -26,    24,    -9,    -3,    18,   107,   -40,   -72,   108,    33,    -9,    37,    37,    37,    -9,    10,    -7,   -22,   -11,   -57,  -100,   -25,   -79,   -94,  -112,  -200,   -58,   -32,   -34,    58,    78,   -27,    66,   -23,  -137,  -177,  -108,   -69,    14,    31,     0,    85,    79,   -22,   -25,    12,   -20,     5,   -34,   -10,  -110,   -13,   -81,   -66,   156,     2,   -12,     8,    70,    83,    48,    -2,  -217,  -162,  -233,  -135,   -74,    15,   -18,    50,   -27,   -49,    10,     4,    -2,    41,    20,    54,   -83,   -49,  -126,   -67,    56,   -14,     0,    30,    99,   -11,  -100,   -31,  -150,   -51,  -167,  -308,  -373,  -153,  -168,  -166,   -91,   -64,    43,    38,    43,     3,   -26,    47,    13,   -66,  -125,  -128,   -56,   -23,   -38,    25,   133,    33,   -76,    57,    20,    93,   -11,   -41,  -128,   -88,  -189,  -179,   -72,    31,   -32,    -1,   -26,    39,    68,    50,   -10,  -164,  -231,   -83,   -54,   -46,   -16,   -21,   -90,   152,    23,    24,    43,    16,    45,   -40,   -37,   -85,   -66,    40,    -5,    -4,   -19,   -25,    -4,    -4,   -21,   -44,   -77,  -103,  -170,   -70,   -61,   -34,   -18,    13,  -160,   117,   101,     6,    -6,    -1,    61,     9,    44,    36,    36,    37,   -34,   -61,    -5,     3,   -33,   -31,    -7,   -71,  -121,  -155,  -141,   -39,   -34,    -9,   -39,    18,   -22,    55,   120,    -6,   -47,    30,    94,     4,    64,    28,    12,   -55,   -42,   -71,   -84,    24,   -14,  -100,   -47,   -45,   -82,  -166,  -130,   -49,     0,    11,   -10,   -34,   -11,    49,    36,    55,   -38,   -69,   -18,   -54,    -6,   -13,   -61,   -41,   -57,   -32,   -17,    49,   -91,   -16,   -97,  -111,  -163,  -155,  -128,   -56,   -14,   -11,   -20,    12,    88,    81,    14,   109,   -69,    20,   -50,   -14,   -35,    21,   -23,     1,    35,    -8,   118,    -7,    -1,   107,   -54,  -129,  -217,  -164,   -72,  -112,    -9,     0,    -4,     1,   -14,    36,   -44,   -50,    13,   -38,   -41,    26,   -30,   -48,   -47,  -102,   -27,   -68,   -58,   -99,   -40,  -124,  -133,  -110,  -131,   -52,   -66,   -10,     8,    -1,    -4,     6,     7,   -79,   -31,   -13,   -60,  -101,   -66,   -12,    29,   -96,    -7,   -19,   -52,  -147,  -148,  -134,   -51,   -33,     2,   -48,  -120,   -78,     7,   -28,    11,     3,   -13,   -15,    -4,   -60,   -20,    15,   -55,  -101,  -146,  -162,   -60,  -101,    37,    99,    63,    10,   -66,   -81,   -51,   -62,  -105,   -66,   -84,   -12,    15,   -10,     9,   -15,    12,    11,    11,     4,    -7,    -5,   -23,     3,     3,   -46,    -7,   -31,     4,   -25,   -59,    -7,   -63,   -54,     7,   -12,   -42,   -12,   -16,   -12,    -3,    12,   -12,    -3),
		     4 => (    8,    -9,     6,     3,   -10,    18,    13,   -14,    -9,    -7,   -15,     1,   -29,   -30,   -36,   -11,   -11,   -17,    -5,    15,     7,    -2,     9,    -1,   -19,   -11,   -13,    -5,    15,    -4,     5,   -19,    -5,     3,   -55,   -72,   -25,   -30,   -69,   -26,   -77,  -131,   -58,   -61,   -69,   -51,   -19,     8,   -48,   -27,   -44,   -56,     8,     5,    17,    -7,    11,     3,   -11,    15,   -70,   -19,   -75,   -86,  -128,   -56,   -61,  -138,   -85,   -89,   -52,   -50,  -121,   -99,   -94,   -22,  -119,  -108,   -95,   -81,   -25,   -69,    19,   -12,   -14,     4,    -9,   -56,  -144,   -70,  -105,   -61,   -65,   -86,   -46,   -90,   -98,   -84,   -81,   -90,  -143,  -173,   -84,   -19,     9,   -14,   -37,   -24,   -80,   -51,   -15,   -10,   -14,   -11,   -36,  -132,   -20,    22,   100,    27,   -42,  -124,   -82,   -42,   -36,  -115,  -195,  -152,   -88,  -141,   -78,   154,    72,    21,    95,   -55,   -67,   -34,   -61,   -16,   -13,    -8,   -67,   -49,   -11,    22,    86,   -31,   -21,   -41,   -38,   -38,   -27,  -168,  -195,    22,   -82,    27,   -65,    22,    11,    16,    18,  -113,   -49,   -34,   -34,   -16,    11,    -3,    -6,   -15,   -50,   -44,    93,   -80,    35,    63,    17,   -66,  -132,  -277,  -256,  -142,   -36,    22,    96,     0,    -3,    18,   -88,  -116,  -127,   -34,    -5,   -48,    11,   -77,   -18,    13,   -23,   -35,    44,    -7,    19,    23,    35,    36,  -122,  -220,  -306,  -123,   -50,   145,    98,   102,    38,   -16,   -77,  -111,  -109,    -5,   -30,  -113,   -72,  -172,    14,   -15,    40,    38,    57,   -17,    36,    96,   -15,   -34,    13,  -240,  -215,   -94,   133,    91,    54,   -34,   -79,    41,   -12,   -43,   -66,    13,  -104,  -154,   -13,  -114,    21,    19,   108,    49,  -130,   -24,    72,    10,    52,    62,    87,  -119,  -169,   -10,   194,    31,    19,     0,   -96,   -34,   -42,    11,  -117,    23,   -97,   -77,    17,   -59,    -2,    49,    36,   -14,  -230,   -58,    32,    81,   -18,    38,    81,  -124,  -136,    90,    90,    14,    68,    52,   -60,  -121,   -76,  -147,  -150,    33,    -6,   -50,     3,   -88,    30,    18,    57,    15,   -83,   -17,    31,    24,    52,    55,    14,  -184,  -188,    17,    48,    -4,    26,   -43,  -112,  -115,   -55,  -106,   -45,    31,   -37,  -116,    14,   -54,    41,    54,    56,    59,    15,    15,   -79,   -49,    46,     2,    17,   -52,  -124,    55,     6,    10,    -4,    18,   -76,     2,    80,   171,   168,   137,  -129,   -90,    -2,   -42,   -78,    -1,    91,    34,   -27,    -4,   -25,    43,    82,    -3,   -10,   -15,   -45,   -54,    31,    -9,    55,     5,    22,    86,   160,    80,    22,   -12,  -124,     3,   -14,   -12,   -80,     8,    44,   127,    20,    81,    39,   -14,    -9,   -25,   -40,   -21,   -87,     8,   -34,    23,    33,    79,    11,   113,    92,   -19,    50,   -45,   -73,    -9,    15,    19,    21,   -21,   102,   -11,   -10,    82,    -1,    11,     2,    27,    12,    71,    51,    72,    54,    26,    33,    78,    -3,   -21,    35,   -69,   -96,  -100,    40,   -16,   -18,   -13,  -113,    61,   104,   -53,   -64,    89,     6,   -32,    15,     7,   -13,    26,    76,    65,    -6,   -46,    51,     1,   -13,    34,   -75,  -104,   -14,   -32,   -46,     3,    -1,   -15,   102,    75,   157,    -1,   -99,    20,   -62,    14,   -92,   -66,   -33,   -45,    19,   -66,   -88,   -86,   -13,  -147,   -51,    26,   -43,   -61,     3,   -24,    13,    11,   -74,   -12,    77,    90,   113,   -80,   -92,  -101,   -55,   -22,   -61,   -85,   -53,   -39,   -47,  -145,  -105,   -49,   -97,  -103,   -39,    14,    17,   -27,   -39,   -55,    17,    -3,    -8,     2,   -26,    38,   -12,  -124,   -21,  -136,   -74,   -26,   -17,   -10,   -79,    -6,    20,   -16,   -96,    36,   -73,   -24,   -37,   103,    33,     7,   -49,   -77,   -18,     0,     0,     0,   -23,   -83,  -186,  -120,  -109,   -26,   -88,  -106,   -67,    80,    29,   -11,    22,   -13,   -18,   -21,    58,     5,   -49,   -33,    -5,   -17,   -13,  -163,   -23,   -18,   -55,   -52,   -32,  -107,   -71,  -115,   -87,   -83,   -32,   -91,   -37,    13,    14,   -29,    48,   -87,    23,   -63,   -35,   -56,   -83,  -129,   -33,    35,    10,  -137,   -76,   -10,   -23,   -48,   -18,   -53,   -23,    -1,     7,  -101,    21,  -139,   -99,     6,    15,   -47,   -18,   -50,    -9,   -43,   -27,   -88,   -74,  -111,    19,    59,    -7,    15,    34,   -11,   -16,   -19,   -28,   -56,     1,   -39,    62,    59,    13,  -170,   -19,   -55,   -57,   -52,   -39,   -60,     5,     6,    79,   -80,  -101,   -19,   -44,    29,   -48,    36,     8,   -11,   -14,    18,    -9,    13,  -140,   -38,   -57,   -38,   -10,   -32,   -80,   -36,   -70,   -51,   120,   -19,    76,    71,    99,   -91,   -11,    16,   -13,    -7,  -118,     6,   -34,   -11,     7,   -13,    -9,   -18,   -10,   -85,  -230,  -133,   -95,   -64,   -95,   -88,   -86,    16,    34,   -76,    -7,    36,     7,   -48,   -15,    53,   -62,    28,   -55,   -24,   -26,    19,   -15,    -8,    15,   -27,   -36,   -16,   -61,  -103,    24,   -22,  -120,  -203,  -177,  -136,   -61,  -102,  -179,   -43,  -110,  -141,  -179,  -169,  -140,   -32,   -52,    -4,    18,   -12,    20,     0,    -8,    -7,   -11,    10,   -61,   -52,   -71,   -77,   -62,  -133,   -72,   -55,  -152,   -44,   -66,   -88,   -68,   -95,  -116,  -102,   -80,   -26,   -11,    -2,     4,    17),
		     5 => (   13,    -6,    -9,    10,    17,     2,     5,     8,   -10,    16,    14,    -1,    -6,     5,    -1,    17,   -11,   -14,     8,    17,   -18,    -6,     6,    -4,    11,    19,    10,    16,    19,     8,    18,   -14,    12,   -18,     3,     5,    14,    19,    13,   -14,   -41,   -38,   -40,   -37,   -25,   -42,   -13,   -10,   -24,    -6,    -5,    -1,   -17,    13,   -16,    20,    17,   -13,    -3,   -20,   -19,   -14,     9,    11,   -23,    -7,   -70,  -141,  -128,  -177,   -62,    66,    60,    76,   111,    91,   115,    87,    85,    96,   -43,   -24,     6,   -20,    14,    14,   -10,    30,    76,   -17,   -46,   -36,   -29,   -99,  -114,   -89,   -36,   -88,    71,   -33,  -133,  -103,   -12,   -25,    36,    57,   -39,   -17,    53,    45,    60,    20,     9,   -30,   -39,     9,  -101,  -101,  -127,  -149,  -210,   -68,  -161,  -106,  -105,     2,   107,     6,    38,    -4,    -2,   -11,    20,    57,    78,    87,   109,   215,    58,   -18,    -3,   -15,   -21,   -15,   -93,   -88,  -183,  -180,  -217,  -113,   -16,    -9,    37,     3,    13,   -27,    32,    80,    46,    12,   154,   130,    72,   129,   141,   203,    96,   -30,     8,    -2,    39,   -31,   -95,  -165,  -166,  -102,   -52,   -96,   -26,    16,    99,     8,    -1,    10,    43,    73,   153,    21,   126,     1,    11,   122,    44,    99,    67,    17,    -6,    18,   -15,   -55,   -81,  -110,   -48,   -10,   -32,     6,    -1,    91,    60,    22,   -36,   -52,    17,    54,    68,     6,    68,    -3,   -72,   -14,   -43,    41,    49,    33,   -18,   -23,   -60,   -49,   -65,   -41,  -101,   -47,   -78,  -109,    37,   110,    61,   -80,   -73,  -123,  -244,  -133,  -125,  -323,  -153,  -176,  -123,   -47,   -28,   -14,    35,     8,     0,   -31,  -122,  -137,  -124,   -18,  -117,  -134,  -114,   -61,   -56,   -33,   -41,   -70,  -133,  -306,  -383,  -440,  -477,  -460,  -323,  -246,  -225,  -125,   -77,   -63,     4,    22,     9,   -25,    -9,   -70,   -12,   -38,   -74,   -47,    -9,   -49,   -59,    12,   -60,    11,   -95,   -29,     7,   -94,  -276,  -284,  -277,  -229,  -217,  -147,   -83,     1,    13,    12,   -12,    -6,    -9,   -45,   -15,   -49,   -83,   -84,   -66,   -78,   -61,   -36,   -35,     0,   -45,   -41,    34,    10,    40,   -45,  -138,  -231,  -168,   -77,   -89,   -16,    27,   -37,    11,   -14,     0,   -44,   -11,   -38,   -36,   -69,   -39,   -67,   -32,    33,    30,    26,    28,    11,    20,   -44,   -42,     2,   -43,   -79,  -122,   -86,   -34,   -30,     0,   -56,    -7,    -1,   -15,   -18,    -7,    35,   -53,    12,   -85,    31,    64,   116,    47,   -24,    45,    11,    -9,   -23,   -59,    19,     9,    45,   -50,   -32,   -67,     4,   -10,   -33,    34,   -18,   -11,    13,    67,   -67,  -114,   -97,   -20,   -32,    70,    10,     4,   -40,    17,   -77,    63,    12,    10,   -71,     2,    12,    -2,     2,   -28,   -20,   -35,   -31,    -3,   -56,   -36,   -27,    60,   -69,  -113,   -82,   -98,   -52,   -51,   -27,    42,   -48,   -92,   -25,   -73,    40,   -26,   -18,   -54,    18,   -10,    23,    19,   -17,   -18,   -10,    -1,    13,   -50,    17,    -1,  -100,  -106,  -158,  -162,  -261,  -207,  -128,    23,    17,   -69,    29,    24,   134,   -28,    43,    28,    35,    47,   -65,   -85,   -53,   -56,   -57,   -11,   -39,  -107,    26,   -51,   -62,   -76,  -161,   -75,  -202,  -276,   -93,  -113,  -149,  -116,    32,   -36,   -54,   116,    60,    70,    45,   -32,   -48,  -122,   -62,   -23,   -37,    -5,   -27,     7,    58,     4,   -53,   -84,   -22,    65,   -39,   -11,   -74,  -206,  -107,    -9,   -49,    27,     1,    79,   -39,    -9,    32,    -7,   -40,  -117,    16,  -100,   -77,     3,    -3,    84,    -7,    14,   -69,   -14,   -27,    43,    69,    21,    63,    46,    28,    40,   -20,    40,   -16,    32,    28,    27,   -39,     2,   -66,  -105,     7,   -29,   -40,   -14,   -10,    56,    29,   197,    -9,    22,    -7,   103,    72,     9,    28,   -76,    84,    76,    31,    10,    -4,   -38,    58,    43,   -52,    65,  -117,   -78,   -51,   -17,     7,     9,   -24,   -53,   -28,   125,   103,     3,   -21,    23,     5,    37,    67,    34,    45,   -18,    31,    39,   -45,   -69,    44,    69,    81,    71,     9,   -40,   -62,    -5,   -15,    14,     7,   -76,    17,   -57,   -34,   -58,   -32,   -43,   -32,   102,    19,    50,   -45,    -6,   -41,     8,   -22,    31,    12,    98,   -38,   -38,   -49,   -70,   -59,    -4,     6,     4,   -15,    37,    49,   -61,   -54,    23,    11,   108,    58,    17,   -90,   -36,   -35,    -4,   112,   -17,  -112,   -96,   -79,   -96,   -78,    10,    34,  -158,  -163,    22,    -3,   -19,    -3,   -69,    -7,    90,    74,   220,   106,   -19,    65,   133,    -1,    36,    23,    80,   -68,  -107,   -52,   -84,   -97,   -19,    55,    72,   -13,     4,   -47,   -55,    14,   -16,    -3,    -9,    85,   -41,    -8,    76,   105,    28,    88,    72,    60,    31,    13,   -54,   -24,   -46,  -107,    24,    51,    14,    25,    55,    11,   -11,     7,    -9,   -12,   -11,    13,    19,     0,   -42,   -46,   -25,    -9,     6,   -19,    45,    40,    34,   -33,   -42,   -24,   -15,   -23,   -26,   -13,    18,    10,    34,   -17,     8,     7,    11,    -1,    -2,    -6,    11,   -16,    -6,     2,   -19,    11,    -4,   -17,    20,    -9,     4,    17,   -23,     6,   -19,   -19,   -29,   -36,   -30,   -30,   -27,    18,     9,     0,    13,   -14),
		     6 => (  -12,    -8,    10,    11,    12,   -18,   -12,   -13,     7,    13,     7,    13,    48,    26,    -4,     4,     6,    -5,   -14,     3,    -3,    10,   -12,    -9,     8,    -9,    13,    -6,    17,    16,   -16,   -18,    11,     5,    33,    40,    72,   101,    86,    38,    91,    63,   -31,     3,    40,    82,     5,    66,    77,    66,    58,    77,    20,    12,   -12,    12,    15,    10,    27,    60,    87,    51,    61,    68,    15,   -13,   -53,    72,   114,    52,    54,   143,    79,    35,    50,   -18,   -25,    -6,    14,    -6,    29,    33,    -7,   -18,    11,    -7,    -3,   176,    97,   -22,    84,   119,   -24,    19,   -53,    32,    32,    79,    38,   -34,   -30,     4,   -67,    -9,    58,    -3,   -12,   -27,   -25,     3,    14,   -19,    -1,    12,   -60,    84,    -7,    46,    48,   -38,     9,     2,    37,    53,   -62,   -11,   -15,   -85,   -50,   -53,   -66,   107,    87,    41,   -50,  -103,   -55,   -60,   -13,    37,   -14,    10,    15,   -31,    -2,  -118,   -91,   -38,   -63,    71,     2,   -54,    43,    62,   -29,   -40,   -95,    24,    32,    58,    25,    -2,   -56,   -89,   -63,   -27,    20,    42,   -15,   -20,    23,   -87,   -81,  -153,  -122,   -20,   -60,     1,   -97,    70,    99,    15,   -14,   -30,   -29,   -77,    32,    -8,   -86,    -9,  -105,  -136,   -28,   -37,    58,   -17,    -5,   -20,     7,   -84,   -74,  -191,  -122,   -59,   -27,   -27,    20,   112,    81,     8,    48,   -64,   -80,   -73,  -190,  -152,  -151,   -86,  -131,  -163,   -98,   -66,    38,   -97,     6,    -5,    20,   -88,   -66,  -208,   -29,   -35,   -92,    53,    26,   -19,    86,    15,   -69,  -139,  -132,  -224,  -203,  -196,  -132,  -149,  -250,  -190,  -161,  -113,   -35,   -87,    15,   -13,   -38,   -54,   -48,  -221,    -9,    16,   -18,   -67,   -55,     8,   -40,   -90,   -85,  -169,  -160,  -229,  -230,  -199,  -121,  -218,  -204,  -146,   -39,   -42,   -51,   -32,   -17,     6,   -28,   -61,  -105,  -199,  -119,     9,    50,     1,   -59,    -6,    46,   -68,  -200,  -185,   -44,    56,    -6,   -98,   -68,   -53,   -95,   -39,   -31,    59,   -72,   -86,    12,     1,    14,  -118,   -87,   -33,   -86,    -1,    66,   -47,   -12,    20,    43,  -159,  -146,   -39,    46,    62,    52,   -59,     0,  -134,   -66,   -93,   -89,   -15,  -119,   -62,    13,   -19,    20,   -67,   -83,   -91,   -48,    77,    50,   -15,   -58,     4,   -56,  -214,   -64,   -13,    83,    32,    -4,    59,    68,   -13,   -47,   -63,    92,   -29,   -71,   -67,     6,     2,   -50,   -37,  -140,  -117,     1,    99,    49,  -122,   -91,     4,   -41,   -92,   -73,     9,   -19,   -21,    -9,    80,   123,    56,   -23,    34,    22,   -33,   -70,    52,     3,     8,   -12,   -93,  -162,   -62,    84,    56,    26,   -31,    35,    95,   -22,   -26,    43,   -20,    38,   -62,    57,    50,    29,    63,    83,    27,   -22,     9,   -46,   -15,     8,    -3,   -22,   -81,  -120,     2,   120,    70,   -21,    -1,   -23,   127,    16,   -59,    83,   -32,     5,   -36,    48,    13,    12,    49,    99,    43,    -1,    31,   -99,  -129,   -19,   -18,   -23,   -66,   -45,    70,   143,   -18,   -25,  -111,    62,   106,   -18,   -70,   104,   -21,   -24,     2,   -19,   -20,    37,    89,    59,    10,    24,    -1,  -124,  -109,    20,    -1,     4,   -44,    -5,   -44,    65,    35,   -60,   -62,    -5,    45,    22,   -21,    15,   -11,   -27,   -65,    32,   -43,   -65,    76,    87,    10,   108,    96,   -49,  -103,    11,     1,    19,   -73,    -1,   -37,    27,    64,    -1,   -87,    11,   -12,    79,    28,    56,   -83,   -33,   -76,   -23,    40,   -24,    97,    35,    75,    66,   129,   -65,  -108,   -16,    -3,   -11,   -73,    55,  -110,   -84,    37,   -13,   -51,   -68,    14,    57,    52,    81,    67,     9,     5,   -56,    28,   -61,   -36,   -83,    69,    29,    87,   -30,    -9,    12,   -25,     2,   -75,    36,   -49,   -82,    -1,  -115,   -47,   -32,    -1,   -43,     9,   110,   118,    26,     9,    85,   -24,   -28,   -33,    35,    63,    86,   108,    -6,    11,    -9,     4,     0,    -8,     7,   -33,    18,    -7,   -97,  -116,   -19,   -81,  -127,   -98,    75,    78,   -27,    32,   -10,    18,    55,   -59,    62,   107,    41,    21,    39,     6,    17,    11,   -16,   -33,   -34,   -43,    54,  -130,  -233,  -233,   -18,   -59,   -70,   -67,   -84,   -48,  -126,   -80,    44,   -85,   -84,   -83,    29,   -40,  -189,  -124,    38,   -15,   -14,   -11,   -18,    -2,   -65,     0,   -60,   -77,   -98,   -45,   115,    30,  -178,  -139,  -158,  -173,  -173,  -211,  -195,   -43,   -51,  -126,  -105,  -151,  -174,   -57,   -56,     3,    12,     7,   -12,   -12,   -18,   -23,   -30,    -9,   -32,   -35,   -64,    -1,   -45,   -98,  -156,  -113,   -69,  -104,  -117,  -192,   -84,   -87,   -39,   -58,   -94,   -65,     6,    -5,     0,    -8,    15,   -14,    -5,    13,   -23,   -31,     8,   -37,   -14,    34,    48,    14,    -3,    -9,     1,   -30,    -5,   -55,   -89,   -65,   -58,   -95,    -8,   -11,     3,     1,   -14,    10,   -10,     6,    -6,   -14,    -9,   -20,   -10,     1,     8,   -24,   -10,   -26,     1,     4,     8,     1,    -9,   -11,   -27,   -22,   -16,     7,    15,    10,    -9,     2,     3,    -5,     3,    18,   -13,    -4,   -20,   -12,     8,     2,     6,    -9,    -6,    16,    -3,    10,    13,    -8,    -7,    14,   -10,     2,   -23,    11,     2,   -10,    10,    -5),
		     7 => (    5,     5,   -14,    -5,    19,   -17,   -18,    19,     3,    14,     5,     6,    -9,   -10,     5,    -7,   -11,     7,    -6,    10,     7,    -3,    15,    18,     0,   -18,    -7,    11,    -3,     7,    -9,     0,     3,   -19,     5,     5,    -9,    15,   -26,   -45,   -17,   -41,   -49,   -50,   -85,   -89,   -55,   -17,    -9,    22,    28,   -13,    18,     3,   -16,     7,    -1,   -17,    11,    -9,   -13,   -18,     4,   -32,   -46,   -15,   -93,  -168,   -79,   -47,   -35,   -25,   -43,   -23,    -1,    -8,   -40,    -9,   -18,    32,     8,   -22,     9,    -6,    14,     3,     3,   -20,    -4,   -63,   -97,   -78,   -94,   -14,   -18,   -62,  -113,  -143,   -74,   -63,   -65,   -32,     0,   -45,   -29,   -21,   -53,   -34,    -7,     3,    20,   -15,    14,    -6,   -17,    -6,   -37,   -40,   -40,  -122,  -161,   -80,  -165,   -46,    19,   -12,   -85,  -129,  -150,  -167,  -113,   -88,   -65,   -51,  -106,  -151,  -105,   -92,   -61,    -1,     4,    -9,    -2,  -125,   -35,    87,   131,    75,   121,    38,   -61,    24,    22,    34,    70,    40,    17,   -24,   -92,  -121,  -198,  -132,  -117,  -179,  -270,  -185,   -51,    19,   -16,    10,   -26,   -87,   -12,    62,    64,    62,    28,    -8,    64,     1,    97,    41,    44,   -50,   -73,   -48,   -92,    -1,     3,   -40,  -104,  -101,  -206,  -108,  -114,   -38,    -9,    51,     1,    28,    26,    60,    29,    -5,    -7,   -65,    15,   -58,    46,   -25,   -66,  -114,   -56,   -68,  -102,   -93,   -20,   -85,    23,    32,   -34,  -119,  -130,   -47,   -58,   113,    58,     8,   102,   132,     0,    64,    17,    40,    20,   -74,   -48,   -35,   -47,    41,    30,    23,   -11,   -16,     7,     3,   -13,   -52,     3,  -173,  -160,   -58,     0,    83,    20,    58,    91,   123,    37,    25,   139,    42,   -68,   -87,   -67,    -6,   -15,    24,   -46,     1,    47,   -19,    43,    43,    50,   -41,   -57,    -5,   121,   164,    14,   -12,    11,   -39,    45,   -16,    65,    84,    74,    -4,    -8,    17,   -50,   -10,   -39,   -22,   -21,    51,    80,    35,    58,    42,    27,   -20,     0,    79,    52,   143,    -1,   -49,    28,    82,    -9,   -35,   103,   152,    98,    77,     8,    -1,     4,    17,    19,   -16,   -48,    94,   -49,    94,    48,   -34,   -58,   -73,   -37,  -117,   -31,   109,     1,    18,    19,   -55,   -92,  -158,    -7,    -7,    17,     4,   -63,   -51,   -49,  -116,   -70,   -17,   -44,   -82,     9,     1,    -6,   -16,   -52,   -34,   -22,    20,    83,   131,   -17,    32,    82,  -101,  -108,  -123,   -43,   -42,   -93,  -118,  -135,  -126,  -194,  -207,   -29,   -18,    -3,   -29,    80,    32,    50,   -32,    25,   117,    48,    50,   -91,   -81,   -31,   -30,   -29,   -89,   -79,  -133,   -93,  -134,  -214,  -169,  -150,  -152,  -179,   -99,    17,    10,    41,   -12,    48,    80,   103,   -52,    18,   -20,   -60,  -147,  -104,   -22,    -3,     2,   -47,   -12,  -145,   -66,   -59,  -181,   -95,   -70,    -8,   -20,    30,    -4,    57,    66,   -37,    37,    25,   -28,   108,    16,    57,   -24,   -37,  -182,   -73,   -32,   -16,   -32,   -36,   -29,   -99,   -88,   -90,  -121,     8,    74,    72,    67,    75,    47,    49,   -68,   -55,    -6,   -20,    25,    -4,    32,    55,   -62,  -204,  -200,   -86,   -54,   -11,   -18,    -6,   -67,   -63,   -79,  -113,  -141,    -3,    19,   -83,    -4,     6,    37,    40,   -66,   -46,   -92,    31,    47,    18,   -28,    34,   -49,   -80,    14,   -20,   -39,    25,   -23,    95,   -49,   -95,  -157,  -173,  -111,   -68,  -183,  -121,   -21,    95,   103,   -96,   -95,   -73,   -29,   -19,   -82,   -62,   -92,   -46,   -84,   -74,   -42,    65,   -32,   -12,    36,    15,   -30,   -77,  -194,  -102,  -112,   -91,    29,   -58,   -53,    -5,   -25,   -62,   -52,   -19,   -94,   -59,   -40,   -49,   -85,   -70,   -91,  -156,   -19,   -81,     0,    15,   -24,     4,   -38,  -107,   -20,    12,    50,   -41,   -23,   -20,   -14,    23,    26,   -88,  -108,   -85,  -138,  -135,  -102,   -38,     7,    35,    -6,   -69,   -32,  -129,   -13,   -24,   -20,    -7,  -111,   -79,    84,    98,   -54,    31,     0,   -27,   -61,   -30,    31,  -194,  -129,  -176,  -188,  -111,  -123,   -99,   -15,   -25,   -91,   -75,   -21,   -33,   -27,   -45,   -34,   -29,  -172,    58,    90,    85,   103,   127,    37,    37,     3,   -44,   -76,  -125,  -120,  -130,  -103,  -144,  -104,  -110,    13,    30,  -189,  -109,   -13,   -39,     4,     0,    15,   -48,  -198,    50,   -11,    65,   167,    11,     3,   -27,    44,   -64,   -44,  -121,   -56,  -137,  -227,  -178,  -163,  -155,   -13,     3,   -85,   -64,    -8,   -93,     2,   -19,    -1,    40,   -11,    81,   122,    84,    29,   102,    18,   -39,    31,   -30,    40,   -72,   -57,  -195,  -200,  -165,  -102,  -140,    10,   -38,  -149,   -21,   -56,   -15,    16,   -17,    -5,   -34,    75,   -81,    15,    -4,    36,   -44,   -90,   -16,    51,   -21,  -108,  -140,  -108,  -129,   -74,   -47,   -70,  -178,   -16,   -26,  -115,    21,     2,   -22,   -18,    19,    10,    -9,   -89,  -104,  -114,   -28,    56,    96,    36,   -53,    -3,    30,    62,   -70,   -24,    -6,   -40,    20,    -7,   -53,    54,    78,    35,   -29,     3,    14,   -16,    -1,    -6,     1,    15,    83,    77,   -17,    -9,   -21,     1,    52,    38,   -37,   116,    77,     6,    30,    15,    18,   -17,    23,    93,    69,    82,    -5,    13,     2,     5),
		     8 => (   -9,     7,     3,     7,    -8,    12,   -13,     2,    16,   -10,    -5,    16,    -4,    -3,    -3,   -13,   -16,   -13,    -9,    -7,   -18,   -12,   -11,   -14,     0,    -1,    -6,    11,    11,   -11,   -11,    13,     6,    16,    17,   -17,    14,    19,     3,     6,    -3,   -24,   -16,   -21,   -56,   -47,   -25,    12,   -11,     1,    12,     9,     0,    16,    14,    -8,     8,   -15,   -16,    15,   -19,    16,    -7,    -6,   -20,   -57,  -145,  -126,   -34,   -32,   -20,   -60,   -80,    61,    94,    32,   -61,   -60,   -57,   -59,   -21,   -29,    17,    -3,    -6,   -19,   -44,   -40,   -34,   -58,   -35,  -113,    79,    60,   -34,   -92,   -84,   -62,   -60,    24,    18,    16,   128,    63,     1,   -44,    83,   113,    -3,   -27,   -40,    18,     3,   -12,   -41,   -60,  -109,  -146,    -1,    60,   -14,   -87,   -77,    46,   -26,    -5,    24,    29,    37,    11,   -19,     4,   -46,     1,    46,   -51,   -88,    67,    77,    -2,   -10,   -11,   -30,   -63,   -65,  -108,     4,    -7,  -108,   -59,   -37,     0,   -12,    42,   -10,    32,   -38,  -110,  -134,    78,   -15,    78,     7,   -36,   -38,   -10,   -37,   -29,    11,     1,   -63,  -113,   -81,    14,   -16,   -50,   -89,   -40,    19,   -42,   -35,   -38,   -95,     1,   -57,   -57,   -59,    36,     5,   -32,   -30,   -83,   -75,   -54,   -12,   -10,    13,   -88,   -26,   -42,    -8,   -10,   -42,   -43,   -10,   -16,   -68,   -16,   -49,  -109,   -64,    28,   -21,   -78,   -55,    13,     6,   -19,   -80,   -66,   -68,    -6,    24,    56,   -38,   -66,   -19,   -13,   -45,    -7,   -76,   -33,    13,    37,   -96,   -74,   -49,   -14,   -41,   -39,   -65,   -86,   -50,    11,    18,    31,  -106,  -120,   -37,     8,   122,    60,    -7,   -26,   -64,     8,   -31,   -33,   -63,    27,    -4,   -41,   -98,   -11,   -34,   -62,   -92,   -85,   -45,   -46,   -98,    46,    19,  -106,  -114,   -98,   -82,    -5,    41,   -61,    17,   -28,   -55,     0,   -26,    19,   -55,   -54,   -15,     4,    44,   124,   -38,   -50,    29,    11,    11,    10,    31,    53,     5,   -38,   -80,  -124,   -55,   -72,    16,    26,    -2,   -24,   -26,   -61,   -42,    50,    31,     0,    30,    76,    42,    13,   -49,   -86,   -34,   -24,    39,   -20,     7,   -73,   -81,    81,   -52,   -53,   -26,  -159,    -9,   -79,   -11,     5,   -58,    -3,    58,    78,    51,   -16,    22,    69,    53,   -74,   -45,   -82,   -67,   -88,   -50,   -35,    -2,   -86,   -10,    42,    46,    70,    23,  -137,  -143,  -109,    19,    -9,   -74,  -117,    15,    43,   -29,  -106,    53,   158,    60,    47,   -17,   -53,   -74,    -7,     8,  -125,   -37,     4,    40,    97,    71,    72,   -11,  -122,  -189,    24,     0,     5,    -4,  -142,   -66,   -22,   -42,  -116,    23,    18,   -15,     2,    20,    -7,   -49,   -46,  -170,   -74,    56,    82,    82,    66,   -35,  -108,  -153,  -115,  -181,     2,   -20,     6,   -32,    38,    17,   -73,   -59,   -53,     7,   -12,    44,    68,    -7,    -9,   -63,  -139,   -51,   -28,   -56,    21,   -24,   -96,  -113,   -58,   -44,     1,   -92,   -72,     8,   -10,   -16,    72,   -12,   -61,   -70,   -65,  -159,  -107,   -32,    40,    50,   -57,   -41,   -35,    -6,   -18,   -10,   -60,   -15,    23,   -55,   -18,    11,   -18,  -103,   -56,     8,   -11,   -37,    53,   -48,   -69,   -88,   -49,  -139,  -251,   -97,    25,    75,   -13,   -11,    13,    15,   -42,  -103,   -95,    16,   -43,   -47,   -45,   -39,   -20,    13,   -30,   -22,     8,   -45,   -52,   -30,   -56,   -74,   -75,   -48,   -85,    -5,    -6,    41,    28,   -43,    51,    38,   -31,   -27,   -33,     7,   -59,   -31,   -62,   -26,   -11,   -17,   -46,    11,    -9,   -36,   -29,   -17,   -49,  -100,  -121,    34,    39,    -5,   -28,    50,    31,   -23,    69,   -58,   -14,     0,     4,   -70,   -59,   -48,   -42,     1,    -4,   -62,   -69,    16,   -10,   -29,    -1,   -43,   -35,  -116,  -128,   -29,    32,   -24,   -26,   -22,    40,   -56,    11,   -89,   -91,   -31,    -7,  -120,   -47,   -12,     6,     2,    -2,   -45,    -2,   -34,   -16,   -38,    -3,   -51,   -64,   -93,   -20,   -73,   -66,   -39,    31,   106,    32,    38,    17,   -47,   -46,   -33,   -38,   -67,   -54,   -33,   -30,   -48,   -23,   -58,   -20,   -33,   -46,   -20,   -30,   -42,  -126,  -143,   -79,   -52,   -50,  -115,   -54,    60,    45,    48,   -76,    -9,     5,    -3,     4,   -31,     2,    -3,    -6,   -30,   -21,   -55,    -5,   -13,     2,   -49,   -14,   -15,   -67,  -122,  -160,   -53,   -10,   -58,    -4,   -57,   -24,   -82,   -34,    16,   -56,   -47,     4,    38,    39,    11,   -24,     2,    -4,   -63,    -3,    19,   -10,    -9,   -14,   -27,   -45,   -44,   -76,   -59,   -55,  -141,   -46,   -60,   -64,   -32,    51,    41,   -42,    69,    38,     5,   -11,   -29,   -32,  -108,   -76,   -28,    16,    -7,    15,   -28,   -10,   -26,   -70,   -49,   -26,   -48,   -52,   -79,  -101,   -16,    28,   -23,    46,   -11,   -12,    43,    40,    15,   -79,   -28,   -31,    -3,   -32,   -12,    10,     6,   -10,    -9,   -28,   -22,   -48,   -75,   -26,   -22,   -37,   -58,  -123,  -147,  -118,  -123,  -180,     3,   -16,   -19,  -150,  -135,   -77,   -53,    20,   -18,   -10,    18,   -13,     4,    -8,   -13,     6,   -29,    -9,   -25,   -13,    -3,   -37,    -9,   -43,    12,   -39,    -2,    -3,     1,    10,    -3,    -7,    -4,     8,   -19,   -10,     9,    17,    -7,    10),
		     9 => (   -5,   -11,    13,   -12,    -9,   -18,   -12,    16,    11,     3,   -16,    -2,     4,    -1,    19,    20,    -9,    -2,   -20,    11,    -2,   -13,    10,     9,    19,   -20,    -5,     2,    20,   -10,    17,    14,   -15,    11,   -22,   -10,    17,    -4,    -9,   -11,   -54,   -30,    -7,    -4,   -20,   -19,   -36,    15,     1,   -27,   -13,   -21,    -3,    -6,    -8,    -8,    -2,     2,    13,   -11,     9,    17,    -2,    -2,   -14,   -22,   -27,    -3,    -5,    -9,   -55,    -9,   -24,    -8,   -18,    -4,   -50,    23,   -20,   -24,   -20,    18,     0,   -10,    -2,     0,    12,   -34,    -4,   -32,   -23,    -4,   -64,   -28,   -40,   -88,   -55,   -20,   -47,   -49,   -55,   -25,    50,   -29,   -50,   -67,   -53,     4,   -29,   -22,     3,   -10,     0,   -17,    -1,   -32,   -30,     9,   -86,   -22,   -24,    -9,   -36,   -44,  -119,  -156,  -177,  -171,   -91,   -11,    62,   -85,  -129,   -91,   -65,   -57,   -51,  -113,   -81,     8,    -2,    11,   -17,   -26,     6,   -18,   -36,   -45,  -114,   -65,   -99,   -30,   -32,    37,   -43,   -68,  -141,  -150,  -144,  -123,    17,   -64,   -82,   -95,   -60,   -53,  -126,     9,   -19,   -25,     1,   -29,    33,   -53,   -19,  -122,   -96,   -94,  -126,   -46,   -57,   -93,   -31,   -36,   -36,   -92,     5,   -63,    29,    57,     2,   -38,   -56,   -67,   -86,   -79,    -8,   -30,   -47,   -42,   -64,  -107,  -114,  -139,  -161,  -222,  -181,  -142,   -68,   -57,   -72,  -135,    42,    27,   -11,   -17,   167,    64,    63,    46,   -28,   -81,   -32,   -52,   -65,   -22,    17,     0,   -78,   -61,   -75,  -103,  -121,  -173,   -56,  -113,   -49,   -23,  -108,   -42,    14,    63,    65,     7,    11,   -11,    -7,    70,    27,   -50,   -74,   -38,   -15,   -37,    97,    -9,   -42,   -70,   -41,   -17,  -133,   -25,   -28,   -45,   -56,  -106,    20,    82,    15,     6,   -19,    54,   -68,    13,    31,    -2,    57,    53,  -160,   -76,     0,   -25,   -66,   -56,    -9,   -47,   -89,  -112,   -42,    -5,   -17,    35,   -49,    34,   -20,   -75,   -76,   -62,  -146,  -131,   -65,   -27,   -51,   -14,    90,   192,   -67,  -117,    18,  -162,   -35,   -26,   -44,   -73,   -67,   -21,    93,    49,    64,   -23,    19,   -30,   -84,  -143,  -159,  -183,   -83,   -33,    49,   -18,    45,    20,   135,   180,   -14,  -102,     8,   -16,    14,   -96,    42,   -46,   -84,    -8,    42,    22,    73,   -36,  -108,   -77,  -135,   -95,   -42,  -141,     0,    -3,    87,   -26,    58,    72,   -27,  -137,  -118,  -116,   -15,   -30,   -42,   -69,    45,   -61,    -7,    28,    15,    46,   103,     9,     9,    19,   -61,    53,   100,     6,    -4,   108,    38,   114,    18,   -41,   -92,   -60,   -65,     8,     2,   -30,     7,   -64,    52,   -56,    -6,   -46,   102,   105,    93,     0,    43,    49,    41,    63,    10,    14,    -6,    50,   -32,  -115,   -45,  -142,  -130,   -27,    17,     4,   -12,    14,  -117,   -76,    54,   -59,   -83,   -67,    20,   -51,    15,    48,    51,   111,     4,    30,   -13,     4,    63,    27,   -93,  -112,  -154,  -119,   -97,   -21,   103,   -20,   -22,   -30,   -76,   -67,    37,   -39,   -13,    -5,   -54,   -26,    26,    38,   -37,    20,   -77,   -89,     2,    44,    21,   -11,  -135,   -48,   -44,  -143,   -70,    -6,   -17,    -8,     9,   -22,   -63,   -18,   -53,   -61,   -41,    58,   -56,   -98,   -69,   -51,   -36,   -19,   -49,   -23,    -4,    71,    54,   -55,   -70,   -33,   -71,  -143,   -60,    79,    -8,   -30,    -2,    13,   -66,   -28,  -133,   -97,    -1,    51,   -64,  -106,   -23,    28,   -40,   -24,    44,   -51,   -13,   -31,    32,     7,   -62,   -49,   -11,   -54,   -33,    94,   -54,   -53,    -4,   -17,   -74,   -49,  -141,  -119,   -53,   -45,   -87,  -130,   -82,  -106,   -12,   -57,   -11,   -68,   -77,   -50,   -22,     5,  -133,   -61,   -10,   -26,    30,   109,   -71,   -50,    12,    -1,    49,   -40,  -102,   -60,  -178,  -138,    42,   -53,  -119,   -19,    67,    49,   -25,   -79,   -26,    -9,     4,   -28,   -75,   -67,   -50,   -13,    26,    94,   -20,   -14,    -5,   -15,   -17,   -51,  -108,   -52,  -125,   -92,    31,    43,     7,   -46,   -23,   -58,   -48,  -150,     6,   -36,   -34,    28,   -71,   -55,   -74,   -32,    21,    78,   -79,    -8,    14,    12,   -64,  -103,  -126,  -102,  -162,   -54,    33,    53,    59,    42,   -22,   -68,  -108,   -79,   -47,   -31,  -115,     3,    17,   -67,   -35,     5,    31,    -9,   -44,   -16,     1,    12,   -58,   -74,  -159,   -78,  -102,    17,    89,    65,    19,   -66,   -20,  -100,  -101,   -26,     7,   -15,   -22,   -20,    22,    -5,    12,   -63,   -22,    32,   -40,    15,    13,    15,   -33,   -55,   -73,     1,     7,    49,    20,    64,    22,   -23,     1,  -102,    19,   -71,   -63,    -2,   -54,    37,     8,    -3,    33,     2,   -12,   -10,   -27,    -2,   -20,    17,    63,   -28,    28,   -12,   -33,    -6,    39,    22,    65,    -7,    55,    -3,   -60,   -57,    18,    81,    51,    14,   -28,   -40,   -50,    44,    11,    -9,    -9,     7,    16,    20,     1,   107,    50,   -20,    61,    53,   -42,     5,    32,    97,    16,    78,    62,    35,   110,   139,    74,    52,   104,    17,   -43,    30,   -23,     4,     7,   -17,   -12,    11,    18,   -10,   -31,   -21,    28,   109,    95,    67,    63,   134,    70,    60,    50,    50,    25,    49,    78,   102,   -38,   -48,   -25,   -27,    20,    -5,   -19,    -6),
		    10 => (   10,    16,     6,   -19,     8,    -7,   -16,     3,    15,   -10,     7,    -4,   -17,     3,     1,     4,     6,    -9,   -15,    -9,     3,    -9,     0,    10,   -17,    -2,     0,    11,    -2,   -18,   -14,   -17,    11,    19,    -8,     9,    18,   -22,   -21,    20,    46,     6,   -33,    65,    82,    90,     2,    13,    13,    -1,     1,   -10,    -4,     1,   -10,    11,    18,    19,   -24,    75,    67,   -20,   -18,    15,   -26,   -33,   -59,    -7,    -1,   -43,   -22,   -93,   -12,  -110,   -92,   -99,   -80,   -29,   -93,   -56,   -44,   -13,   -19,    19,    18,    10,    10,    -4,   -22,    -2,   -25,    -6,    37,   -61,  -156,   -93,     7,    21,   -14,   -78,   -64,  -127,   -14,    -3,     9,   -74,   -77,   -42,    -8,    15,  -139,    -1,    15,    14,   -20,   -29,    21,  -102,   -67,   -83,   -56,  -104,  -110,   -90,  -159,  -167,   -34,    31,   -80,    22,   -37,     1,   -13,     5,    31,    23,   -71,  -109,  -117,   -14,   -14,   -19,   -46,   -16,    16,  -119,   -59,  -119,   -37,    -2,  -140,   -58,  -102,   -66,    -9,   -19,   -50,    -4,   -49,   -12,  -139,   -65,    69,     6,  -113,   -74,   -96,   -72,     5,     9,   -81,   -11,   -22,   -11,   -50,   -50,    17,   -14,   -44,     7,   -40,     7,     4,   -45,   -31,     0,    18,    10,   -64,    48,    88,   -51,  -113,  -112,    -6,   -15,    -1,   -96,   -52,   -31,   -20,     9,   -15,   -81,   -13,   -39,   -13,    15,   -15,   -41,   -33,    17,   -54,    13,    55,    21,  -111,    -6,   -37,   -50,  -160,  -115,   -80,    44,   172,  -135,    69,    32,   -22,   -30,   -26,   -93,   -49,   -46,     1,    -6,    27,  -156,    24,    67,    -1,    90,    62,   -80,  -112,   -25,   -50,   -52,  -161,   -64,  -121,   -19,    12,   -28,   103,   -12,   -22,    23,   -62,    19,    35,   -37,    18,   -11,     3,     0,   -43,   -51,    68,    34,    57,   -26,    60,   -30,   -71,   -71,   -67,  -148,  -129,    -1,    -5,     8,    61,    33,   -14,    -9,   -20,   -32,   -28,   -13,    23,   -10,    -3,   -31,    16,  -133,   -46,    46,    -8,    -4,   -31,   -68,     8,   -19,   -96,   -89,  -105,    -9,   -13,   203,   -68,   -70,   -78,    17,    31,   -64,  -131,  -111,   -15,    11,   -28,    30,   -85,  -146,  -115,   -22,    36,    53,    -8,  -119,  -125,   -92,  -124,  -118,   -71,    10,     3,    28,   -33,   -88,    76,    84,    21,   -50,  -182,   -19,    31,    14,    67,    -8,  -115,  -155,   -65,    12,    68,    89,    27,   -96,  -116,   -46,   -97,  -123,   -46,   -17,   -13,    47,    55,   -73,   147,    71,    44,    10,   -67,    58,    30,   -18,    10,   -80,  -193,  -261,   -99,     7,    22,    94,   131,   -83,   -45,    52,    12,    -8,   -77,   -30,    14,    11,   -20,   -99,     6,    86,   -68,    18,    47,    50,    23,   108,    86,   -22,  -139,  -107,   -86,   -64,    51,   131,   115,   -88,    -2,    77,    -8,   -46,   -43,   -25,    15,   -14,   -68,  -120,   -78,   -47,   -47,   -18,    40,    15,    51,    94,   194,   -74,  -196,  -100,   -36,    -7,   106,   -24,    46,  -107,    -9,    47,   -27,   -30,  -159,   -29,    16,     9,   -57,   -72,   -54,   -21,   -80,   -84,    59,   -17,   -31,    46,    58,  -142,  -206,   -20,    33,    39,    44,    38,   -83,  -139,   -94,   -29,   -66,   -91,  -135,   128,    12,   -30,   -66,   -88,   -20,   -58,  -109,   -35,    22,   -28,     4,    -2,    29,  -116,  -112,   -13,    39,    33,   -34,    33,   -12,  -134,   -54,   -62,   -64,   -80,   -79,   200,    -5,   -28,   -74,   -73,   -69,  -140,   -88,   -47,     6,   -25,    32,    16,   -81,  -100,   -68,     7,   102,    31,    19,   -45,   -66,   -83,    -1,   -67,   -35,   -59,   -97,   -47,     4,    58,     0,   -54,   -78,   -83,  -121,   -48,    75,    14,    -5,    17,   -16,    19,   -42,   -35,   -95,   -51,    65,   -34,   -34,     6,   -61,   -70,    -9,  -107,   -61,   -22,   -20,    71,   -28,   -66,   -20,   -80,  -141,   -62,    28,    14,    52,    58,    71,    43,   -13,  -126,   -93,   -20,   -64,     7,   -37,    28,   -72,   -22,   -84,     8,    48,    14,    15,     6,   -38,   -86,   -99,   -49,   -88,   -59,     5,    20,   106,    10,    94,    41,   -63,   -60,   -53,   -53,    13,    49,     3,   -43,   -76,   -14,    -1,    22,   249,    58,    14,   -19,   -80,  -133,  -109,   -58,  -100,   -75,   -41,    67,    -6,    -4,     5,  -106,    24,    48,    51,   -62,  -114,   -21,  -103,   -84,   -59,   -37,   -11,    40,   137,    55,   -19,    11,    -8,   -87,  -103,  -167,   -70,   -56,   -64,    73,   138,    45,    26,   -25,   -12,   -68,    12,   -42,     0,   -22,  -103,   -82,   -24,   -27,     0,     4,  -112,     2,   -10,    -4,   -31,    -1,    54,    37,  -108,  -139,  -150,  -113,   -99,   -59,   -16,   -72,   -96,   -58,   -70,   -30,    49,  -127,   -78,   -69,   -47,   -16,    16,    23,    12,    10,    20,    -4,   -25,     0,   -77,   -66,   -73,  -113,   -31,   -57,  -145,  -169,  -281,  -271,  -281,  -218,  -127,  -105,  -106,  -102,  -127,  -102,   -56,   -47,     5,    -6,    -8,     8,    19,   -18,     9,    14,   -51,   -74,  -180,   -54,   -71,  -138,   -91,  -103,   -71,   -75,   -28,   -99,   -95,  -100,  -133,  -116,  -102,   -84,   -40,   -44,     2,     9,     9,     7,    -6,   -15,   -18,    18,    -8,    12,   -17,   -33,   -41,     2,    -9,    -7,    -1,   -21,   -25,   -26,   -14,     0,   -18,    -4,     9,   -22,    -4,   -21,     8,   -13,   -13,     4),
		    11 => (    3,     4,   -15,   -19,    16,   -18,    19,    12,    -2,    10,    18,   -19,   -12,   -14,    15,   -17,     5,    14,   -10,    -4,     2,   -14,     6,   -15,    14,    -4,    17,   -14,     3,    -5,   -15,    20,    -1,   -18,     2,     9,    19,     1,     2,   -20,   -10,   -36,     2,   -27,   -38,   -32,    -3,   -16,     4,   -15,   -11,    14,   -13,    17,    -9,   -14,   -17,   -19,   -15,   -18,   -17,     2,    14,     6,   -33,   -15,    27,    18,     4,   -14,   -22,   -65,  -148,  -178,  -143,    37,    47,   -61,   -27,   -48,   -18,   -17,     4,     5,    11,   -20,    53,     9,   -10,   -17,   -20,    66,    60,    81,    64,    16,    13,    -2,    17,   -92,  -149,  -112,   -15,   -51,   -48,   -81,    22,    61,   -58,     0,    -2,    17,    -9,    14,    46,    41,    18,    40,    58,    51,   -19,     4,   -56,   -46,   -41,   -54,   -60,  -118,   -90,   -44,    16,    36,    79,    -1,    -1,   -32,   -93,   -70,  -102,   -85,    -6,   -10,     4,    87,    67,    68,   -14,     4,  -104,   -58,   -86,   -95,   -41,   -30,  -178,  -193,  -125,    14,    37,    20,    -4,    77,    64,    27,    16,   -62,   -74,    -6,    -5,    -2,   -13,    78,   138,   -23,   -52,   -10,  -116,    73,    57,    -6,  -177,  -202,  -256,  -209,  -100,   -65,    -2,   -21,   -24,    15,    -1,    14,   -54,   -84,   -59,   -39,    10,   -30,   -48,     4,   -59,   -68,   -52,   -65,  -133,     0,    84,     6,  -111,  -161,  -178,  -140,   -46,   -26,    51,     0,     9,   -12,   -12,    23,  -113,  -166,  -101,   -28,    -1,   -71,   -56,   -16,   -29,   -40,   -40,   -81,   -81,   -29,    10,  -110,   -87,   -99,  -175,   -86,    -2,    37,    23,    -5,    37,   -25,    -5,   -11,  -112,  -135,  -103,   -31,   -10,     6,   -52,   -20,   -30,   -45,   -35,   -38,   -38,    -7,  -146,  -163,  -173,  -280,  -247,    -1,    65,    12,    28,   -14,   -20,   -26,     6,    -6,   -27,   -82,   -30,   -59,   -13,     8,   -26,    -9,     0,    -1,   -90,   -94,  -131,   -80,  -146,  -143,  -192,  -235,  -116,    -9,   108,    18,   -36,   -13,    -4,    32,    24,    -8,    18,   -40,   -48,   -37,   -17,     8,    24,    12,   -27,    17,   -40,  -107,  -120,   -95,  -123,   -76,  -114,   -85,   -56,   127,    48,    44,   130,   -26,    -4,    12,   -73,  -107,   -68,    10,   -60,    10,    -9,     4,   -57,    31,    -3,    38,    13,   -86,     9,  -143,   -91,   -99,   -35,   -61,    36,    96,     6,    49,    17,    32,   -96,    -6,   -80,   -17,   -55,     8,   -29,     2,   -16,     6,   -44,    -1,     4,   -46,   -24,   -48,   -38,   -81,   -36,   -20,   -66,    15,    95,    61,    16,    60,    42,   -42,  -219,   -95,   -95,   -33,   -42,   -22,    -2,     5,   -11,    -6,    -7,     0,    25,   -31,   -25,     1,   -14,    59,    71,   -27,    -6,    66,    26,    31,    54,   -87,  -119,  -255,  -279,   -35,    38,    -3,   -21,   -48,   -29,   -12,     4,   -20,    50,    94,    -6,  -105,    -5,    16,   139,    55,    45,     9,   -20,    18,    16,    47,    16,   -79,  -230,  -286,  -168,   -26,    27,     4,  -182,  -136,   -86,    -1,    14,    -1,    19,   -28,    29,   -25,   -60,     4,    56,    52,   -83,    -8,   -29,    -5,   -68,    43,    44,   -18,  -163,  -154,   -22,    43,    52,   107,   151,   -59,   -94,   -26,     0,    -1,    -5,   -52,    -1,  -116,   -52,    30,    -3,     4,   -22,    63,    55,    -7,    13,   -76,    19,    -9,    27,    61,    76,   134,   169,   158,   119,    -9,  -170,   -63,     3,    -2,   -12,    -5,   -73,  -191,  -118,    16,    10,    -9,   -24,    54,   -25,   -13,     6,   -23,   -58,    -7,    29,    46,    46,    -9,    98,    77,     1,    31,   -10,    49,    -7,    15,    14,   -69,  -116,   -34,     9,    30,    22,   -13,   -38,   -15,   -12,   -75,  -153,  -114,   -76,  -111,   -89,   -56,   -48,   -30,    58,    78,    75,    82,    -5,    25,    -8,    -7,    -1,   -56,    28,    61,    53,    11,    25,     3,   -43,    48,   -54,  -109,  -113,   -78,    38,   -53,  -117,   -72,   -77,   -26,    64,    60,   111,    -1,    17,    30,    43,    48,     7,     2,   -17,     1,   -10,    20,    14,   -31,   -32,   -12,   -40,   -20,   -36,    23,    59,    44,   -63,   -55,   -80,   -36,    19,   114,    93,    43,    13,    16,    60,    46,     5,     6,    24,   105,    31,    -4,    27,    61,   -35,   -55,   -87,    -8,   -74,    66,    82,    -1,   -67,   -86,   -78,   -79,    11,    15,    21,     3,    21,     6,     2,     2,   -28,    51,     8,     7,     8,     4,    86,    49,   -28,   -76,    17,    33,    40,    70,    26,   -44,   -56,   -69,   -32,    -7,   -12,   -18,    53,   101,   122,     9,    -4,     6,    13,    33,   -93,   -67,   -94,  -124,   -24,    75,   -18,   -55,    70,   112,    12,    12,    -8,     4,     0,   -31,    -2,    14,    19,    13,   -61,    15,     2,    12,    -3,    -8,    17,   -43,   -78,   -78,   -26,  -166,   -41,    33,   -33,    26,    85,    24,  -121,   -74,   -62,  -109,   -63,   -39,   -22,   -60,   -46,   -38,   -42,   -12,     0,   -10,    -5,   -18,    -6,   -11,   -74,   -57,   -60,   -88,  -114,   -94,   -65,   -32,   -60,   -60,   -49,   -53,   -74,   -81,   -32,     4,   -11,   -12,    -8,   -11,     9,    -3,   -17,   -15,    11,     0,   -19,    10,    -7,   -10,     4,     7,     9,   -13,   -62,   -28,   -16,    -9,   -37,   -20,    16,     7,   -19,     1,    -1,    -1,    14,   -12,    -9,   -10,   -16,    17),
		    12 => (   19,   -17,    18,   -13,     3,    -5,    -5,    19,     6,    12,   -15,    13,    11,   -16,    35,    19,   -20,   -12,     8,    -7,     5,     7,   -12,   -13,     6,     5,    11,   -10,   -19,   -15,   -13,   -11,     1,     1,     3,   -29,   -63,   -24,   -27,   -35,   -32,   -54,   -17,    15,    20,    -7,   -20,   -63,   -40,   -34,    -6,    19,    -3,     8,   -20,    -7,    16,    -6,   -25,   -59,   -42,    15,    -6,   -21,     5,    14,    22,    65,    21,   -31,   -26,   -58,   -69,   -41,    21,    22,    10,    12,   -54,   -19,   -32,    14,    14,    13,     1,    19,   -23,  -115,     5,   -59,   -29,   -56,    -7,    60,   114,    83,    64,    14,     5,     9,    -3,    -3,   -31,     1,    12,    20,   -56,  -100,   -51,   -47,   -14,     8,     0,    -6,    -7,   -45,    13,    34,    72,   100,     8,    -3,    29,    90,    83,    99,     2,   -15,    -4,   -45,   -11,   -68,   -36,   -56,   -65,   -61,  -107,   -88,   -87,   -18,    19,    14,   -69,    -9,     5,    39,    74,   135,    66,    33,    30,     8,    23,    22,   -43,   -31,   -49,   -34,   -44,   -21,     8,    19,   -27,   -53,   -92,   -41,   -49,   -18,   -20,   -12,     1,     0,   -11,     5,    97,    79,    52,    50,    18,     5,   -25,    -3,   -32,   -44,   -33,   -30,   -12,   -56,    -9,    25,    14,   -60,     1,    88,   -46,     5,    14,   -16,    -9,    -8,   -24,    18,     5,    26,    -2,   -50,   -38,    -1,   -29,   -42,   -23,    20,    23,   -63,   -57,   -72,     9,    40,   -23,   -63,    28,   105,  -136,   -57,   -58,    39,   -25,     4,   -16,     4,   -23,    13,   -67,   -83,   -41,   -47,   -12,     8,    -5,    11,    16,   -21,   -47,   -23,   -15,    -6,   -21,    25,    15,   -11,  -127,   -63,    11,   -55,    66,     1,   -30,   -23,   -43,   -34,   -57,   -74,   -38,   -49,    -7,   -20,    70,    14,   -50,   -18,   -40,   -31,   -10,    24,    22,    -4,   -36,   -71,     0,   -46,    13,    -9,    20,   -18,   -65,   -26,   -47,   -83,  -121,  -104,  -117,   -42,   -14,   -34,   -30,     3,   -71,   -21,   -78,   -20,   -67,    25,    40,   -38,   -78,   -31,    37,   -71,    -8,   -41,   -23,   -67,   -52,   -39,     3,  -112,  -119,  -119,  -110,   -38,   -10,    13,    32,   -28,   -81,   -51,    23,   -10,   -34,   -33,   -21,   -30,   -55,   -27,    -2,   -30,    -9,   -27,   -71,   -78,   -31,   -14,   -52,   -63,   -27,   -31,   -29,    17,    56,    -2,   -11,   -19,   -43,   -25,   -43,     6,   -72,   -79,   -30,   -67,   -85,     5,    33,    17,    13,   -26,   -42,   -51,   -55,   -84,   -30,   -74,   -50,   -21,     1,   -16,    -4,   -11,   -14,   -24,   -53,   -44,    21,     0,   -29,   -29,   -58,   -68,   -20,    24,    67,     3,    -4,   -48,   -35,   -21,   -61,   -91,   -18,   -59,   -42,   -48,   -42,   -71,   -68,   -43,   -38,   -56,   -70,   -76,     6,   -19,   -16,   -87,   -65,   -59,   -20,    50,    85,    51,     3,   -59,   -39,     5,   -49,     8,   -46,   -33,    -4,   -51,   -26,   -39,   -58,    -8,   -19,   -60,  -113,   -82,    -6,    -3,     7,   -35,   -60,   -74,    33,    79,   104,    77,     7,   -30,   -13,    58,    52,    -2,   -29,   -38,   -23,   -19,    20,     6,    20,    21,    13,   -40,   -61,   -58,   -67,   -45,   -31,   -24,   -47,   -60,     8,    63,   125,    82,   -18,   -18,    19,    62,    54,   -16,    -8,   -70,   -31,   -21,   -35,   -34,    54,    12,   -34,   -37,   -76,   -72,   -45,   -71,   -85,   -51,   -52,   -92,     0,   100,    82,    96,    17,     1,   -20,    17,    65,     1,   -66,   -28,     1,    12,    -9,   -54,    -3,   -15,    -3,   -13,   -84,   -35,   -69,   -59,   -29,   -33,     8,    -3,    61,    58,    63,    75,     4,    -6,    -4,    27,    14,   -34,   -10,   -28,   -12,   -33,    13,    22,     4,     7,   -47,   -37,    -8,   -23,    42,   -98,   -40,    27,    49,    73,    74,    79,   137,   148,     6,   -28,    14,    -9,    30,    28,   -22,   -24,   -36,    -4,     7,    49,    -4,   -28,   -41,   -51,   -24,   -38,    38,   -64,   -13,    38,    60,    82,    92,    50,    43,   -16,    10,     8,    32,    42,   -26,    14,    -6,   -44,   -59,   -47,   -44,   -17,   -44,   -30,   -52,   -30,   -10,    13,   -21,   -40,    22,    46,    89,    84,    42,   -11,    15,   -29,    -1,    10,     8,    24,    43,   -29,   -14,   -36,   -15,   -31,   -59,   -32,   -20,   -21,    27,   -38,    30,   -28,   -49,    -2,    10,    34,    80,    75,    21,    59,   -65,   -33,    -3,     8,     9,    22,    18,     0,   -13,    -2,    29,   -40,   -22,    40,     4,    15,    25,    22,     2,   -58,   -76,   -55,    11,    34,    83,   100,     3,    46,   -33,    12,    -8,    18,   -42,   -20,   -41,   -45,   -44,    -7,   -22,   -15,   -54,     3,    41,     2,    50,    -2,   -58,   -39,   -41,    -3,   -49,   -20,   -52,    37,    26,    14,     4,    -4,   -14,     8,   -72,   -18,   -10,   -13,     3,   -13,   -49,   -65,   -70,   -23,   -60,  -110,   -42,   -50,   -77,   -13,   -52,    -3,   -53,   -49,   -57,   -38,   -27,   -11,     4,    15,     1,    18,     2,     9,   -35,   -63,   -43,   -49,   -60,   -89,   -80,   -38,   -30,   -53,  -102,   -77,  -160,  -171,  -147,  -119,   -63,   -46,   -80,   -54,     5,    -6,    20,   -20,    11,     7,    10,    -6,    -2,    12,   -23,   -29,   -44,   -24,   -47,   -56,   -28,   -88,   -55,   -52,   -59,   -51,   -69,   -25,   -43,   -30,   -46,    15,     4,    -8,   -19,    18),
		    13 => (   -9,   -20,    18,    -9,   -15,     6,   -20,   -18,    18,     8,    15,   -13,   -20,   -20,    -6,     0,    14,    19,    -6,     7,    18,     9,    -9,   -19,    10,    -5,    -6,     7,     9,     5,   -13,    14,     4,    -9,   -15,    -5,    17,    -1,   -11,     9,    -1,   -10,   -30,   -18,   -38,   -11,    14,    -8,   -15,    -1,   -11,     9,    -8,   -14,    19,     4,     8,     8,     1,    -8,    15,    -9,    11,    -2,   -46,   -87,    68,    44,    79,   -28,   -32,   -41,   -22,     4,   -10,    -7,   -42,   -27,   -63,   -34,     2,     0,     6,    17,     0,    11,    -8,     7,     4,   -30,    17,   -26,   -51,   -79,   -97,   -61,   -78,  -198,  -283,  -219,  -177,   -24,    25,    -5,   -74,   -63,   -51,   -89,   -10,   -12,     0,   -18,    19,    54,     4,    29,   -72,   -89,   -55,   -42,    86,   -54,    49,    90,   -72,   -45,     3,   -24,   -75,    64,    19,   -73,   -33,    54,   -37,   -39,   -72,   -35,   -27,    -1,    13,    -5,    78,     0,   103,   122,    68,    55,   -50,   -78,    -1,    -2,   -12,   -29,    15,    -1,   -43,   -34,   -22,   -16,  -108,  -103,   -49,   -89,   -35,   -86,   -44,   -17,    -5,    -2,    19,    32,    85,    98,    31,     4,   -37,    -1,    -7,    66,     0,    59,    31,    18,    -7,    45,     5,  -188,   -11,   -63,  -132,   -71,   -29,   -36,    -8,   -19,   -15,    18,    34,   -48,   119,   -46,   109,    34,    13,    58,    11,    40,     8,    37,    37,   -92,   -49,    -2,    15,   -47,   -32,     0,  -126,   -84,   -54,   -48,   -61,   -19,    -8,   -15,    29,   -51,   110,    23,    16,    35,     0,   133,    72,    39,   -32,   -11,   -47,    -1,    -7,    31,    52,   -39,   -83,     6,   -72,  -189,  -117,   -36,   -81,    17,    14,   -54,    71,    32,    83,     8,   125,   144,    66,    65,    -4,  -117,   -86,   -14,    16,    47,    -4,    10,     9,    42,    17,   -30,  -139,  -141,  -154,   -57,   -42,     0,    15,   -69,    80,   121,   103,    60,    71,    39,  -124,  -181,  -246,  -124,   -99,    24,    36,    79,   -20,   117,    -8,    13,    19,   -41,  -105,    -4,   -83,   -56,   -50,     5,    14,   -42,     7,   117,    44,   -62,  -119,  -195,  -309,  -163,   -35,   -40,    51,   106,     9,   -10,   -62,   -51,    21,    -9,    33,    -6,  -139,  -100,   -57,   -48,   -15,    -4,   -11,   -10,    96,   110,   -70,  -155,  -253,  -154,  -155,    14,    89,    56,    82,    64,    16,   -55,   -97,   -76,   -77,  -157,   -98,  -202,  -100,  -156,   -68,    -3,     3,   -28,   -16,     8,   -27,   -35,   -23,  -100,  -155,  -124,   -62,     8,    80,    25,    43,    26,    23,   -75,   -30,   -54,   -88,   -86,  -119,  -131,   -52,   -36,   -33,   -67,   -51,   -30,   -19,    37,     7,    49,     2,   -75,   -89,   -54,    94,    -4,    25,   -11,    15,    -7,    60,   -31,   -31,   -40,  -109,    26,   -75,   -68,   -78,    33,    -9,  -152,   -74,   -39,   -32,    34,    31,    82,   -48,   -68,   -36,   -23,   -14,    47,    78,   147,     3,    17,    23,    41,    -5,   -82,   -89,     1,     6,    72,   -86,    98,   -11,   -76,   -31,   -49,    20,    13,    38,    75,   -88,  -119,   -70,   -49,    33,   101,     3,     4,    78,    70,    58,   -22,     5,   -14,    -3,   -54,    18,   115,    47,    57,   -18,  -110,  -113,   -48,    11,    24,    40,    82,   -94,  -173,  -170,  -146,   -63,   -37,  -104,   -17,    19,    51,     7,    10,    50,    10,   -15,    17,   -39,    89,    95,     9,   -52,  -171,   -79,   -31,   -29,    -5,    70,   138,   -31,   -98,  -140,  -181,  -288,  -383,  -317,  -334,  -318,  -240,  -161,  -211,   -55,   130,    13,    40,    42,    32,   146,    80,   -59,  -137,   -69,   -56,    -1,   -24,  -116,    75,    63,    72,   -60,   -70,  -121,  -169,  -258,  -280,  -255,  -219,  -174,  -196,  -104,   -45,    18,    89,    82,    62,    94,   106,   -20,   -90,  -115,   -61,     9,    20,   -81,   -45,   -19,    74,    27,   -21,    -9,   -88,   -90,   -76,   -62,   -16,   -24,  -105,  -120,   -20,    -3,    62,    54,   -20,    13,   201,   -12,   -89,     6,     6,   -11,    10,    53,    60,    45,    -8,    59,    36,    -9,   -24,    11,    -5,    40,    50,   -36,   -19,   -50,    -8,    36,    21,    92,   -51,   -55,   -18,   -69,   -80,   -24,    10,    16,   -14,    83,    77,   108,    63,    31,    51,    91,    35,   -10,   -42,    -5,    50,   -65,     8,   -11,   -61,    23,    13,    41,    32,    -4,    36,  -134,   -97,     2,   -15,    -5,     8,    85,   112,   101,   -10,     4,    41,    34,    22,   -19,    45,   -40,    36,   -37,   -28,   -41,   -40,  -104,     0,   -77,   -33,   -80,    -5,   -89,   -15,    16,    17,    19,    19,    27,   -14,   122,    78,    32,   114,    80,     0,    84,    65,    36,   -14,    22,   -40,   -49,    16,   -23,   -76,  -129,     7,    52,    12,   -83,     5,    -3,     1,    17,     4,   -19,   -70,    25,    93,    23,    47,    75,    43,   -17,   -46,   -67,   -87,  -110,   -70,   -24,  -123,  -125,  -124,   -89,   -74,   -42,  -221,   -95,   -19,   -15,     4,    15,     0,    17,   -50,     6,     5,   -66,   -29,   -90,  -105,  -119,  -123,  -106,    40,   -37,   -80,    88,    -4,    22,   -17,   -12,     8,   -61,    -9,    -6,   -16,    12,     2,    20,   -18,    -5,   -10,   -22,    13,   -13,    15,    -5,   -98,   -72,   -53,     6,   -65,   -40,   -49,   -25,    -5,   -30,   -73,   -82,   -14,   -36,   -12,    -6,   -14,   -17,     7),
		    14 => (    0,   -19,    14,   -15,    11,    14,    10,   -19,     1,   -11,    -1,     1,   -54,   -36,     0,    -5,     6,   -18,    -7,   -16,    13,    -1,   -12,    20,    18,    12,    12,    13,     7,    -6,    15,    12,     8,     1,    -3,   -36,   -16,   -27,   -61,   -55,   -75,   -50,   -20,  -168,  -139,  -108,   -31,   -23,   -62,   -32,   -18,   -14,   -11,    -5,     0,    13,    15,   -20,    -7,   -60,  -168,     4,   -14,   -54,   -93,   -69,  -136,  -132,  -136,    -4,    32,    33,  -131,   -88,   -44,   -43,  -126,   -65,    12,    -9,   -14,   -85,    -3,   -14,    -4,     1,     3,   -59,  -167,  -131,   -56,   -26,   -29,   -51,  -122,  -131,   -89,     5,    48,     5,   -98,  -123,     1,    62,    88,    71,   -33,   -84,  -132,   -71,     7,     0,    12,    -7,   -25,  -116,   -51,   -62,   -34,    27,    52,    75,    -8,  -128,  -133,     8,    12,   -21,   -35,   -37,    48,   -13,    71,    16,   -10,   -66,  -128,   -79,   -96,   -15,     2,    14,   -47,   -18,   -43,     0,    50,    32,    82,    43,   -13,  -109,  -110,   -72,    -5,   -50,   -85,    20,    24,    56,    -8,   -14,     3,    -5,   -39,    47,  -106,   -27,   -10,     2,   -81,   -33,    53,    57,    14,    24,     3,   -46,    10,   -43,    50,    40,    94,   193,   193,   144,    91,    80,    16,    92,   -47,   -12,   -27,   -57,     6,   -43,    -5,  -143,   -37,    24,    30,    39,    90,    87,     4,    32,    38,   -11,    48,    56,    49,   126,   144,   114,    13,   -23,     3,    -3,     9,     9,   -39,    24,   -19,  -147,   -68,  -168,   -16,    11,     5,    12,   103,    67,    85,   -18,   -76,   -13,   -43,    -7,   -32,    19,     5,   -34,     1,     3,   -17,    13,   -17,    -8,    25,    54,   -11,  -125,    -8,   -75,   -88,     8,    -1,    21,    -5,   -11,   -15,  -127,  -129,   -23,   -71,  -112,  -133,   -61,   -49,   -52,    -5,   -54,     6,    55,    14,    20,   -44,   -23,   -47,   -93,     7,   -61,    13,    -4,   -44,   -30,   -62,   -45,   -70,   -76,   -50,   -48,   -65,  -162,  -181,  -116,   -99,   -65,    14,   -29,   -70,    70,   -28,  -128,  -153,   -97,   -56,   -29,    -5,   -57,   -47,     1,   -70,     2,   -61,   -32,   -75,   -75,   -60,   -76,     3,   -65,  -147,   -13,   -56,    25,    23,    37,   -29,    36,   -62,  -187,  -178,  -118,   -78,  -121,   -11,     9,    12,    33,   -37,    26,    48,    -9,    40,    43,    48,    15,    69,    54,   -86,    40,    32,    -6,    -6,    31,    46,   145,    35,   -40,  -107,   -67,  -141,  -150,   -11,   -26,   -62,    -5,    76,   -16,     1,   -12,    51,    33,     5,    67,    39,   -24,    27,   113,    56,    64,    69,    81,    54,    35,   -28,   -29,  -113,   -50,  -105,    -5,   -13,   -28,  -166,   -33,    76,   -25,   -18,    -9,   -19,    -1,   -58,   -22,   -75,   -28,    18,   107,    29,    72,   108,    73,    82,    23,     4,   -46,    11,   -63,    95,    15,    10,     3,    83,    21,    58,  -101,   -46,     3,   -27,   -71,  -157,   -92,   -55,    51,    87,   149,   136,   118,   117,   -13,     4,    25,    34,   -34,   -83,   -90,   100,   -81,     8,    -4,    13,    52,    58,   -73,   -76,   -41,   -55,   -94,  -125,   -15,    24,   115,   170,   138,   161,    39,   104,   -39,     7,   -16,   -33,   -48,   -41,    13,    11,   -34,    18,    -5,    40,   -35,   121,   -95,   -40,   -46,   -10,   -89,   -21,    44,   119,   115,   101,   116,   162,    50,    76,   -63,   -33,   -14,    14,     6,   -65,    11,    69,   -84,  -108,   -17,    -5,   -16,    99,   -67,   -41,   -53,  -176,   -40,    24,    40,    89,    17,   103,    98,   114,    38,    -9,   -80,    17,    10,   -18,   113,   -95,  -118,   -32,   -13,    -3,   -28,   -66,    77,    -6,   -19,     6,     6,   -12,    40,    51,   135,     1,   -66,    56,    59,    -8,   -53,    60,    24,   -30,    19,    -9,    -9,   -73,   -59,   -37,   -13,    14,     9,   -33,   -68,  -112,   -93,   -71,    11,    82,    64,    81,    79,    68,    72,   -19,    30,   115,    12,    84,    41,    66,    27,    14,    -7,   -96,  -143,   -82,     4,   -17,   -27,  -106,   -52,  -130,   -14,  -144,    -8,    40,    25,     5,   -47,  -103,   -97,   103,    73,    40,    31,   -16,    40,    29,   -30,    47,    21,   -33,  -214,  -125,     6,   -20,   -31,   -20,   -88,  -264,  -123,   -25,   -18,    13,  -129,    10,   -43,   -58,   -29,   -24,    56,    -7,   -84,   -36,    33,   -21,    42,     3,    47,   -65,  -111,   -47,   -35,     5,     0,    -4,  -146,  -225,  -197,    59,    -6,   -86,   -91,   -41,   -63,   -69,   -30,    29,   -32,   -39,   -37,    22,    75,    12,   -36,   -73,   -10,   -49,   -15,   -28,   -11,    15,     0,   -25,   -29,  -161,    27,    -7,   -57,  -107,   -86,   -96,   -56,   -46,    12,   -15,   -55,     6,   -50,     3,   107,   -66,   -92,   -25,    24,  -102,    55,   -74,     9,     4,    19,    -6,    -8,   103,    76,   -95,  -111,   -89,    -4,   -98,    28,    -9,    58,    27,    25,   -13,   -75,   -45,   -27,   -93,  -121,   -42,    47,   -27,   -80,   -78,   -14,   -18,    12,    17,   -77,   110,     9,   -64,  -151,   -89,   -81,  -102,   -65,  -178,  -136,  -155,  -160,  -108,  -156,  -120,   -59,  -169,  -255,  -268,     5,    -8,    -9,   -17,    -4,     9,     5,   -10,     6,   -14,   -30,   -39,   -68,   -79,   -75,  -140,  -108,   -80,   -90,  -158,   -18,   -87,  -114,   -69,   -94,  -110,   -89,  -107,    -7,   -13,    -6,     8,    12),
		    15 => (   -6,   -19,    -1,    20,   -13,    -8,     6,   -16,    17,    17,    -5,     0,     7,    -3,    -5,    -8,    19,    19,    -7,    -5,   -18,    -7,    12,    -1,     5,   -17,    -1,   -10,   -12,    -2,    -9,     0,    15,    19,   -18,    12,    18,     2,   -16,   -20,   -43,   -51,   -43,   -31,   -42,   -77,   -42,   -29,   -35,   -18,     9,     6,    -4,   -20,     0,   -16,   -20,   -20,   -13,   -25,   -12,    15,   -25,   -58,   -52,  -109,   -50,   -18,   -47,   -86,  -103,  -137,   -59,   -34,     9,    -1,   -25,   -60,   -14,    10,   -31,   -22,   -20,    -9,     4,    -6,   -39,    36,    16,   -43,    -2,   -85,   -86,   -85,   -87,   -45,   -36,   -92,   -93,  -144,  -168,   -92,   -39,   -18,   -18,    29,    28,   -19,   -41,   -49,    10,   -15,   -15,     4,   -23,    25,   -24,   -20,   -10,    33,   -36,    21,   -85,   -70,  -114,  -118,   -22,    29,   -86,   -37,   -47,   -35,   -77,   -18,   -48,    35,    42,   -49,   -87,   -91,     5,   -16,   -27,    -1,   -13,    22,    52,    43,   -79,   -74,    18,   -18,   -58,  -103,    12,    31,   -28,   -64,   -60,   -48,    18,   -20,   -89,  -126,   -96,   -23,   -44,   -61,    12,   -22,   -10,   -51,   -38,    49,    38,   -13,   -56,   -65,   -46,    17,   -38,    -9,    70,   -53,   -83,  -112,   -89,   -11,   -12,   -44,    -8,   -19,   -55,    -5,    -4,    66,    12,   -27,   -23,   -75,   -16,    19,    19,   -51,   -64,  -106,    17,    10,   -38,   -71,    28,   -68,  -102,  -101,  -197,  -185,  -160,   -61,   -10,   -28,    29,    25,    27,    50,    -5,   -89,   -83,   -88,   -65,    74,     2,   -27,  -128,   -36,    51,   -63,   -24,     7,   -82,  -163,   -87,   -71,  -160,  -149,   -80,   -68,   -65,   -19,     8,   -66,  -150,    -3,    -3,   -19,   -30,   -77,   -45,    62,   -64,  -120,   -43,    -9,    32,     1,     6,  -134,   -33,  -118,    34,    34,    42,   -44,   -58,    -7,   -35,    16,    94,    28,   -33,   -24,   -13,   -33,    -7,   -16,   -71,   -31,    -6,   -94,   -16,   -11,    43,     6,   -29,    63,   -21,    27,    93,    94,   103,   106,    84,    47,    60,   178,   114,   147,    35,   -28,     8,   -16,   -23,   -24,   -39,   -47,    52,   -48,    -7,    13,    38,    84,    10,   -27,   -24,   -22,    81,     6,    59,    69,   123,   145,   161,   174,    45,    77,     6,     2,   -14,    -5,   -10,   -60,  -104,   -39,    -9,   -35,   -11,    85,    83,    15,    28,    -1,    51,     7,   -29,   -18,     4,    28,   144,    74,   121,    87,    19,    76,   163,   -20,   -12,   -11,   -13,   -31,  -129,   -25,   -69,   -59,    32,    23,    69,    18,    14,   -18,   -44,  -138,   -30,   -20,  -199,  -124,   -79,  -107,   -17,   -39,   -17,     8,   145,   -45,     1,   -11,   -42,   -98,    62,    48,   -20,    -8,    85,    31,    41,    99,    40,    55,  -127,  -139,  -113,  -100,   -65,  -141,   -47,   -73,   -34,   -68,   -87,   -98,   -51,     6,    22,    16,   -28,   -55,   140,    -8,    27,   -17,   -27,    56,   -14,    21,    98,    -7,   -96,   -75,  -125,  -125,   -38,   -89,   -61,   -42,   -55,   -93,   -12,  -142,   -29,   -41,   -25,   -34,   -36,    -7,  -118,   -76,  -125,   -46,   -92,   -60,   -29,   -31,     6,    -1,   -31,   -16,   -11,    -6,   -15,   -79,  -100,   -28,  -101,   -25,   -51,  -127,   -66,   -47,   -16,   -21,   -30,   -48,   -71,  -102,  -112,  -168,  -141,   -28,  -123,    -4,   -28,   -92,    11,    -7,   -43,    -9,    -5,   -37,    -7,   -32,  -132,    62,   -84,  -149,   -80,  -134,   -13,     3,   -28,    17,    -8,   -16,    -2,   -29,  -102,   -55,   -50,    39,    32,   -60,   -92,  -108,    61,    32,    10,   -63,   -14,   -58,   -61,    37,   -56,   -34,   -86,   -69,    -6,   -16,    41,   -84,   -17,   -85,    56,    50,   -64,   -37,   -11,    16,   -32,     0,    37,    14,    77,    14,    46,     8,   -32,   -83,    27,    74,   -31,  -100,   -91,   -79,   -11,   -51,    30,   -83,   -64,   -44,    46,    79,   -12,    34,    70,   -45,   -13,    21,   -60,     7,    60,    52,   -25,   -22,   -65,    25,    66,    16,   -26,    -7,  -119,    19,     1,   -17,   -14,    -7,   -61,    30,    82,    90,    15,    -2,    21,   -54,   -85,    34,   -69,    28,    27,    -9,    63,     9,    55,    43,    -4,    -8,   -95,   -20,   -92,   -13,     2,    15,   -17,    50,    -9,   -25,    31,   -26,    43,     6,    44,    40,    89,    29,    46,    46,     7,    34,    -1,    33,    54,    16,   -32,   -14,   -82,    -6,   -33,    -9,     4,    11,    41,   -36,   -70,   -93,   -32,   -19,    72,    30,    34,    16,    54,   105,    68,   -38,   -14,    13,   -62,    33,    45,   -33,   -64,     8,    -6,     4,   -16,    -4,   -19,   -13,   -43,    -9,   -12,   -88,   -88,   -81,    69,    78,    56,    27,    12,   -26,    62,    24,    20,    68,   -32,    25,    12,   -89,   -43,    23,    -9,   -92,   -27,    19,     3,   -17,   -18,    15,   -48,  -121,   -62,  -142,   -89,  -133,   -89,   -61,   -84,  -116,   -80,   -49,   -99,  -134,   -86,   -66,   -34,   -26,   -34,   -18,    -8,   -11,    18,   -13,    -3,    14,   -12,   -24,   -18,   -86,  -108,  -101,     1,   -45,    26,   -29,   -80,  -147,  -135,  -139,  -114,   -61,   -90,   -18,   -26,    13,     3,   -50,    -3,    13,     9,   -16,    16,   -11,    -8,   -18,   -29,    -2,   -17,   -27,     2,     6,     5,   -11,   -22,   -25,  -118,   -55,   -41,   -11,    -9,   -47,   -57,   -78,   -76,   -23,   -14,   -10,     0,   -12),
		    16 => (   11,   -17,    15,    -1,    16,    -9,   -10,     1,    20,    -2,    -1,    -8,    30,     6,   -13,     3,    -4,   -11,    16,    13,    -3,    -4,     3,   -14,    -6,    -6,    13,   -17,    -3,     7,     7,   -12,     9,   -15,     5,    56,    18,    15,    18,    23,    70,    31,   -54,     5,    31,    29,    13,     4,    89,    17,    27,    18,    12,     5,    -1,    19,    -7,    -8,    36,     7,    20,    24,    37,    44,    44,   -26,   -33,    -8,   -71,   -55,    33,    27,   120,   137,    14,   -68,   -93,    48,    81,    56,    26,   -24,     1,    -3,   -16,     0,   -22,    -3,    29,    59,   -14,    -8,    -3,   -38,   -30,   -14,   -87,   -25,    59,    69,   124,    53,   -22,    26,   110,    52,   -45,   -15,     7,     1,    -6,   -18,    14,     5,   -57,   -54,   100,    89,   -18,   -21,   -52,   -31,   -28,   -79,   -91,   -39,   -80,     7,   -20,     4,   -52,   -25,     8,   -79,    11,   -70,   -62,   -35,    49,    46,    15,    -5,   -38,    -8,   111,    98,    11,   -10,   -20,    -8,  -103,  -166,   -55,  -102,   -24,   -28,    48,    46,   -31,   -22,  -128,  -105,   -10,   -73,   -14,    -1,    42,    20,     9,    -2,    10,   -53,    68,    56,   -12,    -3,   -26,   -50,  -142,  -156,   -96,   -18,    22,    86,     8,   -91,    48,    43,   -19,  -127,   -23,   -26,     5,   -10,   -18,    23,    16,    -9,    -1,   -98,    50,    68,    -5,   -50,   -40,   -64,  -116,  -154,   -87,     6,    15,  -117,   -69,  -122,   -72,     9,    12,    48,    54,     7,   -16,    28,     9,   -30,    -5,     5,   -15,   -97,    53,    61,    15,    -4,   -61,   -73,  -110,  -164,   -40,    19,    17,   -82,   -44,   -74,  -115,   -77,   -35,    87,    34,   -29,   -22,    -9,   -68,   -94,     9,     1,    -6,   -47,    94,    74,    11,    26,   -35,   -79,   -87,   -21,    29,    42,   -20,    16,   -80,   -55,   -93,   -80,   -78,   -74,   -70,     6,   -19,     6,     2,   -27,    18,   -16,   -31,   -60,    89,    98,   -24,   -34,   -54,   -25,   -16,   -63,    44,    -1,    -6,  -129,   -80,   -92,  -165,  -120,   -98,  -111,   -59,     9,    18,     6,   -30,   -15,   -11,    12,     3,   -71,   114,   107,   -19,   -28,   -54,   -90,   -69,    20,    -7,   -42,   -65,   -92,   -59,  -111,  -149,  -122,   -81,  -124,   -94,    21,    29,    10,   -22,   -45,     7,    -4,   -17,   -53,    62,    91,   -30,   -67,   -64,   -32,   -10,    87,    28,   -47,   -36,     0,   -90,  -137,   -95,   -54,   -43,  -111,   -93,    60,    50,     0,   -57,   -41,     8,     4,    19,   -47,    68,    67,    -5,   -42,   -34,   -47,    -8,    41,   -11,   -10,    22,    32,    87,    26,   -49,   -47,   -27,   -84,   -74,    31,   -59,   -75,   -56,     1,    14,    14,   -18,   -13,     0,    53,    40,    10,   -15,  -108,     2,    -7,    -5,   -32,   -59,   -16,    70,   -55,   -90,     0,    50,   -65,   -70,   -14,   -34,   -35,   -37,   -22,    19,    -2,   -20,   -59,   -20,    15,    24,     0,   -42,   -76,    -5,     6,    -4,  -138,   -22,   -21,    25,    89,    -2,    92,    73,   -54,   -17,   -29,   -53,   -54,   -27,   -75,   -10,    19,   -13,   -63,   -25,    26,    -6,    42,    36,   -81,    -8,   102,    87,   -77,   -22,   -94,   -16,    24,   -56,    49,    -5,   -83,   -38,   -66,   -33,   -19,   -39,   -32,     7,    19,     9,   -68,   -44,   -21,    14,    25,    30,   -82,    53,   128,    32,  -142,  -128,   -48,    14,   -56,   -11,    40,    -6,   -69,   -58,   -30,   -54,  -102,   -18,   -56,    17,     2,    -2,    17,   -52,     1,     1,    -1,   -92,   -70,     3,    14,    54,     5,  -106,   -77,     1,    36,    28,    36,  -107,   -64,   -92,   -76,   -94,  -106,   -15,   -53,     8,    -8,     4,     4,   -25,   -49,   -58,   -61,   -67,   -94,   -11,   106,    60,    64,    -3,   -36,   -66,    49,    21,    23,   -62,   -43,   -81,   -72,   -75,   -56,   -58,   -24,    12,   -12,   -17,   -16,    -2,   -31,   -48,   -76,   -84,  -128,  -110,   -10,    31,    70,   -15,     5,   -24,    76,   -12,    41,    25,   -43,   -35,   -39,   -28,   -29,    -9,     2,    -8,     4,    11,    -8,    15,   -17,   -25,   -54,   -72,  -114,  -107,  -107,     1,    52,     7,   -17,   -40,   -18,    -2,    -8,   -90,   -51,   -29,   -23,   -44,   -53,    -2,    12,    14,     2,     1,   -26,     5,   -18,    19,     0,   -56,  -128,    15,   -43,    -1,    16,    61,    65,   -41,   -93,  -103,    32,   -20,   -28,     9,   -27,   -78,   -22,    14,     8,    11,   -16,   -11,   -27,    10,   -11,     1,   -20,   -21,   -82,   -99,   -58,    15,   -27,     8,   -27,   -35,   -41,    -9,    11,   -39,   -30,    10,    -8,    -7,   -24,    15,     4,    18,    10,    -2,   -21,   -27,   -31,   -24,    -1,   -47,   -26,   -53,    15,    26,    29,     1,    87,   153,    65,  -102,  -151,   -42,    -4,    -3,    -9,   -12,   -26,     1,     5,     7,   -19,     1,   -17,    13,   -21,   -16,   -17,     4,   -29,   -18,     7,    44,    29,   -18,    -8,   -26,   -10,   -17,   -26,   -52,    -8,   -22,   -32,     5,    17,    11,     2,    -3,     9,     9,     6,    -9,    -6,    15,     8,     9,    -4,   -18,   -23,   -12,     7,    13,   -20,     3,     0,     8,   -17,    -6,   -32,     4,    -4,    17,    16,   -19,    11,    -9,   -11,    16,    16,     3,    -2,   -14,    -9,    10,   -13,    -6,    11,     1,     5,     6,   -23,   -13,    -1,    13,    -7,     4,     6,     7,   -13,    14,    -1,     0,     0),
		    17 => (   -5,     5,   -14,    11,    -1,   -12,   -16,   -18,    13,    12,   -14,    17,     5,    19,    17,   -14,    -2,   -13,    17,    -8,   -13,     8,   -11,    19,    -7,     3,     6,    12,   -10,     1,    19,    -3,    20,    16,     5,    -6,   -10,     8,   -16,   -80,   -72,   -50,   -12,   -62,   -66,   -49,     5,     8,    13,    10,     2,   -13,    18,     5,     8,    -4,    -5,    12,     6,   -44,   -33,     4,   -18,    -4,   -29,   -21,   -20,   -61,   -36,   -30,    -1,   -46,   -50,    -7,    -8,    12,   -11,     6,   -19,     1,    15,     6,    20,    -5,    11,     0,    11,   -69,   -13,   -25,   -28,   -52,   -72,   -55,   -44,   -34,   -37,   -54,   -30,   -54,   -15,   -15,   -29,   -20,   -21,   -32,   -93,   -39,    -6,   -28,    19,   -14,     6,    -6,   -16,    -6,   -92,   -44,   -14,  -125,  -120,   -61,  -125,  -204,  -175,  -160,  -123,   -64,   -37,    -8,     7,   -14,   -78,   -96,   -53,  -100,   -25,   -43,   -23,     4,    13,    20,    -7,   -20,   -97,   -47,   -31,    28,    25,   -16,   -81,   -49,    12,     5,  -109,  -133,  -148,  -273,  -311,  -290,  -277,  -164,   -17,  -100,   -65,   -47,   -20,   -11,   -15,    14,    94,   101,    -8,   -16,    -2,   -51,   -50,   -92,  -129,    44,    74,    38,   -45,  -161,  -121,    -2,   -17,   -13,   -38,    99,    59,    22,   -72,   -81,  -132,   -40,   -14,   187,   170,   113,    15,   -17,    -2,    83,   -20,     0,    16,   -50,    41,   -14,   -58,   -84,   -82,   -26,   -10,   -28,   -63,    10,   -22,    48,    41,    -8,   -99,   -46,  -118,   198,    61,    18,   -41,   -66,   -51,   -19,   -86,   -12,    81,     7,    33,   -69,   -57,   -38,   -58,    38,    45,     6,   -25,   -70,   -30,    77,   125,    35,   -76,   -64,     9,   113,   -86,    -9,    31,     6,    48,   -19,   -45,    15,    16,    39,    21,     5,    89,    -7,   -57,    30,    66,    55,    10,    20,    19,    46,   139,   -20,  -128,    -4,    17,    86,    61,    15,    35,    17,    78,    31,    38,    -5,     7,    75,    74,   101,    -7,   -83,   -61,    28,     1,    54,    82,    70,   -55,   -38,   -59,   -44,  -106,    33,    -6,    18,    73,    92,    35,   111,    22,   -45,   -80,    81,    29,   136,   154,    -6,  -125,   -82,   -47,   -19,   110,    58,    78,   -28,   -70,     0,   -34,   -89,   -45,    14,    20,    27,    43,    60,     9,    58,    22,    84,    53,    41,    87,    46,    93,  -246,  -265,   -43,    40,    37,    59,    -1,    31,   -35,   -80,   -81,   -50,   -65,   -10,    56,     2,    33,    92,   -24,   -19,    93,    63,    87,    70,   -11,    12,     8,   -54,  -336,  -227,  -118,    53,    -8,    62,   -55,     0,    38,   -72,  -132,    -7,  -106,   -28,   -16,   -20,    65,   176,    66,   -47,   105,    31,   -27,   -12,    69,   101,    22,  -156,  -441,  -203,   -74,    43,   -12,    87,    47,   -13,   -19,   -20,   -14,     6,   -65,   -49,   -11,   -18,     1,    46,    66,  -160,    40,    59,    52,   -72,   -44,   114,   -57,  -384,  -270,  -143,   -62,    54,    51,    35,    79,     3,   -30,    10,   -64,   -88,   -87,   -10,   -33,   -25,   -25,    28,    26,   -78,   -60,    14,   110,   -18,   -10,   122,  -164,  -372,   -48,     5,   -23,   -28,    15,    70,    62,   -76,    -8,    51,   -47,   -47,   -78,    -5,   -74,   -20,    10,    52,   -29,    14,   -53,    14,    -9,   -62,  -126,  -188,  -257,  -203,   -18,    25,   -15,   -25,   -44,    64,   -55,    19,   -11,    62,  -189,  -246,   -41,    -2,   -91,    45,   -16,   107,  -162,   -68,   -16,    38,     9,   -95,  -191,  -320,   -84,   -26,    51,    91,   -15,    33,    45,    46,   -52,    60,   -44,   -68,  -239,  -227,    25,    -1,   -29,   -15,    60,    39,  -131,   -20,    26,    31,  -201,  -201,  -235,  -248,   -81,    -8,     3,    22,    -4,   -27,   -48,    37,     2,   -37,   -96,  -151,  -177,  -110,    78,    -2,   -19,     1,    70,    -7,   -77,   -46,   -44,   -80,  -190,  -193,  -252,   -55,    93,    66,   -49,     1,   -66,   -43,    13,   -52,   -16,   -63,  -151,  -132,  -187,   -69,     2,    -8,    -6,   -12,     1,   -28,   -93,  -184,   -49,  -168,  -157,  -142,   -55,   128,    41,   -43,   -67,   -40,  -115,   -63,   -10,    53,    13,    -9,   -33,    -5,   -28,   250,    12,   -19,     8,     2,    19,   -18,   -48,  -118,    12,    11,     0,    19,    44,     8,    27,   -51,    -1,    10,     3,   -23,    12,    24,    48,    12,   -42,    -4,   -29,   -16,    -4,   -52,    -8,     9,     9,   -19,  -118,   -64,    69,    88,    55,    61,    -6,    33,  -129,     5,    41,    -1,     0,   -52,   -39,    43,   -81,   -40,   -17,  -171,  -110,   -20,   -37,   -15,   -13,   -13,     1,    28,    30,    -6,    84,   -33,   -96,    59,    -8,    15,    33,    22,    -2,    56,   -34,   -53,   -41,  -123,   -78,   -38,    27,  -138,  -139,   -32,  -116,    17,     6,    13,     0,   -15,    -5,  -140,  -178,   -66,   -47,    -2,   -15,    30,    25,    39,     7,    60,    -3,    37,    54,   -83,   -27,   -35,    35,    -7,   -89,    39,   -21,   -16,    10,     7,     5,    16,    -9,  -156,  -144,  -119,  -129,   -54,   -79,   -74,   -95,    16,    76,    83,    10,    52,   -23,     1,    37,   -34,   -40,   -23,     1,   -38,    13,     0,     6,    16,    17,     9,    -9,    47,    45,    17,    41,    78,    28,    42,    21,   -25,   -17,    21,   -41,   -45,    93,    86,   -73,    43,   140,    35,    75,    -9,    15,     1,    -1),
		    18 => (   14,   -15,     4,     1,    14,    -2,     3,   -15,    -3,   -12,   -18,   -12,    -4,    15,    -7,     7,     7,     6,    -6,   -17,     6,    14,   -17,   -16,     3,     6,   -17,     9,    14,   -16,    -4,    -6,   -13,    15,   -13,    -8,    13,   -18,     8,     4,   -19,   -31,   -49,   -87,  -138,   -64,   -25,   -32,   -26,   -44,   -37,    -2,    15,    16,   -10,    -1,    17,    -4,   -26,    -1,    -2,    -8,   -52,   -33,   -41,  -117,  -147,   -80,   -20,     5,   -27,   -99,   -64,   -24,    28,   -50,  -155,  -128,  -142,   -43,   -30,   -26,    14,    11,   -11,     7,   -59,   -63,    -1,   -52,   -70,  -163,    30,    17,   -19,   -69,   -76,  -116,  -171,    -8,    24,    15,    59,    36,   145,   120,    54,    48,   -52,   -19,   -43,     3,    -3,    18,    -7,   -99,   -90,  -151,    -3,     0,   -63,  -102,    14,   -49,  -134,  -112,    55,     5,    21,   -20,   -20,    46,   106,   116,    67,    44,     1,   143,    62,   -23,   -18,     7,   -75,  -104,  -155,   -51,    -9,    10,    42,   -14,    -6,    -2,   -56,   -53,   -47,    15,    -1,   -65,   -82,   -33,   102,    56,    27,   132,   133,    58,   -52,    -6,     6,     5,   -57,   -94,   -26,   -83,    23,    37,    41,   -11,   -30,   -54,    34,    -3,    21,    -4,   -93,   -99,   -32,    53,     4,   -46,   -97,    33,   -12,   162,    12,   -81,    -8,  -109,   -61,   -19,    -3,   -95,    37,   107,    -5,   -56,   -39,   -24,     8,    -1,    12,    38,   -93,   -20,    66,    28,   -51,     7,    46,    47,    36,   -12,   -18,   -91,   -36,   -31,   -60,    33,   105,   -40,    77,    81,   -75,    41,   -22,    13,    18,    85,   -39,  -131,   -56,   -42,   -49,  -108,    10,    95,    57,   -10,    19,    63,    54,    28,    -7,    20,   -16,    66,    33,   -95,   -41,   -27,   -45,   -32,    32,    77,   -27,   -31,   -95,  -134,    -5,   -19,   -75,    37,    39,    32,    14,    81,    18,    22,   -93,  -217,    10,   -22,   -28,   -65,    -7,   -93,   -66,  -109,    21,    58,    77,    17,   -19,   -76,   -83,   -79,    17,    81,   -30,   -40,   -25,   -35,     2,    53,     2,  -150,   -81,  -170,    -5,   -16,   -59,   -81,   -79,   -55,   -28,    12,   -47,    55,    -2,    92,    76,   -16,   -32,   -58,    -3,   -46,   -30,  -135,   -68,  -160,   -75,    73,   140,    14,   128,   -99,     3,    10,   -92,   105,   -53,    96,    11,    28,   -93,   -44,     2,   -67,    42,    74,   -17,   -55,   -62,    -2,    23,    60,   -96,   -24,    86,   169,   161,    48,    37,  -175,     1,    -5,   -88,    84,   -27,   -53,  -164,   -63,   -75,   -84,   -17,   -18,    16,    46,    10,   -16,  -108,    24,   -12,    44,    59,   136,   196,   170,    86,   -48,   -52,    27,   -29,    -2,    -2,  -144,    -1,  -137,   -66,   -66,  -110,  -141,    -2,   -60,     0,    87,    27,    13,   -99,    72,   -91,    40,     2,    92,    16,   140,    84,   -49,  -117,    -1,    -1,    11,   -21,    53,   -16,    31,    11,   -41,     2,  -125,   -33,    16,    51,    24,    -4,   -39,    57,  -172,   -58,    27,   -61,  -125,   -31,   100,   104,     0,  -144,   -95,    -6,   -16,   -41,    70,  -100,    95,   -24,    22,   -78,   -92,   -46,   -11,    83,    16,   -11,    20,   -83,   -38,   -32,  -110,  -141,  -106,   -72,    51,    19,    38,  -108,   -81,    -3,   -13,   -46,    43,  -150,   -24,   -12,    62,   -47,   -74,     9,    64,    73,   -52,    80,    72,   -26,   -25,  -142,  -119,   -61,  -107,   -67,     0,   -14,    13,   -20,   -52,   -34,   -12,   -20,   -58,  -102,   -50,   -29,   -63,   -77,    77,    58,   110,   -54,  -176,   -35,    86,     3,   -21,   -40,    45,   -33,  -175,   -45,     7,  -111,    13,   -10,   -55,     6,   -17,   -41,   -39,  -119,   -47,   -45,  -103,    84,    29,    93,    88,   -82,  -165,   -75,    29,    20,    65,   -78,   -18,   -53,  -105,    -7,   -68,   -75,     2,   -70,   -27,     1,    16,   -21,   -53,  -179,   -19,   -87,    59,    43,    42,    80,   104,    17,   -47,   -19,    12,     2,   -43,     0,    10,   -54,   -52,   -58,   -72,    -1,    21,   -83,     8,   -17,   -59,   -47,    -8,  -152,  -183,    16,    33,    34,    34,     7,   -12,    32,   -78,   -68,    40,   -88,   -45,    27,   -45,  -173,   -97,   -13,   -63,   -28,    44,   -98,     1,   -22,   -18,   -27,   -71,  -107,  -220,  -105,    27,   -26,    10,    -4,    47,   -22,    48,   -59,   -15,  -162,     0,    14,  -150,  -236,  -106,   -62,   -66,    11,    50,  -140,    -3,     4,     6,   -57,  -100,  -125,  -152,   -54,     5,    89,   -58,   -98,    11,    49,    22,    33,   -75,   -26,    94,  -105,  -230,  -209,   -94,  -100,   -33,    49,    42,  -136,    10,    -9,    -4,   -16,   -12,  -137,  -185,  -100,    -8,    46,     5,   -14,    21,    83,    83,    43,   -20,    40,   -77,  -110,  -136,   -68,   -51,   -63,   -20,   -51,  -111,  -106,     2,     0,    -6,   -67,   -41,   -65,   -98,   -36,   -20,   -77,   -76,    84,   -99,  -115,   -50,   -20,    57,   -38,     2,    32,    62,    61,   -27,   -69,   -33,   -91,   -49,   -51,    -6,    -8,    -3,    15,   -13,   -24,   -72,  -107,   -11,     8,   -58,  -146,  -102,   -83,  -113,  -163,  -152,   -60,   -29,    -8,   -32,   -55,   -60,   -54,   -18,    -7,     9,    14,     8,    -6,     3,   -17,    12,   -35,   -13,    -5,   -52,   -61,   -28,   -29,   -30,   -11,   -38,   -32,     5,   -13,   -16,     3,    -9,   -13,   -12,   -19,     7,    -2,   -13,    14,    -2),
		    19 => (   -7,     7,    -5,    -7,    -2,     5,     0,   -13,    12,    18,    -6,   -10,   -11,   -10,    14,    -1,    17,    13,    -4,    -4,     8,     7,     1,    -9,   -15,     4,   -19,    18,     6,    17,   -13,    -5,    13,    -2,    19,   -13,   -20,   -16,     0,    22,   -24,   -27,    -1,   -47,   -43,   -65,   -25,   -19,     6,   -25,    -3,     3,    17,    14,   -15,    -3,   -16,    16,    20,    -5,     1,    -5,   -10,    -4,    -4,   -23,   -13,   -18,     9,    -7,   -46,   -23,    -3,   -15,   -43,    -9,   -35,    12,   -11,   -20,   -19,   -19,   -10,    14,     3,    10,   -14,    -4,   -21,   -87,    -5,   -12,   -62,    -4,   -12,    -3,    -9,    -2,   -55,  -129,   -65,    27,   133,    48,   -77,   -36,   -45,    -3,   -11,   -27,   -17,    15,   -16,    -5,   -20,   -25,    -2,   -50,   -51,     2,   -24,     7,    17,   -14,   -67,   -89,  -116,  -185,  -204,  -207,  -126,  -152,  -183,   -97,   -91,  -113,   -72,  -103,   -54,   -11,    10,     7,   -36,   -11,   -19,   -11,   -23,    -7,   -85,   -11,   -34,   -75,  -175,  -200,  -259,  -255,  -203,  -173,   -55,   -51,     9,   -23,   -78,  -147,  -107,   -80,   -96,    11,   -11,   -32,   -61,   -61,    41,    -7,   -51,   -58,   -66,  -136,  -106,  -239,  -268,  -144,    -9,   -31,   -11,    82,    67,   -64,   -21,   -39,   -85,  -132,   -73,   -65,   -81,   -91,     8,   -52,   -72,   -33,   -43,   -30,   -60,   -83,   -32,  -189,  -267,  -156,   -51,    40,    42,   115,   100,   -50,    56,   -10,    76,   -60,   -37,    35,  -110,   -80,   -68,   -51,   -82,   -57,   -64,    12,   -19,     1,   124,   -53,    -9,   -86,  -108,   -56,    35,    45,   -42,   -75,    -5,    19,    31,    63,  -114,     5,    95,    69,  -129,  -130,   -69,   -25,    -4,   -61,    66,    59,    72,    17,   -24,   -58,  -150,   -47,    23,    45,    56,     0,  -105,    -4,  -111,  -189,   -63,     1,   -63,   -58,   155,   -59,   -67,  -138,   -24,   -57,     6,   -86,  -151,    69,    78,    23,   -70,  -128,   -56,    36,    43,    81,    26,    18,    10,   -10,   -90,  -107,    -3,    -3,   -35,    12,     1,   -69,   -28,  -112,   -87,   -51,     3,   -37,   -61,    12,   -17,   -12,   -39,    -9,   -51,   -43,   -13,    70,    10,    46,     1,   -10,    26,   -45,    68,     6,   -33,    13,    22,   -48,   -33,   -45,   -92,   -47,    -1,     0,    34,    10,    27,   -67,   -81,    -6,   -12,   -49,    34,    16,    24,     4,   168,   110,    74,   -16,    16,  -108,  -200,   -36,  -111,   -32,   -78,  -127,  -106,  -114,    14,   -40,   -37,   -31,   -23,   -49,    10,   -78,    12,   -38,    86,   121,    63,    52,    49,    57,   -32,     4,   -27,  -249,  -232,   -81,  -112,   -31,     9,   -58,   -54,     4,   -25,   -19,   -60,   -35,   -27,   -19,   -27,    17,   -61,   -59,     9,    15,     1,    16,    75,    26,   -11,   -15,     1,  -207,  -142,  -103,   -63,   -41,    13,     0,    -4,   -15,   -11,    -8,   -81,   -21,   -35,   -78,    -9,    -5,    18,   -49,    40,    14,    30,    32,    60,    38,    99,    36,    59,  -277,  -185,   -58,   -84,    38,    39,   -28,   111,    15,     5,   -15,   -58,    -4,   -18,  -169,  -121,   -45,     7,     6,   155,    68,    62,   -69,   -49,    -9,     9,    15,  -233,  -321,   -97,    83,    26,     7,   129,   -77,   -26,     6,    14,   -26,   -42,   -22,   -28,  -146,  -142,   -77,   -96,   -47,    68,    30,   -95,    -1,    74,    -8,   -49,   -63,  -146,  -150,    53,   110,   -90,   -56,   100,   -37,   -86,    -4,    57,    -9,   -51,   -34,   -57,   -60,   -43,  -194,  -207,   -80,   -12,   -43,  -119,    25,    43,    39,  -103,   -74,  -122,  -127,    95,    95,    10,   -25,    -4,     7,  -102,   -59,    -1,   -53,   -62,   -30,   -87,  -119,   -97,  -146,  -255,  -203,  -154,  -146,   -18,    12,   -28,   -14,  -105,   -51,  -140,   -29,    49,   127,    17,   -42,   -24,     0,   -39,   -53,    -8,     2,   -46,   -49,   -87,   -14,   -57,  -168,  -124,   -64,   -93,     0,    -2,   -56,    -7,  -117,   -85,   -81,  -105,    75,    23,   -25,   -20,   -29,    75,    44,   -15,   -12,   -19,     0,   -61,   -62,   -77,   -36,    28,   -31,    11,   -13,   -13,   -52,    11,   -22,   -34,     2,   -39,  -120,   -66,    84,    86,   -10,     0,    89,  -134,    82,   -57,   -18,     0,    13,   -46,   -91,    -7,    28,   -61,     9,    37,     8,   -45,    18,   -74,  -105,   -54,   -47,   -52,  -158,   -63,    60,   121,    -3,   -35,    79,   122,    -5,     9,   -11,   -11,   -12,   -33,   -27,   -91,    16,   -29,    86,    15,    25,    13,   -86,   -29,   -61,   -80,  -110,   -63,  -101,   -83,    45,   146,    21,    -5,   -31,    85,   -59,    10,     7,     1,    -1,   -19,   -63,   -42,    35,     7,    62,   -10,    15,   -21,   -74,    -7,   -50,   -62,   -85,   -49,   -37,  -128,   -74,    48,   -12,    -2,    10,   -82,   -51,   -68,   -15,   -18,    -3,    55,   -21,    96,   -28,     4,    73,     7,   -98,   -59,    58,   -35,    34,   -74,   -52,   170,    56,   -73,   -43,    29,    34,   -23,    27,  -103,   -86,   -63,     3,   -19,    -7,     9,   110,   122,    13,   -16,    77,   -20,    49,   -44,    67,   120,    51,   111,    26,   214,   193,     6,  -131,     9,    48,   -35,   -31,     6,   -20,    -2,   -15,   -20,    19,    -4,    -8,    -5,   -12,    12,     8,     5,     8,    68,   135,   115,   116,   148,    87,    51,   -24,   -39,   -25,   -42,   -33,     7,   -20,    10,     3,     6,    15),
		    20 => (    4,   -17,    -8,     0,   -16,   -19,    12,    16,    -4,    13,     4,   -19,   -17,   -26,   -15,   -22,    -8,    12,    11,    18,   -15,    -4,   -17,   -10,    -6,    -1,    19,   -13,   -20,   -20,    -8,     4,    15,    19,    -2,   -35,   -61,   -79,   -85,    22,    20,     5,    -8,    74,    43,    42,   -20,    -7,    -7,    -5,   -18,    -9,   -15,     8,   -16,    -6,     3,    14,    -6,    28,    55,   -19,   -28,    -7,   -42,   -80,   -53,   -10,    10,   -34,   -88,   -69,     7,    -6,    12,   -15,    -5,   -21,   -85,   -72,   -27,   -30,     3,    17,     0,    11,   -14,    33,     6,   -74,   -43,   -15,   -83,  -156,   -52,   -57,   -51,  -124,   -89,   -37,   -36,    11,   -39,   -25,  -105,  -100,   -77,  -125,   -51,   -60,   -88,     5,    10,     1,   -34,   -57,   -52,  -136,   -46,   -32,   -45,   -29,    -1,     4,   -80,   -65,   -53,   -27,    46,    67,    48,    46,   -29,   -74,   -64,   -76,     8,  -152,   -64,    19,     5,    -4,   -43,   -19,    26,   -66,   -29,   -80,   -76,    -3,    18,    14,   -26,   -48,    11,    33,    98,    77,    98,    49,   -28,   -19,  -120,   -92,   -10,  -138,   -66,    -2,    -3,   -11,   -50,    -1,   -11,     0,   -10,   -34,   -82,   -69,   -21,   -23,   -56,    10,   -20,    52,    68,    66,    79,    41,    82,    38,     0,   -14,   -42,   -86,   -23,    48,   -17,   -61,   -91,   -63,   -46,   -27,     2,    11,   -96,   -47,   -26,   -14,   -24,     7,    36,     4,    16,    48,    11,    33,    46,   -27,    35,     7,     0,    35,   -77,    13,    37,  -120,    16,   -54,   -71,   -36,   -79,   -45,   -84,   -60,   -51,    -5,     3,    -9,   -30,   -58,   -34,     7,    40,   -16,    10,    48,    13,     9,   -14,   -53,   -72,   -16,   -24,   -26,    21,   -11,   -71,   -66,  -118,   -28,   -78,   -58,   -76,    -5,   -27,   -39,  -103,   -82,   -45,   -71,   -97,   -93,   -59,   -58,   -45,   -44,   -18,  -105,  -111,     1,   -16,    15,    58,    -5,   -82,  -106,   -47,    -2,   -73,   -76,   -94,  -112,  -127,  -125,   -60,   -84,   -55,   -38,   -88,   -81,  -147,  -162,   -47,   -34,   -60,   -46,   -85,   -15,   -12,    92,   -94,    12,   -68,   -26,    37,   -44,  -127,   -98,   -95,  -103,   -98,   -62,   -66,   -33,   -60,   -41,   -38,   -23,   -58,   -77,   -13,   -36,   -27,   -43,   -32,   -18,    -8,    16,  -121,    32,   -42,    -7,   -10,   -49,   -44,   -12,   -34,    -6,    10,    15,    14,   -15,    -4,   -20,    25,     9,     9,    -9,    16,   -23,   -31,   -59,   -51,   -26,     2,    29,    -5,    21,    -8,   -17,    10,   -25,   -61,    -5,   -49,   -25,   -16,    10,    -4,   -67,   -35,     0,    67,     8,   -62,     6,    16,    24,    -9,   -11,   -83,   -60,     7,    -7,   -28,   -77,    11,    -2,   -14,    18,    19,   -11,  -107,   -70,   -50,   -38,  -117,   -95,   -72,   -10,    -9,   -75,   -29,   -18,    -5,   -61,   -24,    55,   -91,   -11,    11,    11,   -22,  -108,    36,    30,   -69,    21,    23,   -76,  -109,  -125,   -77,  -183,  -186,   -86,   -62,     0,   -17,   -15,    37,     5,   -51,   -76,   -14,    13,  -114,   -40,    14,    -3,   -61,   -21,    85,    -1,   -66,   -73,   -13,  -113,  -143,  -102,  -148,  -172,  -114,    -4,     3,    45,    15,     1,    51,   -33,   -52,   -10,    37,    33,  -152,    23,    -5,   -10,   -66,   -17,    19,     2,    24,    11,   -12,    -7,   -91,   -85,   -46,   -54,   -31,    49,    23,    56,   -11,    33,   -19,   -42,   -28,    45,    31,    13,  -139,    27,   -27,   -12,   -48,   -15,    36,   -26,    18,    22,    23,    21,   -23,   -69,   -90,   -64,    -4,    75,    56,    42,    -8,   -38,   -41,   -34,    10,    35,     9,    -6,   -83,   -58,     7,    11,     2,    -2,    14,    12,   -19,    60,    35,    34,   -23,   -24,    -3,   -77,     2,    47,     5,   -78,  -120,   -76,    -8,    72,    36,    13,    70,  -132,   -54,   -46,   -12,    32,    34,    17,     8,    17,   -29,   -23,   -14,   -31,    -5,   -33,   -38,   -68,   -12,    -3,   -48,  -101,   -44,   -11,    -7,   -19,   -10,    40,    35,   -38,   -19,   -19,    16,    12,   -28,    -2,   -14,    -9,   -24,   -15,     6,    -2,   -29,   -97,   -63,  -113,   -52,    10,   -41,   -52,     4,    12,    12,   -69,   -15,    42,    39,     1,    29,    11,    -1,   -19,   -76,     0,    39,     4,    -7,   -12,   -16,    -9,   -84,   -27,   -44,   -25,    -5,   -80,   -13,   -68,    -1,    -1,   -42,    -3,    35,    19,    12,   -19,     2,     8,   -16,    -2,   -69,   -63,   -55,   -35,   -21,   -20,   -88,   -67,   -21,    14,    11,     7,   -45,   -32,   -23,    12,    36,    22,   -25,    36,    43,    15,  -107,   -75,   -45,     5,   -13,     9,    -6,   -47,   -57,    27,   -85,   -31,   -35,   -69,  -151,  -109,   -81,   -75,   -91,   -64,   -45,    25,   -14,    -6,   -31,   -30,   -27,   -43,   -40,   -11,   -11,    11,   -11,     7,     3,   -61,  -104,   -59,   -61,   -52,   -53,   -42,   -66,  -111,  -120,  -144,  -128,   -92,  -101,   -39,   -26,  -122,   -77,   -74,   -83,   -48,     5,    -5,    14,    -8,     4,   -10,   -14,    11,   -77,  -100,  -120,   -57,   -39,   -71,   -76,   -17,   -34,   -72,   -68,   -96,   -83,  -121,  -123,  -136,  -101,   -97,   -77,   -29,    14,     3,     2,     5,    -1,    -4,     5,     1,    -3,     8,   -37,   -65,   -58,   -46,    -9,     7,    -9,   -46,    14,   -23,   -30,   -49,   -31,   -46,   -17,   -35,   -49,   -29,   -12,    -6,    20,   -17),
		    21 => (   16,    -6,   -18,     7,   -11,   -16,     6,   -15,   -17,   -17,   -15,    20,    16,    16,    -1,    11,    -3,   -16,    12,    -5,    13,    -5,    -8,     2,    17,     2,    -9,   -19,    11,    12,     8,    15,   -13,     5,    14,    -4,    18,   -10,   -16,    16,     2,   -50,    87,    93,   -14,   -72,   -26,   -40,     4,   -12,    -8,    17,    13,     9,   -10,   -20,     8,     3,     4,   -17,   -19,     5,   -12,    -6,   -15,   -97,   -90,   -62,  -158,   -44,   -89,   -84,   -16,   -85,   -44,   -24,   -28,  -112,  -141,   -82,   -62,   -30,     8,    -8,    -3,   -20,   139,    90,   -10,   -76,   -17,    86,    74,    90,    25,  -123,   -84,   116,   -19,  -113,   -88,   -32,   -38,   -70,   -24,  -190,  -126,   -80,   -73,   -25,    15,    13,   -15,   -19,   122,   122,    15,   -40,    -5,   117,   116,   106,    70,   -31,   -10,    41,   -12,     1,   -92,   -96,   -29,    10,   -51,  -128,   -66,   -70,   -68,  -142,  -152,  -115,   -12,     4,   112,    17,    33,    60,    60,   115,    38,    94,   151,   157,    78,    82,    10,   -45,   -52,   -35,   -56,    22,   -43,   -94,   -74,    55,    12,  -240,  -109,   -99,     1,     4,   -52,     7,    51,    22,    77,   142,    36,    46,   173,    76,    28,    62,    14,     1,   -25,     1,    -8,     3,   -13,   -86,   -51,    65,     4,  -106,  -132,   -65,    -7,   -98,  -136,  -115,  -171,    67,   105,   167,   -53,   -62,    76,    25,    74,   -35,    74,    -2,    35,    28,   -77,   -61,    55,   -47,    62,    54,   -32,   -87,  -218,  -137,   -25,   -97,  -127,  -183,  -177,   -16,   111,   120,   -65,  -141,    70,   -71,    26,    93,    63,    48,    18,    67,    89,    31,   -31,   -13,    45,   -16,  -107,   -92,  -232,   -90,    17,   -39,  -128,  -174,  -125,   -59,     0,    85,   -32,   -42,   -81,  -107,   -43,   110,    21,    26,   -11,    83,   115,   -25,    18,    37,     9,   -65,   -91,   -95,   -89,  -132,     6,   -62,  -112,  -164,  -134,   -80,   -76,     2,    56,   -65,   -93,  -111,   -22,    69,     1,    -7,   111,   127,    38,   -25,    -8,   -59,   -77,  -113,  -127,   -80,  -144,    13,    -2,    -8,   -43,  -101,     6,   -28,   -45,   108,    41,     9,   -56,   -80,   -20,    25,     2,    17,   144,   212,    59,    -4,    87,  -102,  -135,  -107,  -134,  -116,  -145,   120,     7,    17,  -173,   -72,   -11,    17,    90,    97,    20,   -52,   -47,    -3,    38,    -4,    43,    93,    91,   126,    79,   -24,    14,  -119,  -125,   -34,  -132,   -43,    12,   110,     5,   -19,   -87,     3,   -52,    49,    89,    42,   -53,   -89,   -37,   -53,   -19,   -39,     5,   -33,     9,   150,   -76,    12,    -3,   -92,   -96,  -190,  -150,    37,    90,     9,     3,   -16,    13,    32,   -68,    17,   -61,   -80,     1,   -58,   -84,    24,   -19,   -18,    75,   -10,   -40,   -12,  -168,   -56,    27,   -33,   -36,   -76,  -136,    51,   161,    -1,     6,   -16,    13,   -46,  -126,   -88,   -43,    -1,   -37,   -12,    26,   -61,    -3,    13,    45,     9,   -46,   -98,  -163,  -116,   -33,    25,  -125,  -129,  -180,   -69,    -7,   -38,    -3,    -6,    23,  -118,  -109,    22,     9,   -80,   -81,    50,     3,   -43,    -3,    62,    55,   -97,  -160,  -158,   -48,   -64,     4,    -6,   -28,    -8,    65,     7,   -53,   -38,     2,   -14,   -27,  -180,   -92,    44,   -19,   -61,   -58,   -98,   -78,    60,    68,    47,    70,  -153,  -127,  -169,  -113,   -10,    24,    60,   105,   112,    90,     0,   -81,  -104,   -19,   -12,   -46,  -175,  -119,  -113,  -193,  -123,  -102,   -67,   -42,     0,   -19,    21,     8,   -47,   -95,   -91,    97,   106,   116,   101,    20,   -11,    43,    70,   -57,    38,    15,    -2,    26,  -208,  -154,   -53,   -30,   -22,   -11,    17,    58,    60,   -49,   -67,    47,   -29,   -36,     5,    12,    70,   194,    99,    13,    82,   113,    92,   -37,    13,   -15,    -5,   -94,  -170,   -31,   -11,    53,   -23,    39,    88,   125,    41,    -9,   -46,   -33,    12,    -4,    52,   126,   114,   181,    66,     9,   -11,    50,    31,    -8,     0,    41,    32,  -139,    -7,   -31,    34,   -12,    13,   -17,    42,    84,   -42,  -100,   -67,   -39,    67,    44,   -25,   150,   139,   169,   140,   -19,   -37,    59,    44,   -56,     5,    14,    14,  -122,   -95,   -42,    37,   -16,   -26,    79,    24,    37,   -35,   -73,    -1,   -72,    85,   -21,    40,   244,   162,   100,   143,    31,     1,    54,    84,   -14,     2,   -14,    15,   -41,   -10,   -93,   -26,    13,    10,  -102,   -24,   -47,    -7,   102,    29,    54,   161,    62,    96,   114,    74,   107,    33,    -9,   -89,  -121,   -72,    71,   -20,    -7,   -15,     3,   -21,  -104,   -92,   -99,   -13,  -128,  -142,    31,   -72,    12,    19,    16,    75,    47,   126,    38,    45,    15,    82,    37,   -92,   -80,    38,    19,     6,     6,    -2,   -11,   -53,   -96,  -177,  -198,  -206,  -122,  -300,  -286,  -234,   -26,    -7,   -55,    11,  -109,  -218,  -203,  -251,  -210,  -161,   -65,   -64,   -68,   -59,   -45,    17,     9,     1,    -7,   -45,  -132,  -248,  -229,  -161,  -308,  -302,  -164,  -114,  -152,  -193,   -17,   -18,    37,  -119,   -93,   -32,   -52,  -111,   -11,   -14,    14,    14,    -7,    -8,    15,    13,    -1,   -15,   -28,   -34,   -31,     4,    -9,   -26,  -135,   -77,   -28,   -42,   -64,   -35,   -17,   -10,    24,   -19,   -23,    11,   -11,    -1,     0,    11,    17,   -19),
		    22 => (   -1,    -7,    -8,    -4,     3,    -3,     1,   -16,    12,    10,     4,     7,   -36,   -50,    35,    34,    -5,   -12,     0,   -19,   -16,    -2,     4,    -4,    12,     1,     0,   -18,   -17,     3,    10,    13,    12,    -8,   -47,   -50,  -114,   -86,   -50,   -71,   -51,  -106,   -35,    -1,     2,   -21,   -51,  -194,  -112,   -61,   -66,   -42,    19,     3,    -1,    20,     0,   -11,   -18,   -34,   -64,   -26,   -15,   -64,    43,    86,   103,    94,    78,    54,   -53,   -39,   -23,   -57,  -100,  -119,  -114,   -69,   -47,   -17,    14,    86,    14,    -1,    12,     8,   -40,  -108,  -107,    89,    72,   -58,   -10,   164,    61,   110,   111,    36,    20,   -37,     0,   -14,  -108,   -81,   -41,    71,    -2,  -106,    11,    27,   -14,     6,    -9,    -7,    -3,   -42,    87,   -31,    37,    81,    48,   130,    82,    72,    76,    63,    -6,    22,    40,    62,    29,   -17,    -9,   -76,   -37,   -61,   -44,   -57,   -43,   -45,    -9,    11,    33,    21,    68,    55,   -17,    38,    50,    21,    -8,    -6,     3,    18,    27,    34,   114,    39,    84,   -44,   -31,   -18,    27,   -55,   -57,   -52,   -41,   -41,    -2,     2,    21,     8,    -2,    35,   -32,    13,    79,    26,    17,   -15,    43,     4,    86,   153,    93,     8,    21,    16,   -96,   -64,   -49,  -109,  -187,    -8,   -27,   -32,   -12,     0,    22,   -58,     9,   -22,    68,    65,    54,    64,    -1,    21,     3,    38,    13,   -76,     2,   -14,   -25,   -32,   -74,   -98,   -59,  -184,   -70,    14,   -51,   -10,   -62,    51,   -76,   -85,   -14,   -50,   -22,     5,   -32,    -2,    87,    24,   -71,   -35,   -23,   -26,   -27,    12,    51,    48,    13,    -3,  -120,  -115,   -68,   -68,   -22,   -50,    10,     4,   -15,  -101,   -98,  -129,  -111,   -89,  -137,  -137,   -12,   -15,   -10,   -64,   -88,   -90,    -3,   -36,   -15,   -52,     4,   -37,   -41,  -130,  -147,  -107,    18,   -22,     4,    -3,   -10,  -134,   -83,   -29,    20,   -59,  -121,  -147,   -94,  -132,   -86,  -179,  -129,  -125,   -48,    36,    42,    52,    25,   -64,  -183,   -64,   -20,   -31,   -15,   -49,   -14,   -60,   -55,  -109,   -80,  -133,  -136,  -246,  -213,  -220,  -214,  -210,  -182,  -128,  -130,  -174,   -90,   -11,   -65,    55,   -16,   -52,   -39,    48,    50,    -3,  -129,   -38,    -2,   -87,   -96,   -86,  -175,  -159,  -158,  -244,  -191,  -124,  -106,  -162,   -47,    -2,   -34,   -63,   -33,   -43,   -28,    52,   -29,   -18,   -37,   -63,  -160,    32,   -93,   -24,   -11,   -82,   -30,   -65,  -121,  -138,   -75,    -8,   -38,   -77,   -72,    57,   149,   109,    68,   -48,   -27,     6,    74,   -23,   -17,   -92,   -49,     2,    70,    68,    67,    26,   -17,   -90,   -81,    92,   -19,   -38,    32,    46,    56,    98,   135,   152,   168,    30,    87,    37,    45,     7,    47,   -21,     2,   -59,     2,    13,    90,    14,    84,    95,     5,   -39,    -3,    79,    71,   130,    77,     9,    46,   115,   107,    81,   -19,   -11,    40,    59,     5,   -23,    23,   -22,   -68,    29,   -19,   -34,   -21,    89,    84,   143,   -15,    13,    71,    12,   110,    39,    72,    46,    11,    30,   -18,    51,    -1,   -25,    27,    25,    44,    82,    58,    54,    85,   107,    51,    19,   -34,   153,   127,    33,    16,    -4,    59,   -36,    36,    51,    91,    -1,    90,    -1,    67,   -36,     1,   -95,    25,    60,   -30,    69,    54,    22,    -5,   -64,    31,   -35,  -155,    96,   -21,    75,   -10,    -2,   -42,  -124,   -56,    96,    65,    83,   132,    56,    10,   -77,   -98,    -1,    22,    29,    56,   -23,   -56,    19,    59,   -63,    82,    11,    45,     3,   -30,   172,    -8,   -54,   -15,  -163,   -37,  -133,    18,    26,    41,     1,   -12,  -116,   -99,   -95,    13,   118,    31,    36,    26,   -62,     1,   -20,    33,   -55,    -6,   -45,   104,   149,    -6,   -78,    69,    -8,    28,    14,  -116,     6,   117,   -14,   -78,   -25,   -51,   -21,   -52,   -57,   -53,   -62,    54,   -36,     7,   -57,   -32,   -76,    90,   -87,    88,    -2,    19,    22,    50,    78,    50,   -18,    -6,    -5,    27,    -7,    65,     1,   -51,   -35,   -41,  -146,  -154,   -79,   -64,    11,   -63,    50,    -1,    23,   -96,   -84,  -197,   -10,    15,    19,    47,   140,    68,    15,    19,   -78,   -55,     5,   -36,   -10,  -116,   -66,  -176,  -266,   -51,  -110,    16,     5,   -93,   -76,    43,    18,   -23,  -130,  -210,    -4,    16,    -4,    21,    35,   -32,   -27,  -104,   -83,   -51,   -32,     3,   -47,   -65,  -188,  -116,  -161,  -124,  -130,   -75,  -216,  -134,   -96,    17,   -87,   -73,  -112,  -200,     4,    -9,    -8,  -107,   -47,  -125,   -80,  -236,  -113,  -133,  -172,  -188,  -128,  -215,  -251,  -227,  -218,  -155,   -81,  -253,  -255,  -163,   -68,   -30,  -144,    20,    30,     0,   -18,    14,    16,    -4,   -13,    -4,   -42,   -51,   -95,  -157,  -193,  -112,   -79,  -120,  -138,  -127,  -137,  -184,  -203,  -140,  -176,  -138,   -66,   -49,    -3,    44,    80,    87,   -11,    11,     0,     5,    -9,   -17,   -36,   -32,   -19,   -27,   -40,    -3,   -14,     5,   -27,   -21,   -50,   -71,   -85,   -61,   -26,   -35,    15,   -61,   -10,   -35,    19,   -14,   -17,   -19,    -9,    15,    -5,   -15,    14,   -11,   -18,     0,     9,   -15,   -20,    -7,    -1,   -28,     4,     0,   -10,   -13,     8,   -21,   -39,   -21,    -4,    20,     1,    17,     8),
		    23 => (    4,    -5,    -8,    -6,    15,   -15,    -4,     3,    -8,     7,     4,     8,    -7,   -27,     7,    -6,     3,     3,   -14,   -15,     2,    -8,    -9,    19,   -18,    19,     4,     8,     8,   -13,    -2,    10,    -7,     1,    -5,     9,    -8,   -11,   -50,   -47,   -57,   -30,   -51,   -52,   -51,   -76,   -68,   -28,   -24,   -23,   -20,   -18,    17,    17,     1,    -3,     9,   -10,    12,    18,   -16,   -21,    -1,   -20,  -101,   -80,    11,     1,   -62,   -50,   -67,  -101,  -160,  -110,   -78,   -90,   -55,   -27,   -38,   -84,    -5,    11,   -10,    -7,    13,     5,   -28,    31,   -30,    69,   109,   161,    75,    41,   -61,   -15,    -6,    15,   -55,    22,    57,   -31,  -194,  -116,   -41,  -128,   -79,  -136,   -40,   -38,    19,     2,   -13,    33,     8,    23,    84,    86,    17,    56,   124,    90,     7,   -26,    20,    27,    25,    -8,     1,     8,  -113,  -159,  -219,   -86,  -104,  -190,  -109,   -26,   -24,    -4,    19,     8,    62,    12,    23,    78,    58,     8,    14,     0,    49,    55,    17,    81,    12,    26,    32,   -62,   -75,   -47,  -186,  -168,  -211,  -178,   -86,   -77,   -42,   -17,    19,    22,    28,    56,    21,   105,   100,    24,    70,    98,   105,   -28,    -6,    45,     7,    34,    26,    17,    47,   -26,   -56,  -179,  -186,  -171,   -47,   -50,   -95,   -16,    -3,    10,     2,    80,   128,   130,    44,    24,   -23,   -13,     3,   -24,   -53,    52,    17,    -3,    73,    40,   -28,   -26,  -146,  -184,  -191,  -208,  -104,   -13,   -90,   -45,   -35,   -12,    25,    45,     8,   103,    93,    70,    -9,  -146,   -57,  -248,  -160,   -45,   -39,    36,    59,     8,     9,    87,  -120,  -137,  -194,  -212,  -147,   -47,  -102,    -3,    18,   -28,   -21,   -38,   -36,   -28,   -43,  -188,  -304,  -269,  -167,  -171,   -47,   -27,    63,    75,    43,    25,     0,  -125,  -264,  -188,  -171,   -99,   -76,   -50,   -94,     9,    -6,   -52,    26,     5,  -115,  -197,  -338,  -360,  -219,   -78,    76,     8,    15,    65,    94,   -10,    -8,    40,  -117,  -209,  -265,  -209,   -46,     8,   -79,   -39,   -58,   -29,    16,   -28,   -15,   -29,  -207,  -222,  -201,  -154,    99,    65,    86,   143,    77,    99,    48,     2,  -123,  -124,   -91,  -155,  -133,  -129,   -86,     7,  -104,   -23,   -55,   -14,    15,   -30,   -46,   -73,   -66,   -13,   -33,   100,    90,   140,    61,    20,     2,    20,   -18,    36,   -94,  -126,   -60,   -89,   -75,   -82,   -44,   -56,   -95,   -11,   -45,   -20,    14,   -13,   -33,   -63,     3,    32,    89,   218,   145,    54,    -1,   -61,     1,   -17,   100,    14,    -4,  -112,   -47,   -27,    -4,    -9,   -60,   -17,  -105,   -97,   -70,   -44,     3,     9,     6,   -77,    18,   -42,   -37,    -2,    41,   -17,   -21,   -57,   -61,     6,     3,   -61,   -26,   -42,   -41,    44,     4,    92,    15,    44,    -5,  -204,   -17,   -56,   -25,    48,     3,   -51,   -10,    -9,   -38,  -155,   -63,  -111,   -63,  -110,   -49,    -8,    -3,  -128,     2,    53,   -14,   -23,   -11,   100,    25,    46,    78,  -112,   -16,   -23,    -1,     5,     9,   -65,   -58,   -52,  -116,  -200,   -48,  -119,  -126,  -203,  -290,  -170,   -57,   -86,   -13,    45,     5,    45,    20,    98,   110,    72,    52,  -212,  -173,   -40,   -12,    32,    53,    42,   -64,   -51,   -33,    18,    98,    17,   -38,  -198,  -248,  -183,  -189,   -93,    -5,    34,   -82,   -94,   -19,    28,    47,   -81,   -40,  -216,   -37,   -53,   -22,    37,   -23,    96,    54,    63,   149,   -63,   152,    28,   -34,   -17,   -40,   -86,   -63,   -45,    66,   -53,   -51,    -6,    11,    11,    -9,  -100,   -83,  -108,   -67,   -47,   -18,    -6,  -108,    24,    46,    43,   -38,   -40,    53,   -29,   -37,    55,   100,    83,   -33,   -19,   -91,   -34,   -24,     7,   -43,   -77,     6,   -33,    23,   -65,  -103,   -52,     8,   -10,   -91,    32,   -58,    23,    45,   -23,    32,    46,     1,   -65,   -53,   -57,     8,   -46,     8,    -8,    17,   -70,    11,  -109,   -86,   -32,    38,   -30,   -86,   -20,   -21,    -2,    29,     5,     3,     7,    20,    32,    28,    54,     5,    39,    71,    10,   -70,   -71,    14,   -57,   -16,     9,   -29,   -82,   -25,   -26,   -61,   -21,   -56,    -1,    -4,    -2,    -1,    61,   122,    33,    87,    21,    -2,    33,    28,    18,    -7,     3,    -6,    -2,   -78,   -31,   -29,     5,   -34,   -14,    29,    40,    32,   -81,    -4,   -14,    -7,    10,    39,   163,   164,    34,    22,    76,    24,    19,    20,     4,   -52,    59,   -28,     8,   -21,   -42,    37,     3,    23,     9,   -60,    14,    68,     9,   -18,     5,    -1,    -5,   -41,    30,   -20,   -12,  -117,    57,   -44,   -52,   -42,    39,     0,   -10,   -10,   -46,   -49,   -43,   -17,   -58,   -54,   -97,  -107,   -88,   -56,   -24,     5,   -11,   -12,    -4,    17,   -31,   -24,   -40,    67,    99,    90,   -21,   -39,   -83,  -186,   -77,   -96,   -58,    42,     9,    -6,    82,   -21,  -105,  -148,   -99,     8,   -28,   -14,   -18,    -2,   -14,    16,   -37,   -47,   -57,   -44,    -8,   -53,   -83,   -51,   -66,  -108,  -117,  -144,    -1,    29,   -29,   -21,    13,   -48,   -71,  -104,    -2,     1,    -8,     6,    -4,     5,     7,   -13,    12,    -8,   -14,   -15,    -4,     2,   -22,   -36,  -113,   -70,  -133,    -4,   -30,   -12,    12,    -8,    14,   -28,   -19,   -40,   -19,    18,   -19,    16,     3),
		    24 => (    1,    -5,   -19,    11,    14,   -10,    19,    -8,   -12,     0,   -14,    -7,   -57,   -54,   -28,   -35,    -9,    16,     5,     5,     9,   -20,     5,    14,    11,   -19,    -2,    -3,     7,    -5,     5,    18,     5,   -11,   -55,   -64,   -34,   -86,  -113,   -50,  -168,   -27,    56,   -59,  -111,   -67,   -86,   -31,   -62,   -19,   -30,   -68,   -10,     1,    -7,   -10,   -18,    -1,   -23,  -180,  -199,   -44,   -67,  -137,  -144,   -96,  -130,  -177,  -175,   -60,   -21,  -128,  -108,  -101,   -62,  -136,   -61,   -27,   -18,    -1,     3,   -22,    11,    -3,    18,    -6,   -18,  -153,  -148,     1,   -69,  -144,  -121,  -176,   -18,   -97,  -199,  -119,     3,     3,    72,    49,    53,     2,   -51,    -6,    57,    47,    79,   -50,     6,   -12,   -15,    17,    -6,   -40,    35,  -119,   -17,   -51,   -41,    -9,   -24,    21,   -47,    45,   -77,   -13,    36,   -13,   -68,   -96,    73,    62,   150,   173,    94,    16,   -79,   -23,   -16,     0,   -36,    46,   -65,   -19,   -55,   -86,   -72,   -51,     7,    52,    24,   -43,   -61,   -63,  -133,  -150,   -75,   -31,    47,    -6,    -8,    25,    13,    -4,     9,    13,   -16,   -14,    11,   -30,   -40,    38,   -68,  -107,   -34,    45,    34,   -63,   -80,   -22,   -57,   -45,  -292,  -362,  -156,    -9,    93,    24,    61,    23,   -89,   -35,    10,   -79,    -6,   -17,   -15,   -57,   -25,   -41,   -57,   -48,    25,    12,     6,   -10,    15,    24,   -23,  -186,  -336,  -299,   -86,    56,    45,    85,   160,   114,   -61,  -115,    90,   -68,   -33,   -56,    52,   -39,   -92,   -83,   -55,   -29,   -32,   -96,   -16,   -55,   -31,    53,   -61,  -167,  -295,  -229,   -42,    41,     8,    17,    91,    79,   -48,   -17,    49,   -88,    -4,   -34,    59,   -58,   -58,   -40,   -31,   -57,    11,    16,   -24,   -54,    29,    26,  -115,  -257,  -308,  -183,   -34,   127,    62,    -9,    83,    47,    10,   -10,   -72,   -27,    10,    -4,    47,    75,   -44,   -50,   -79,   -42,    23,     2,   -17,    37,    42,   -13,  -217,  -285,  -194,  -100,   104,   100,    21,   -20,     2,    25,    18,   -26,   -27,   -54,    -9,   -39,   -28,    23,   -45,   -50,   -25,   -49,    -5,   -41,    37,    28,   -14,   -36,   -89,  -180,  -122,   -22,    26,   112,   -40,    -4,     0,    27,   -23,   -56,   -56,   -96,     1,     5,    48,   -60,   -45,   -82,   -43,    15,    15,   -21,    -3,    -7,    38,   -56,  -196,  -107,  -123,   -25,   104,    52,     9,   -52,    -9,    21,   -74,   -89,   -60,  -104,   -17,   -36,   -30,   -61,   -29,    -3,   -16,   -16,    44,   -17,   -10,   -48,     2,   -82,   -93,   -88,   -84,     0,   -45,   -36,   -18,    42,    41,   -15,  -150,   -20,   -63,     1,     0,    -3,   -83,   122,    24,   158,   -24,    32,   -88,    42,    10,     3,   -61,   -93,   -53,   -72,   -51,     2,   -82,    26,    -9,   -32,   -14,   -47,   -56,  -114,    -7,    -8,    -2,    20,   204,   108,    31,    55,   -53,   -14,   -13,   104,    84,    11,   -63,   -29,   -85,   -84,   -81,    44,   -14,    -6,   -13,   -85,    51,   -35,  -196,  -114,   -80,   -27,    13,    19,    66,     4,  -158,   -27,    70,    89,   155,    95,   181,    -9,   -49,    -2,   -64,   -18,    12,   -12,     4,     1,    22,     0,    62,  -118,  -112,  -116,   -51,   -56,   -19,    -9,   -13,  -100,  -102,   -49,    34,   104,   142,    77,   116,    55,   -66,    -9,    19,     2,   -18,    20,   125,    84,    42,    76,    48,    -7,  -133,   -85,    46,   -59,   -20,     9,    -6,  -203,    25,    16,   -16,    25,    23,    11,     9,    14,    72,   -12,    34,    61,    39,    65,    84,    60,    32,    49,    32,   -73,  -146,   -84,     1,    -8,     1,     1,   -19,  -130,   -29,    65,    82,    15,   -14,    14,   -32,   -47,   -76,   -26,     4,    59,     5,     0,    33,    85,    -9,   -89,   -50,   -75,   -14,  -145,   -46,    -9,   -10,   -15,    11,  -148,  -121,   -32,   -77,   -58,   -81,  -135,  -146,  -130,   -29,   -59,    29,   -16,   -59,   -27,   -77,    89,    33,   -46,    18,    18,    26,  -111,   -52,    -1,     2,    -1,   -32,  -121,   -36,   -53,   -60,   -33,  -119,  -226,  -217,   -82,   -62,   -35,     1,   -47,    -9,   -14,   -10,    51,   -16,   -47,    67,    58,   -13,  -128,   -61,   -12,   -17,     3,   -17,  -102,  -117,   -70,   -95,  -138,  -175,  -159,  -172,    79,   -12,   -56,   -71,   -25,    -7,   -56,   -41,    12,   -70,    56,    70,    91,   -54,    13,   -31,   -15,   -12,   -19,   -10,   -30,   -86,   -48,   -96,  -121,   -48,   -46,     1,    63,    29,   -26,   -13,   -69,    28,   -22,   -17,   -26,  -112,    64,    11,    23,   -82,   -48,   -27,   -10,     6,     9,    -5,   -23,   -46,    16,   -13,   -87,   -24,    -2,    -9,   -24,   -18,     3,   -63,   -10,    53,    42,   -98,   -51,  -128,    -6,    82,    54,   -97,   -63,   -23,     6,   -17,    11,   -47,    17,   -22,   -18,   -32,    -2,     9,   -26,     5,   -52,     4,    15,  -134,    -8,   -47,   -89,    21,   -22,  -106,  -122,   -28,    20,   -57,   -11,   -16,   -11,    12,    -6,     4,   -19,    -7,   -22,   -22,    -2,   -14,    43,    50,    33,    55,    24,  -209,  -140,   -55,   -71,  -102,   -23,  -127,  -152,  -133,   -52,   -35,    -5,     6,    13,    16,    13,   -17,   -18,    -7,     5,   -40,   -55,   -67,   -25,   -55,   -48,   -23,     8,    -3,   -15,   -81,  -105,   -24,   -55,   -40,   -87,   -73,     1,     1,   -17,   -17,     2),
		    25 => (  -16,    12,    10,   -17,     5,    -2,     8,    17,     0,   -16,    -7,     5,     4,   -20,   -14,     4,    -3,    19,    -5,     6,    17,   -17,   -13,    -8,    16,   -17,    -8,     6,     6,   -14,    20,    18,   -10,    18,    -6,    -4,     2,    14,   -21,   -40,   -17,   -31,   -14,   -41,   -50,   -68,   -59,   -31,    -1,    -2,     0,    -7,    12,     5,    19,     6,   -16,     8,     3,   -18,     6,    -2,     5,     1,   -32,     3,   -45,   -50,   -37,   -22,   -61,   -10,   -49,    85,    67,   -71,    26,    -9,   -23,   -20,   -26,   -55,   -11,     9,     3,   -13,   -16,    24,    43,   -61,   -31,   -44,   -22,   -22,   -29,   -60,   -80,  -131,   -37,    27,    19,    59,    71,   -50,    35,    72,    27,   -72,   -59,   -27,    65,     9,    11,    -8,   -28,    37,   -24,     8,   -14,   -15,   -22,   -13,   -60,  -183,  -131,  -142,    -5,    62,   -55,    39,    64,    -2,   -43,    -8,   -46,    37,    41,    34,     9,  -111,     1,     5,   -45,    10,   -19,    -9,   -28,   -25,   -28,   -65,  -143,  -168,   -81,   -64,   -53,   -27,    10,   -24,   -40,    -4,     3,   -76,   -31,    76,    33,   116,   -27,   -61,     4,    13,    13,   -20,   -29,   -60,     8,   -49,   -32,   -61,   -82,  -232,   -30,   -36,    80,     7,   -11,   -60,     3,    71,    30,   -20,    91,    81,    97,    93,    -7,    -5,    -4,    -4,     6,   -40,   -33,   -25,    22,    -1,   -50,  -177,   -32,  -170,   -72,   -20,   -13,    23,    38,    14,   -44,     0,   -23,    38,    81,    87,    62,   143,    26,    13,   -19,   -61,   -72,   -30,   -12,   -20,    43,   -51,   -67,   -49,   -17,     7,    90,   -14,   -25,   -13,   -51,   -45,    22,    15,   -47,    44,    86,   133,   119,   130,     4,    65,   -15,    -2,   -79,   -47,   -12,    33,   -51,   -50,    -2,   -16,    49,   -28,    42,   -68,     3,   -16,   -50,    15,   -21,   -37,   -17,   -12,    84,   128,   214,   128,     1,    93,    -1,   -30,   -12,    -4,   -34,    -6,     4,    -3,   -34,  -112,    55,   -41,    34,    43,    99,    -2,   -37,   -58,    45,    50,    61,   -67,    25,    34,   126,    86,    75,    81,   -17,     6,   -27,   -14,    -8,    -4,    27,   -11,    -7,   -26,    56,   -11,    -5,   -19,   -55,   -54,  -141,  -120,  -106,    24,  -140,   -67,   -17,    18,   -23,    31,   108,    30,    13,    11,     8,   -15,   -44,   -11,    26,    18,    57,     3,    23,   -26,    19,    66,   -44,  -139,  -258,  -282,  -257,  -278,  -257,  -259,  -168,   -78,   -85,    -4,    65,  -104,   -12,   -25,     9,     0,   -52,   -12,    60,    47,   -24,    15,    37,   -53,    27,    12,    14,  -109,  -161,  -203,  -271,  -214,  -234,  -230,  -230,  -136,     8,    -1,    94,   -53,    29,     5,   -36,     4,   -27,   -42,   -16,     8,   -14,   -41,    51,   -57,   -12,    -4,   -36,   -43,   -98,  -211,  -255,  -206,  -179,  -151,  -118,  -101,    18,    18,     0,   -55,     8,   -29,   -46,    -1,   -38,  -110,   -94,  -102,    -9,   -22,   -22,   -19,    71,   -42,    19,    28,   -14,    -4,  -113,  -167,  -198,  -146,  -115,   -62,   -35,     0,   -15,   -27,    19,   -28,   -45,    57,   -38,   -87,  -149,  -166,   -68,   -74,   -44,   -24,    -6,    11,    38,    -1,    32,    15,   -91,  -145,  -206,  -140,  -102,   -93,   -28,   -34,   -57,   -22,    14,   -11,  -105,   124,    37,   -88,  -151,  -158,   -70,  -111,  -131,   -24,    50,   -11,    17,   -13,    51,    90,   -94,  -118,  -165,  -104,   -73,  -109,   -90,   -36,   -67,   -65,    -3,   -21,     5,   141,   105,    60,    -1,   -17,  -107,  -126,  -101,   -97,   -55,    21,   -23,   -34,   -49,   -47,   -88,   -56,  -168,   -83,   -56,   -69,   -26,   -28,   -72,   -23,     3,   -11,    25,    14,    97,    74,    98,   122,   -18,   -88,     5,   -71,   -79,    48,   -69,     1,    -6,    78,   -88,   -60,   -77,   -42,   -46,   -63,   -22,  -103,   -52,   -45,   -19,   -13,     7,    17,   -31,    70,    73,   135,    63,    12,   -12,    13,    25,    53,    11,    23,    84,    -7,   -34,  -102,   -68,   -40,   -25,    -4,   -11,     0,   -31,    -7,     5,   -11,    -5,   -26,   -67,   -57,   -75,    65,    75,    34,   -12,    43,    41,    17,    76,    43,    24,   -36,   -16,   -56,   -61,   -19,   -22,   -27,     0,     5,   -23,     3,    -1,    16,   -45,    63,   -11,   -70,     9,    36,     6,    -3,     6,    93,    59,   -11,     7,    19,   -66,     6,   -11,   -58,   -70,     2,     5,   -12,     9,   -37,   -10,   -16,    -8,   -10,    55,    44,    52,   -27,    -3,   117,   105,    97,    42,   107,    63,    22,    41,     0,    -6,    69,     6,   -10,   -33,    -2,    -5,   -12,    18,   -25,   -76,     0,    -7,     2,   -37,   -19,    -2,   -67,    22,    77,    13,   129,    88,    80,    75,    36,     8,   -45,   -60,    37,   -40,    19,    -6,   -13,     4,   -10,   -10,  -109,   -38,    17,   -11,     8,    11,    -3,   -90,   -82,   -13,   -69,   -45,    60,   -16,   -39,   -41,    -7,  -108,   -93,   -62,   -44,    72,    34,    -2,   -34,   -20,   -12,    12,     1,    -2,    -2,   -13,    -9,     0,   -11,   -44,   -42,  -142,  -140,   -59,   -25,    39,    69,    91,    39,  -116,  -141,   -36,    -1,   -40,     3,    11,    14,    20,   -51,    12,    -5,    -1,     1,    11,    15,     8,    -2,   -29,     4,   -30,    -2,   -18,    -9,    -4,    20,    17,   -10,   -25,    -1,     5,    12,    -5,   -20,     6,   -15,   -70,    -2,     2,   -18,   -18,     1),
		    26 => (    6,    -5,    18,    -6,   -14,   -14,     6,    18,    -7,    -6,     6,   -16,    76,    58,    -7,     7,    -6,   -12,     6,     7,     4,    -6,     9,     2,    11,    -6,    15,    -9,   -18,    19,    -7,     4,   -14,    -9,    53,    79,    88,    56,   173,   155,    27,    72,   -74,    14,   -32,     8,    58,    70,   208,    74,    41,    82,    18,    -3,     8,   -19,   -15,    -2,    29,    52,   107,   146,    63,    98,   188,   153,    81,    88,  -146,   -92,    -3,   -10,    -9,    92,    52,    -7,    61,    62,   117,    67,    14,   -83,   -14,     7,    16,     5,  -167,   -32,    -7,   142,   123,    39,    18,    13,   -23,  -106,  -147,   -25,    66,    40,   -23,    62,    61,    45,    -8,   -49,    14,   145,    72,  -114,   -88,    11,    -4,    10,  -152,    -4,    -1,   114,   -12,   -32,    82,   107,   -37,   -84,  -237,   -62,     7,   -69,    33,   -23,   -81,     7,   -37,    62,    72,   135,   -13,  -158,    88,   139,    20,   -11,  -125,   -99,    44,   -55,  -146,    80,    53,    20,   -96,  -209,   -81,   -50,     4,     0,  -120,   -20,  -116,   -68,    -8,     3,    23,    91,    19,   -79,   187,   123,     1,   -17,    51,   -32,    25,   -50,   -96,    52,   -39,  -142,   -87,  -103,    14,  -110,  -104,   -10,   -44,   -32,   -15,    20,   -31,   -68,    79,     3,    43,   -61,    53,    74,     0,     6,     4,   -61,    34,   -21,   -51,   -24,   -67,  -107,  -105,   -17,   -24,   -50,   -36,   -59,   -17,   -33,   -87,   -27,   -37,   -15,    -3,    16,    19,    -7,    34,    59,   -14,    20,   -79,   -67,    45,   -65,   -98,   -92,   -67,  -125,   -13,   -36,   -66,   -47,   -87,   -90,   -60,   -82,  -169,    -3,  -147,    -6,   -36,   -33,    49,  -200,   -38,  -138,    17,     2,   -95,    32,    21,  -152,   -42,  -111,   -99,     5,   -14,    19,   -69,   -53,   -24,  -136,  -211,  -187,  -201,  -112,  -118,  -111,  -295,  -101,    24,    -9,   -47,  -144,   -13,   -12,  -120,   -99,   -60,  -116,  -161,  -165,  -100,    41,   -65,   -25,    16,    -9,   -72,   -89,  -150,  -116,   -73,   -54,   -58,   -55,   -92,    72,    88,   139,   -81,  -177,    12,    -9,     8,   -71,   -46,   -52,   -89,   -10,   -20,    23,    59,    42,    23,    99,    30,   -32,   -17,   -51,  -110,  -139,    31,   -79,   -68,    21,    22,   -37,   -98,   -45,    10,    -2,   -18,   -77,   -60,  -117,    -2,    49,    93,   130,   123,    42,    12,    25,   -12,   -26,    34,   -21,   -88,  -196,  -148,   -37,    68,   139,    95,   -12,  -163,   -31,    16,     3,   -37,   -63,   -66,   -10,   122,    59,    22,    87,   123,    32,    13,   -46,   -29,    -2,    -7,     9,   -74,   -60,  -100,   -57,    38,   141,    91,    46,   -50,    17,     0,    16,   -19,  -127,  -103,    85,    39,    46,    97,   134,    38,    81,    -9,   -75,   -13,   -11,    33,   -28,   -34,   -23,   -29,    55,   107,    86,    29,    43,  -124,   -86,     7,     6,   -50,  -143,  -125,   101,   109,   121,   176,   163,   101,    75,    77,    21,   -38,   -70,   -20,    -1,   -14,    33,    17,   -32,   107,    91,  -106,   -53,  -165,   -85,     7,    -7,    -2,  -121,   -19,    76,    64,   134,   212,   189,   139,   127,   125,     9,    22,   -13,    47,   -26,   -37,    98,    56,    24,    79,   108,   -62,  -108,  -153,   -90,   -14,   -20,    -8,  -114,  -118,    48,    50,    90,    72,    70,   154,    52,   128,   162,    13,    -8,   -22,   -45,   -23,    41,    36,    78,   -10,   -20,   -38,  -117,  -181,  -141,    17,    -5,   -19,   -11,   -68,   -48,   -16,    70,   -41,    46,    43,     3,   113,   160,    49,   -94,     5,    -2,   -56,   -92,    -8,   -24,   -43,   -68,  -190,  -134,   -94,   -95,     9,    -6,  -100,     8,     0,  -137,   -94,   -29,   -83,     3,   -26,    60,    52,    21,    -3,   -28,   -39,    53,   -54,   -43,   -37,    -9,   -18,   -15,   -88,    25,   -72,  -117,    15,   -28,    -8,  -136,    29,  -103,   -90,   -76,   -61,    18,   -24,   -10,   -25,   -78,    63,   -14,   -89,   -57,    -9,   -42,   -21,   -41,    88,     1,    69,   134,   -27,     3,   -16,     2,   -46,   -65,   -62,   -49,   -89,   -28,   -19,    27,    16,   -83,   107,   107,    11,   -67,   -17,     3,    15,    64,   -17,    -6,    82,    94,    88,    38,   -17,   -38,     9,   -12,     0,   -47,   -67,  -177,  -179,  -112,    50,   -63,     7,   -52,    84,   104,    31,    49,    79,    13,    18,    39,   -30,    66,   -31,    -2,   -59,  -145,   -19,   -26,    19,     2,    16,   -19,   -82,  -139,  -166,  -124,   -73,   -39,   -46,     7,   -54,    12,   -17,    34,   -56,     1,    80,   109,     4,   -93,  -151,  -120,  -110,  -109,  -167,     8,    20,     8,    -4,    -4,   -49,   -43,   -22,  -109,  -113,  -164,  -182,  -128,   -46,   -82,    13,    52,    73,    81,    22,  -196,   -82,  -194,  -117,   -91,   -59,   -73,     8,     0,    13,    -5,    -1,   -16,     2,   -32,   -28,  -100,   -51,   -62,   -91,    -4,    94,    -3,   -76,   -32,   -88,   -76,   -28,   -73,  -142,   -45,   -55,   -50,   -39,    -6,    -3,   -11,    15,    -1,     9,   -14,    -2,   -33,   -47,   -21,    -6,   -24,   -61,   -49,   -11,   -19,     2,   -25,   -12,     5,    -8,   -19,   -26,   -33,   -22,   -12,   -22,     9,    -3,    16,   -18,    -3,   -14,    19,   -16,   -17,    17,     5,   -10,    -7,     1,     4,    16,    -4,   -16,    -6,    -1,   -21,     2,   -21,    -4,   -28,    -6,   -10,    -5,   -20,     2,    -1),
		    27 => (   20,     4,    18,     3,    13,    13,    -7,    17,     7,    -9,   -13,    14,   -11,   -15,    -5,    -6,     4,   -18,   -16,     0,   -16,    14,     4,     0,     3,     5,   -13,    -2,   -18,     9,    -2,   -19,   -17,   -17,    -8,    18,    18,    -7,    -4,   -88,   -62,   -78,    -6,   -17,   -29,   -20,    11,   -10,    -6,   -18,   -20,   -18,    -3,   -10,   -12,   -17,   -15,    10,    20,   -25,   -30,     3,     0,   -27,   -20,   -12,   -25,   -51,   -90,   -56,   -19,   -17,    -6,    14,    -8,   -21,     0,    -8,   -28,    -3,    10,   -15,    -2,    12,    18,   -19,    -2,   -40,   -42,   -32,   -31,   -50,   -78,   -73,   -54,  -102,   -73,   -36,   -15,   -27,   -53,   -46,    -6,   -52,     1,   -67,   -52,   -33,   -15,     4,    17,    10,   -15,    15,     2,    -6,  -106,     1,   -27,  -101,   -91,  -127,  -173,  -162,  -146,  -172,  -127,  -138,  -105,   -47,   -40,   -24,    -4,   -73,  -112,   -84,   -69,   -51,   -31,    11,    -6,    15,     9,   -61,    20,    27,   -26,  -100,    78,    64,   -86,   -69,  -116,  -101,   -88,  -118,  -156,  -322,  -388,  -257,  -178,   -66,    -6,  -176,  -134,  -130,   -64,    -3,   -10,     8,    20,   172,   135,   108,   -48,  -101,   109,   -12,   -65,   -10,    53,    68,     6,  -120,   -22,    16,    68,   -14,    45,   156,    -5,  -222,  -165,  -155,  -109,    -6,   -11,   126,     1,   133,   128,   -40,     3,     8,    13,    56,    98,    84,    57,     1,   -18,   -23,    30,    35,    12,    93,    65,    84,   126,   141,    -8,   -64,  -126,   -62,   -94,   153,    35,   100,    52,   -84,   -72,    26,    56,    14,    11,    37,    25,    30,    -8,    30,    43,   -17,    29,    39,    27,    64,    47,    26,    48,   -88,  -170,   -39,    -9,    96,   -48,    17,    56,    43,    -3,    71,    76,    99,    95,    63,    99,     3,   -26,   -12,   -30,    18,    -6,    80,    30,   141,    30,    -4,   -16,   -34,  -158,     1,     3,    57,    -5,   -65,   105,    82,    14,    38,    48,    45,    18,   110,    18,   -36,  -137,   -73,    10,   109,   -19,    59,    76,    41,    30,   -41,   -81,   -98,  -100,    22,     6,   -46,   121,   -20,    99,    32,    36,    77,     6,    16,   132,   167,   -21,  -203,  -304,   -52,    33,    57,   -18,   -12,    74,   -34,   -19,   -35,    24,  -144,   -35,    11,     0,    67,    16,    12,    10,    82,   -65,    49,    12,     0,    80,   -22,  -182,  -458,  -301,   -31,    39,    -9,    30,  -134,    -9,    23,   -16,  -166,    -8,   -53,   -43,    20,   -12,    77,     6,   -16,   -68,   -21,    28,    59,    76,    61,    48,    -4,  -282,  -487,  -180,   -58,    18,     1,   -94,  -131,     7,    18,  -130,  -162,   -57,   -40,   -52,   -28,     0,    15,    71,    13,   -18,   -46,    85,    46,    36,    38,   102,  -148,  -407,  -414,    -7,   -15,    22,   -25,  -111,   -19,     0,   -63,   -63,    10,    64,   -42,   -27,    -8,    -1,   -16,    67,   -18,   -63,    19,    -3,    77,    -4,   -23,     2,  -266,  -452,  -104,   -54,   -91,   -15,   -40,   -27,   -14,    31,   -30,   -14,    26,    68,   -11,     1,   -16,    20,     5,    60,   -59,   -76,     2,   -45,    -3,   -19,  -105,  -124,  -263,  -151,   -51,   -72,   -48,   -74,   -34,   -57,   -34,    16,   -13,   -42,  -125,  -141,   -64,    -6,   -42,    12,     2,    -3,   -50,   -68,   -47,  -176,   -94,   -73,   -71,   -52,   -38,  -139,  -114,   -65,   -42,    12,     5,    68,    28,   -10,    22,    -2,  -129,  -168,   -77,    -1,   -84,    20,   -14,   101,  -113,  -131,   -24,   -74,   -82,   -89,   -15,   -24,  -100,  -122,   -75,   -17,   -80,    12,    40,    44,    30,    -7,  -110,   -54,   -88,  -193,  -151,    -1,   -52,    20,    48,     8,  -128,    20,    64,   -23,  -150,    76,    77,   -45,    -4,   -51,   -31,    28,   -35,   -27,   -68,   -68,   -20,   -11,   -87,    27,   -88,   -95,   -52,   -14,   -17,     3,    97,   -24,   -35,   -52,  -142,  -115,   -33,    -9,    20,    12,   -34,    93,   -44,   -14,   -18,   -96,   -66,   -81,    -5,   -83,  -203,  -153,  -151,  -123,   -12,   -44,    17,    -4,    18,   -11,   -74,  -135,  -113,  -105,  -159,   -36,   -66,    18,    85,    33,    -9,    10,   -34,   -31,   -85,   -31,    12,   -18,    43,    35,   -71,     8,    -9,   -54,    -4,     5,     7,   -23,   -64,   -92,    30,  -105,   -72,   -25,    12,    -7,   -43,   -39,    21,   -23,    19,   -53,   -44,    31,    31,   -76,   -33,   -50,   -72,   -34,     7,  -162,     8,     2,    11,   -29,   -78,    24,    96,    40,    16,   -64,    39,    70,   -50,  -109,    16,   -52,     4,     9,     9,   -50,   -12,   -84,     7,  -102,   -62,   -29,   -12,   -88,    -9,     2,   -11,    51,   107,   223,   133,   -14,   -40,     6,   -59,    81,   -43,   -32,  -123,  -154,    24,   -34,   -23,   -49,   -14,   -72,    17,   -54,   -32,    -7,   -39,    -5,     9,    13,    16,  -101,    77,    17,  -122,   -90,   -14,    30,    -3,  -104,   -46,    83,   -15,    70,    31,    -3,    19,     8,   -32,    21,   136,    68,   -72,   -21,     4,    11,    -1,    -3,     2,   -20,   -62,  -101,  -141,   -59,    84,   112,   -22,  -109,   -89,   -70,    31,    -1,    66,    33,   -44,     0,    94,    65,   -18,    -8,   -25,   -36,   -21,    -7,   -20,    -1,   -16,     7,    -2,    85,    99,    35,     7,    53,    53,    36,     8,    13,   100,    99,   -20,     0,    98,    27,    78,    60,    21,    18,   121,   -19,   -10,   -16,     7),
		    28 => (   -2,   -16,   -11,    -4,     3,    20,   -17,    -5,     1,   -10,    19,   -13,   -18,   -18,    -1,   -12,    16,    11,   -15,    -2,    -8,    18,     0,     2,     0,     1,    -4,    10,     5,   -18,     6,    16,     2,    20,     6,     0,    14,   -19,   -18,   -70,   -71,   -83,   -83,  -154,  -121,  -156,   -23,   -34,   -10,    29,     8,     9,    12,    -1,     6,   -20,    16,     1,    -2,   -15,   -24,   -11,   -39,    -4,   -58,  -136,  -220,  -202,  -101,   -76,   -33,  -181,  -182,  -162,   -70,  -129,   -75,   -87,  -108,   -86,   -31,   -35,    14,     3,    12,   -18,   -70,   -51,   -34,  -134,  -223,  -275,  -325,  -355,  -222,  -199,   -48,   100,   -56,    -9,   -55,  -111,  -225,  -215,   -55,    35,    77,    96,    64,    -3,   -44,    -7,    -6,   -77,   -45,  -134,  -165,  -265,  -124,  -117,   -38,   -52,    -7,   -92,   -87,    48,    43,    -2,   -25,   -59,   -83,    38,    70,   -81,   -62,   -65,    52,   -82,    96,   -13,    11,    -9,  -116,  -102,   -87,  -223,     1,   -14,    25,    -6,   -75,   -12,   -35,    -1,    52,   -57,   -26,   -15,  -120,   -21,   -20,    86,    60,   -31,   147,   122,  -101,    25,    -5,    -3,   -38,  -183,   -67,   -91,    60,     6,    -2,   -13,   -20,    33,    31,   -59,   -55,   -25,    25,   -15,    58,   -51,    40,    67,    75,   107,    37,   -81,   -88,     8,   -17,   -67,   -42,  -160,    10,    38,   -15,    61,    14,   -18,    50,   -10,   -35,   -57,   -97,    10,    11,    -1,    18,     1,   -84,    72,   132,    44,   -39,   -67,  -126,    20,   -63,   -84,  -140,   -10,   -17,   -42,    37,    44,   -14,    69,   -17,   -75,   -46,    26,   -51,  -140,   -92,    26,    62,     6,     2,   -15,    89,    54,    98,   -79,    67,    61,   -13,   -62,  -151,   -15,  -120,   -25,   -24,   -46,    67,   -18,   -44,   -38,   -60,   -28,   -88,  -117,   -48,    42,  -103,    77,   -37,   -47,   -23,    83,   111,    -6,    51,   -61,   -17,   -22,  -205,  -183,    37,   -22,   -35,    54,    -7,    64,   -46,   -15,   -24,   -64,   135,    25,   -37,   -56,   -29,    27,    18,     2,    16,   165,    91,   -95,    34,   -27,     3,   -17,  -125,   131,    42,    35,   -25,   -12,    43,   -10,    16,    -6,    33,    69,   130,   144,    14,   -11,   -28,   -24,    42,    42,   -13,    52,   202,   198,   105,   -83,     5,    -7,   -87,   150,    88,    66,   -47,    11,    -6,   -88,   -90,    87,   139,   143,    78,    91,    46,   115,   -37,   120,    34,    -1,  -124,   -24,    51,   138,    64,   -91,    -5,     4,   -54,   177,    11,    20,   -30,    43,   -59,    10,    26,   132,    85,   133,   116,   107,    69,    60,    73,   100,   -35,  -134,    19,   -62,  -122,   -15,   -46,     7,   -12,   -14,   -24,   129,    39,    22,    38,   -61,   -98,   -17,   162,    97,    73,   133,    65,     8,    66,    53,    60,    43,  -123,  -161,   -91,   -66,  -108,   128,  -127,     3,   -10,    -7,   -47,     1,  -175,  -120,   -43,    39,    19,   103,   113,    84,    72,   128,    86,    43,    79,    57,   -14,   -67,   -88,  -131,    23,    36,  -144,   143,  -286,   -96,   -20,   -18,   -26,   -22,   -39,   -30,    30,    18,    39,    52,   159,    45,   142,   -12,    34,    25,   133,   -85,   -57,    10,  -108,   -55,   -23,   127,  -159,    64,  -236,  -107,   -12,   -14,   -28,  -104,   104,    43,   164,   -27,   -62,    68,   115,   155,   137,   152,   112,     0,   141,     5,   -98,   -44,   -72,   -45,    29,   199,    64,  -118,   -58,  -145,   -18,   -24,   -45,  -127,   119,   -12,   -36,    23,   -27,    18,    70,    99,   198,   237,   107,    87,   -25,   -63,   -49,  -114,   -35,   -65,   -39,    44,   -29,  -139,   -75,   -55,   -17,   -15,  -148,   -61,   -63,    -7,    51,   -31,    53,    27,    27,   -76,    17,   114,    31,   -66,  -145,   -84,    -4,   -35,    20,   -35,    49,   -62,   -27,  -169,  -224,   -52,    -3,    -2,   -58,    -5,   -18,    13,    55,    21,  -112,   -30,   -50,   -86,   -64,   -64,   -29,   -55,   -38,   -86,     2,   -34,    49,   -56,    75,   -87,   -68,  -130,  -133,     5,   -67,   -12,   -93,    20,   -39,    16,   -11,   -59,   -99,     0,  -114,  -157,  -128,   -89,   -74,   -99,  -100,    80,    88,   -46,     7,   -26,   -16,   -86,  -206,  -125,  -225,   -37,   -41,   -33,   -51,   -10,    32,   -93,   -35,     7,    16,   -20,   -47,  -100,   -68,  -116,   -89,   -24,   -77,  -111,   -30,   -45,   -20,    86,   -79,  -112,  -161,    29,  -100,   -10,    -9,    -5,   -68,    33,     9,    -1,  -119,    -8,    27,    57,   -80,   -67,   -75,   -15,   -95,   -12,   -12,     6,     4,    70,   117,   -73,    32,    72,   -74,    31,  -134,    -9,    17,    18,   -60,   -46,  -221,  -169,  -144,  -201,  -118,   -10,    -3,   -33,    -5,   -23,   -85,   -53,  -106,  -141,   -74,    97,   -37,  -129,   -47,    23,   -51,   -75,   -34,   -18,     5,    -9,   -68,   -50,   -48,   -13,    92,    72,   -36,   -14,   133,    19,  -125,   -63,    -9,    48,    75,    -1,    39,   -92,   -50,   -86,  -129,   -90,  -137,   -91,   -56,    -8,    -3,     7,    10,   -56,   -60,  -124,  -159,  -157,  -192,  -280,  -221,  -111,   -97,   -96,  -107,  -276,  -145,   -90,  -116,  -219,  -165,   -99,   -61,   -60,    -4,   -18,    -3,   -18,    -4,    10,    10,    -9,     1,   -19,   -15,   -68,  -120,  -134,   -81,   -18,   -41,  -101,  -119,  -145,   -89,   -96,   -60,   -74,     8,   -17,    -9,     2,    -1,    -3,    13,   -11),
		    29 => (   17,     0,     7,   -19,    -3,     1,   -16,    17,     0,    15,   -20,     2,    18,    13,   -18,    14,    -3,    -8,    -8,   -13,    -9,   -16,    -6,    13,    -4,     0,    -5,   -18,     1,     4,    19,    -1,   -12,    10,     2,     6,    11,   -17,    -3,   -31,   -50,   -33,     4,   -21,   -63,   -84,   -69,   -41,    16,   -32,    -5,    -6,    13,   -12,     8,   -19,     2,    13,   -12,   -26,   -32,     3,    -4,   -39,   -14,   -34,   -35,   -67,    -5,    -5,  -120,   -88,   -72,   -22,   -20,   -16,  -147,   -52,   -96,   -58,   -26,   -12,    -1,    13,    -6,     7,     9,   -26,   -52,  -125,  -117,  -105,  -136,  -133,  -238,  -241,  -161,  -185,  -348,  -138,  -172,  -254,  -189,  -127,  -201,  -217,  -146,   -81,   -54,   -26,   -11,     7,    13,   -11,   -55,   -55,   -65,  -208,  -290,  -107,  -130,  -159,   -76,   -49,   -34,   -25,   -58,    27,   -32,  -118,   -39,  -293,  -254,   -75,  -109,   -58,   -43,  -144,   -94,   -14,     6,   -16,   -10,   -26,   -20,   -78,   -99,   -96,   -52,    15,    21,    81,    18,    58,    40,   -21,    21,    50,    94,    97,    33,  -129,  -133,  -123,   -43,   -98,   -68,    10,   -16,    14,   -16,   -84,   -74,  -138,   -51,  -100,     1,    89,    40,   -48,   -88,    17,    23,    52,    33,    -7,   120,    76,    91,   -29,   -42,    53,    15,   -33,   -69,  -120,    -7,   -18,   -92,   -67,   -94,  -111,  -138,  -117,    -3,    32,    19,   -45,     1,   -73,   -11,   -47,   -30,    -9,    -1,    32,   -43,   -81,   -94,   -24,    19,    55,   -79,   -43,   -63,   -75,   -38,   -31,   -31,  -101,    27,   -21,    40,    98,    61,   -24,   -25,   -14,   -45,   -23,   -15,   -34,    12,   -52,  -134,  -109,  -121,   -71,    36,   -14,   -93,   -32,   -13,   -73,    38,   114,   114,    46,    54,     0,    44,   106,   -13,   -17,   -32,   -52,   -54,   -62,    30,    80,    76,   -37,   -18,   -39,  -107,  -163,   -93,  -132,  -213,   -80,     9,   -99,   -85,    63,   242,   131,   142,    88,    19,    23,   -32,   -41,    32,   -40,   -42,    35,   176,   141,    17,   -49,   -53,   -37,   -74,   -55,   -64,    33,   -63,   -38,    12,  -192,   -16,     5,   131,   137,   126,    19,   -68,   -14,   -20,    21,   -24,    57,    87,    52,   197,   134,    11,   -99,   -52,   -15,    49,    41,    15,   108,   -26,   -55,    14,   -47,    28,   -43,    98,    79,   109,   -29,   -10,   -25,   -34,   -12,    -8,    40,   201,   141,    82,    15,    30,   -31,    38,   -14,    25,    36,   -53,   -67,   -76,   -52,    -8,   -55,   -31,   -52,    73,   113,   -19,     3,   -48,   -54,   -26,    17,     7,   149,   184,   196,    89,    24,    40,   -45,     3,    31,    48,    24,    -7,   -29,   -62,   -29,     5,   -65,   -82,   -59,    13,    16,    71,    11,    14,    24,   -22,    19,    71,   179,   207,   144,   136,    43,    56,    59,    49,    -3,   -50,   -83,   -62,   -62,     7,     7,    15,    16,  -137,   -52,   -27,   -31,    45,   -20,   -75,   -35,   -32,    -5,    60,   192,   193,   111,   117,    38,   113,    62,    94,    38,   -61,  -129,  -133,   -55,   -14,   -35,    11,   -28,  -128,  -109,   -33,   -64,    80,    29,    56,   -53,    66,    45,    89,    92,   166,   118,    12,    56,   114,   100,   147,     6,   -36,   -72,  -171,  -124,   -32,   -49,   -10,     2,  -120,   -22,   -51,  -109,    84,   105,   -21,    35,    12,   135,    97,    62,   152,    55,    26,    62,    90,    61,   102,    -5,   -28,   -72,  -164,   -64,   -98,   -37,    53,   -11,  -125,   -52,  -124,  -131,    98,   119,   113,    75,    54,    21,   -10,    27,    22,    37,    11,   158,    63,   105,    71,   -46,    -9,  -102,  -193,   -92,  -100,   -97,     0,    -3,  -167,   -41,  -146,  -132,    59,   118,    81,    92,    51,    26,   -27,     8,   -71,    14,   134,    97,    56,     9,     5,     6,    41,   -15,   -52,   -34,   -47,   -40,     5,   -19,  -153,   -61,  -146,   -90,   -70,    26,    90,    21,   -41,     7,    39,   -39,   -73,   -23,    58,    32,    -3,     3,   -19,   -46,   -42,     2,   -18,    50,   -54,    10,     3,     9,  -140,   -60,  -120,    -8,   -50,    13,   -78,   -30,   -58,    12,    33,   -64,   -70,    60,     7,     4,   -84,   -60,   -31,   -39,   -71,   -30,    33,    -3,  -126,     1,   -12,    -2,   -98,    77,   -79,  -120,   -37,   -59,   -59,   -24,   -23,    11,    16,  -105,   -29,    17,   -93,  -104,  -117,   -60,   -53,  -114,   -80,   -64,    26,   -90,   -36,    -7,     0,    10,   -67,    23,   -50,   -74,   -17,   -97,  -110,  -101,   -95,   -10,    30,   -12,    11,   -60,  -116,   -88,   -85,   -71,    76,   -77,   -86,  -115,    17,   -25,   -69,   -10,   -15,    13,   -88,  -118,   -35,    26,   -98,   -92,   -42,   -46,   -39,   -37,    12,     1,   -52,  -140,  -112,   -71,   -91,   -84,   -51,   -48,     0,   -48,     3,   -12,    -8,   -11,    -6,    11,    68,   -42,   -20,   -32,  -107,  -158,   -92,     4,   -61,   -53,     0,   -36,   -40,  -135,    13,   -37,   -27,   -85,   -52,   -50,    -3,    70,   -35,     3,   -25,     6,   -16,   -11,    -5,   115,   -54,  -116,   -84,   -95,   -75,   -62,   -71,    -2,    16,    -8,     0,   -31,    90,    58,    50,  -109,    -7,    19,   -16,    18,    18,    14,    16,   -12,    20,   -10,   -11,   -13,   -11,   -31,    53,    67,    31,    43,    27,    11,     4,    79,    34,   -25,   -17,   -68,    -2,     3,   -34,   -69,   -28,   -68,     1,    -3,    -2,   -10),
		    30 => (   18,   -18,    -8,    -3,   -13,    -9,    15,     7,     1,     4,    -1,   -15,    10,    -4,   -35,    -2,     0,    -6,   -12,    -8,   -19,    -5,   -15,    10,     6,    19,   -19,    16,   -19,   -12,     0,     1,    15,    -2,   -11,   -87,   -78,  -126,   -80,    63,    27,    19,   -52,    81,   111,    83,   -47,   -26,   -14,   -26,   -24,   -14,    -3,     6,    -6,     5,     1,    -3,    11,   115,   102,     2,   -15,   -14,   -77,  -100,  -150,  -194,  -110,  -165,  -142,  -245,  -209,  -227,  -146,  -123,  -111,   -96,  -136,   -82,   -45,   -43,    -1,   -10,    10,    11,     3,    71,   -37,   -73,   -68,  -116,  -107,   -37,  -129,    21,    67,    88,   -49,  -166,   -57,   -39,  -147,  -200,   -50,   -88,   -80,   -88,  -114,   -15,   -61,    -5,    15,    -8,   -66,  -136,   -30,  -170,    20,     4,   -21,    13,    38,   -14,    25,    20,   -63,   -72,  -141,    -6,    -1,    62,     6,    -5,   -49,   -89,  -163,  -193,   -79,   -14,   -18,    -8,   -32,   -99,   -22,   -38,    63,    39,    -4,   -52,    36,   -32,  -106,  -107,   -40,   -73,   -93,   -21,    43,    46,   -71,   -68,    12,  -118,   -10,  -243,  -148,   -17,   -13,     2,   -25,    -6,   -26,    -1,     8,    65,    35,  -171,    -5,   -59,  -121,    16,   -38,   -24,   -39,    -8,    -1,    17,   -45,     2,    35,    -6,    51,  -205,   -58,    -9,    16,   -44,    -5,   -63,   -17,   -20,    -2,    -1,   -87,     6,   -19,   101,   -31,    74,   -10,   -57,    24,    -5,    55,    83,    30,   101,    56,   134,    27,    -3,  -127,     0,   170,  -128,    84,    23,   -51,  -138,  -109,   -51,   -25,    -3,    90,     0,    34,   -16,    13,   114,   103,   123,    27,   101,   105,   101,   102,     7,    13,  -105,  -182,   -60,   -15,    -8,   137,  -101,   -94,   -62,   -77,   -93,    -7,    45,    29,     4,    -3,   -11,    60,    48,    70,    50,   -52,    18,   132,    61,   -16,     3,    34,  -151,   -82,   -24,   -34,   -24,   120,    61,  -121,   -64,    50,    -5,   -18,   -17,    15,   -35,   -47,   -27,     3,    90,    40,    96,    12,    -3,    49,    54,    18,   -81,   -68,  -158,  -199,   -12,   -13,   136,  -103,   -27,  -224,     5,    35,    30,    35,   -65,   -45,   -97,   -86,    16,   -50,   -73,   -43,   -38,   -51,   -62,     7,   112,    25,  -128,  -166,  -156,  -130,   -16,    -5,    24,   -92,   -24,   -45,    24,    75,    56,    -6,    31,   -21,  -125,   -47,   -25,  -125,   -70,   -23,   -47,   -58,   -39,    -6,    76,    92,     0,   -86,   -42,   -72,   -53,   -12,    33,     0,    68,   102,    37,   144,    81,     4,    64,     0,   -72,   -28,  -109,   -50,  -120,   -34,    54,    16,    36,  -109,    43,     3,    -6,   -94,   -42,   -86,   -85,    10,     1,    -7,   -19,   171,   192,   196,    91,    67,    91,   103,    36,     0,   -80,   -94,   -13,   -97,    -9,     9,    51,   -39,  -130,    -3,   -57,    49,  -125,  -172,    -1,     5,    -2,   -80,   -65,   123,   219,    60,   127,   146,   212,   127,   -41,   104,   -71,   -73,   -40,   -61,     3,   -14,   -43,   -16,   -91,    14,    30,    -6,   -96,  -187,   -92,   -13,    -5,   -47,  -150,   134,   140,    87,    89,   172,   186,    74,   149,   108,   -63,    21,    42,   -55,   -35,    -5,   -60,   -43,  -110,  -126,    72,  -136,  -207,  -264,   142,    10,   -11,   -46,  -192,    52,    55,   -37,    79,    42,    83,   116,   123,     4,   -62,   -28,   -18,   -11,    10,     8,     5,     2,  -127,    38,   -41,  -140,  -154,  -136,   199,   -15,   -14,   -31,  -214,     0,   -27,   -27,     5,    89,    41,    62,    13,    49,   -12,   -16,     8,   -37,   -67,   -58,   -52,   -55,   -50,     2,   -48,   -68,  -124,  -137,   -49,     4,    48,   -54,  -150,   -68,   -23,   -30,   -19,   -34,  -111,   -57,   -19,    88,    20,   -11,     0,   -43,   -84,   -24,     4,   -59,     5,    11,   -65,   -60,  -215,  -116,   -49,     5,    71,   -50,  -179,   -45,    -9,   -31,   -67,  -101,  -122,   -43,    34,   -19,    27,    77,    38,   -14,   -59,    -3,   -58,   -52,   -37,   -36,   -44,   -76,  -194,     1,   -17,   -15,    12,  -154,  -104,  -112,   -27,    59,    20,   -50,   -51,   -36,   -29,    40,   113,    85,   103,    95,    25,   -44,  -133,  -111,   -45,    14,   -43,   -57,   -55,   126,    43,    -2,    12,  -210,   -65,  -197,   -63,     0,    39,   122,    -8,    49,    48,   167,    67,   131,   112,    14,   -11,   -60,   -70,     7,    42,    71,    76,   -86,   -55,    74,    36,     6,   -13,   -52,  -211,  -169,   -41,    43,   -29,    -3,   -47,    25,    26,    43,    45,    78,    18,    64,   -61,   -56,   -52,   -47,    50,   -32,   -71,   -88,   -62,  -155,     1,    -9,     2,   -22,   -47,   -27,    64,   -55,   -94,  -117,  -186,  -180,  -117,    47,   137,   129,   115,   105,   -14,   -47,  -189,  -134,   -60,   -95,  -113,   -64,     4,   -13,    18,    10,    16,    -2,   -62,  -328,  -261,   -62,   -23,   -25,  -207,  -161,  -109,   -16,   -46,   -61,   -95,   -29,   -14,  -129,  -212,  -157,  -148,   -85,   -38,     8,    -5,    13,    -8,     5,     4,    14,    -8,  -167,  -144,  -208,   -71,  -100,  -166,  -156,   -82,   -92,   -99,  -171,  -140,   -99,  -229,  -225,  -104,  -141,  -157,   -72,   -88,   -29,   -11,    -2,    -7,     4,   -20,     5,    -8,     7,     2,   -21,   -13,   -61,   -39,    12,    10,     9,   -55,    -2,     3,   -34,   -36,   -51,   -50,   -22,   -74,   -78,   -67,    -7,    13,   -17,    19),
		    31 => (   14,   -17,    -7,    -9,     3,   -16,     8,    11,   -10,   -12,     8,   -18,     9,    19,   -12,    13,   -17,   -18,    17,    -5,    -4,   -20,   -16,   -16,     4,    12,    13,    19,    -8,    -6,    10,    13,    12,   -13,    -8,   -19,    -8,     1,   -27,   -27,   -23,   -78,    35,    42,     5,   -45,   -23,    11,    -9,     9,    -2,     2,    17,    20,    10,    -7,   -17,   -14,    -6,     0,   -17,     8,   -14,    17,   -60,   -95,   -64,   -64,  -129,    49,   -32,    -8,    45,    11,    29,   105,   103,  -177,  -146,   -87,   -31,   -37,    18,   -17,     3,    -4,    84,    64,    -2,   -84,  -118,    59,    89,    89,   -10,  -118,   -50,   -68,     6,    85,    14,    -3,    -5,    93,    77,   -43,   -15,   -53,   -81,   -18,   -19,     3,   -10,   -13,    96,    81,    65,   101,     0,     6,    58,    18,    68,   -10,    -8,    54,    -8,   -10,     8,   103,   141,    97,   -13,   -20,    17,   -14,   -54,  -101,  -130,   -93,    14,    17,    48,    28,   106,   124,    91,    97,   -41,   -96,   -40,   -46,    -5,   -17,   -60,    -4,   -30,   -38,     6,   103,    44,   -33,   -32,    61,   -34,  -141,  -101,   -96,     7,   -17,   -83,    31,   118,   102,   115,    78,   -48,   -55,    -7,   -27,   -73,   -44,   -50,   -71,    18,     3,    20,    40,    27,   -66,   -63,     5,    -9,   -60,  -140,   -16,     6,   -50,  -135,   -53,  -189,    15,   103,   113,   -74,   -53,   -67,   -26,     7,    36,    35,     9,    12,   -90,   -11,    40,    40,   -27,    -3,    72,   -23,  -116,  -255,  -147,     5,  -130,  -145,  -184,  -178,   -78,    39,    -2,   -89,   -62,   -10,   -17,   102,    88,   108,   -14,   -23,   -41,    37,    15,   -80,   -42,    54,    11,   -24,  -103,  -356,   -71,    14,   -39,  -118,  -202,  -162,   -82,  -103,   -42,   -92,   -69,   -19,    29,   119,   125,    86,   -32,    -4,   -44,     4,    18,   -58,  -112,     4,   -41,   -90,  -102,  -159,   -89,    -1,   -35,  -115,   -57,  -153,  -116,  -116,   -62,   -81,  -143,   -76,   -38,   144,   125,    74,   -12,   -26,    37,   -43,   -58,   -74,   -83,  -111,  -115,   -99,   -67,   -53,   -21,   -14,    24,   -11,   -89,   -96,  -122,  -161,  -151,  -142,   -98,  -113,   -92,     1,   106,    38,    62,   -50,   -24,   -38,   -77,    15,   -69,   -39,  -135,  -136,   -74,   -80,   106,    -3,   -18,  -169,   -52,   -23,  -104,   -95,  -204,  -142,  -116,   -60,   -58,    11,   112,   -24,     5,    78,    16,   -38,   -35,    40,  -100,   -97,   -56,   -98,   -28,    15,    91,    10,     6,  -144,    47,   -44,  -122,   -68,  -120,   -95,   -75,   -65,   -91,     4,   -16,    41,    47,   123,    87,   -10,   -34,   -36,  -181,  -142,  -137,  -132,    16,    15,    -9,   -19,    -5,    36,    15,   -69,   -82,  -101,   -66,   -94,   -55,  -100,   -88,    29,   -20,     8,    33,    27,    22,   -44,  -113,   -37,  -127,   -98,   -73,   -99,   -94,   -36,   -11,     4,     1,    23,   -69,  -133,  -109,  -112,  -129,   -89,   -17,   -20,   -13,    -6,    42,    35,    13,    52,    49,    25,   -53,  -112,  -207,  -176,  -135,  -338,  -166,   -92,   -63,   -15,    -2,    40,  -144,  -128,   -13,   -49,   -90,   -50,    28,   -38,   -55,   -28,    17,    13,   -10,    49,    -2,   -24,   -28,   -82,  -145,   -81,   -62,    28,  -108,   -65,   -80,    17,     1,   -55,  -153,   -71,   -49,   -85,  -157,    28,     5,    52,    57,   -48,   -45,    95,    73,    57,    27,    -8,    -3,   -34,    47,    42,   -28,    36,   -57,   -88,   -87,   -11,    10,    14,  -174,  -110,  -112,  -235,  -155,    -4,    66,    75,   -36,   -91,   -53,    27,   117,    95,   -35,    26,  -115,   -62,   -31,   -26,    33,    36,   -10,   -79,     6,   -19,    -3,   -34,  -181,  -202,    10,     8,   -10,    60,    85,    82,   -27,   -54,    28,    48,    44,    43,   -46,   -64,  -137,  -104,    -2,    76,    78,   104,    46,  -100,   -23,   -13,     9,   -67,  -184,   -35,   102,   120,   163,    30,   108,    97,    10,    50,    69,    41,    27,    27,   -67,    27,   -33,    34,    51,   102,    88,   101,    12,   -33,     1,    57,    37,   -24,    -9,   -34,    59,    87,   111,   149,   149,    69,     3,    60,   133,     4,   -56,    23,   -44,    23,   -10,    54,    70,    80,    19,    24,    45,   -64,    10,    27,    33,   -52,   -18,   -23,    92,   107,   109,    89,   143,    68,    62,    59,   123,  -125,   -83,   -16,   -30,    21,    56,   104,    74,   -75,   -32,    57,     4,    13,     2,     4,    10,   -27,   -27,   -48,    33,    33,     4,    33,   147,    87,    80,    93,    -7,  -108,   -60,   -92,    37,   -36,   -31,    47,     6,   -33,   -90,  -104,   -78,   127,   -19,     6,   -14,    19,   -23,   -82,    10,   -40,    13,   -27,    50,    44,  -104,   -29,   -10,  -119,  -112,  -111,    22,   -24,  -106,   -37,    54,   -13,  -130,  -128,    12,    21,    19,   -19,     4,     0,   -31,   -90,  -148,   -85,  -200,    17,   -82,   -20,   -87,    66,    -3,  -103,  -126,  -148,  -205,  -234,  -177,  -325,  -118,   -78,   -57,   -28,   -32,   -37,    -5,    -4,   -13,    -5,   -26,  -102,  -216,  -306,  -331,  -231,  -214,    33,     7,  -131,  -130,  -125,  -132,   -86,  -169,   -88,   -27,   -59,   -65,   -16,   -22,    -3,    -6,    -9,    14,   -17,    -4,    -4,    12,   -14,   -26,    -2,    15,    10,   -17,  -126,  -104,    10,   -30,   -93,   -35,   -40,   -10,     2,     2,    18,   -17,   -10,    15,     6,   -18,    14,    18),
		    32 => (   -1,    15,     5,   -12,    -9,    -3,     2,     9,     2,    -8,    -5,   -17,   -40,   -30,    19,     1,    -1,   -16,    -4,     1,   -11,    13,    15,    -6,     6,    10,    14,     7,     0,   -17,    -6,    18,    -3,    -2,    15,     6,   -78,   -50,   -41,   -18,   -31,   -34,  -121,     6,    18,   -31,   -17,   -96,   -48,   -30,   -53,    -5,    17,   -20,    -8,    -5,     9,   -14,    -6,   -21,   -25,    -9,    -9,   -59,   -24,    19,    27,   -27,    20,   -28,   -18,   -47,   -59,   -74,    25,    -6,   -82,   -32,   -28,     5,    -2,    32,    18,     2,   -11,   -19,    -9,   -35,   -68,    53,    35,    27,   -58,   -56,  -104,   -61,  -114,  -145,   -87,   -45,  -149,  -179,  -124,   -37,  -117,  -123,   -46,   -12,    -3,    -9,     7,    -9,   -20,   -11,   -35,   -28,    75,    90,   122,    93,    97,    68,     2,    26,    45,   -50,   -58,   -30,   -29,  -111,   -36,   -18,   -91,   -86,  -121,   -58,   -43,   -30,   -58,    -3,   -15,   -20,    26,    23,    32,    -7,    26,    22,    45,    76,    49,    44,   -17,   -66,   -96,  -132,   -29,   -18,   -76,   -61,   -51,   -30,   -87,   -64,   -12,     4,   -42,   -39,    10,    -6,   -49,    76,    72,    74,   118,    -6,   -25,     5,    -8,    11,   -50,   -40,   -49,   -53,   -10,    -1,    -8,     3,   -70,   -31,   -23,   -82,   -33,   -60,   -32,    -2,    11,    -2,    13,   117,   119,    41,   118,    56,   114,    -8,   -51,    -6,    56,   -17,   -83,   -27,   -23,   -77,    -3,   -28,   -38,   -35,   -67,  -174,  -108,   -53,   -68,   -27,   -49,    29,     4,    44,    59,    40,   102,    80,    57,    65,    21,   -17,    51,   -28,    53,   -28,  -124,   -52,   -76,   -28,   -39,  -104,     6,   -62,  -122,   -67,  -103,   -37,    16,   -24,   -14,   -33,     9,    61,    17,    22,   -22,   -38,  -128,   -72,   -49,   -57,    21,     7,   -31,   -88,   -32,   -10,    -4,   -26,    27,   -31,  -109,   -54,    31,   -10,     0,   -18,     9,  -118,   -63,    -3,    49,     4,   -35,  -110,   -92,  -212,  -203,   -91,   -18,     1,   -29,   -41,   -33,   -30,    35,   -70,   -77,    -6,   -47,   -44,   -53,    -9,    18,   -18,   -50,   -71,   -87,   -72,   -23,   -30,   -40,  -108,   -28,   -59,  -191,   -96,   -50,   -26,    -7,   -66,   -44,   -10,   -32,   -71,    -8,   -35,    -4,    11,  -133,   -30,    10,    -6,   -17,     5,  -108,  -194,  -142,  -125,  -107,  -107,   -71,   -30,   -63,  -101,   -56,  -101,   -43,   -19,   -71,     4,   -55,   -44,    59,    19,   116,    35,   -22,   -20,   -15,     0,    -7,   -31,   -31,  -181,  -220,  -193,  -136,  -129,   -84,     9,    -7,   -19,   -41,  -118,   -70,   -80,   -54,    -2,    45,   -25,    84,   120,   166,    94,    11,   -38,    19,   -38,   -38,   -22,   -84,  -150,  -217,  -152,  -120,   -68,    61,    26,   -48,  -103,   -13,   -62,   -84,  -123,   -30,    96,    14,    27,    80,    52,    36,    18,    47,    78,    19,   -52,    59,    54,   -63,  -142,  -122,   -24,    -3,    30,    68,   -12,    29,    67,    57,     5,   -34,    17,    24,   157,   121,    62,    11,    74,   103,    98,    70,   120,   -10,   -26,    75,    10,   -51,  -151,   -21,     9,     2,     4,    29,    15,    19,     9,     0,   -36,  -110,    16,    88,   126,    24,    86,    91,    99,    25,   160,    48,    59,    16,   -17,   104,   -24,   -84,   -33,    29,    78,    42,    95,    -9,     0,   -63,   -60,    37,   -24,  -132,    79,   126,   -24,   -11,    56,   -19,   -14,  -107,    95,   -15,    72,     6,    14,    20,    81,  -118,    11,    54,    44,    44,   -18,   -59,   -41,    18,   -72,     7,   -46,    38,   102,    69,   -71,   -92,   -31,   -51,   -46,    44,   121,    18,   170,   -14,   -80,   -48,   -39,  -118,     2,    29,    80,    26,   -46,   -65,   -11,   -35,     4,   -37,    -7,    67,    82,     8,   -62,   -99,  -120,    15,   -72,  -109,     5,   111,   128,   -18,   -74,    -6,   -11,   -84,     0,    46,    44,    35,   -62,   -86,     4,    14,    55,   -43,    -4,    21,   -21,   -20,   -65,   -94,   -97,   -74,   -92,  -133,   -18,    23,    10,    -1,    20,    26,    17,  -125,   -76,   -24,   -73,    48,   -19,   -26,    24,    -1,    25,    -4,    55,    76,     3,    14,   -50,     1,    15,   -53,    13,   -79,   -19,    34,   -20,    -3,    11,    -9,    54,   -95,  -151,   -76,   -80,   -63,   -61,   -34,    75,    16,    92,    82,    -7,     3,    30,    -5,   -46,    20,     7,  -100,    10,     7,   -13,   -54,     0,     2,     6,   -12,    66,   -93,  -135,   -94,   -69,   -69,     6,    43,    36,   114,    71,    16,    13,    33,    53,   -41,   -35,   -44,   -24,    23,    40,    23,    39,   -63,     4,     4,     9,   -99,   -76,  -154,  -104,  -137,   -56,  -101,  -131,  -117,   -90,   -82,   -89,   -33,   -43,  -120,   -31,    16,    39,    24,   -43,    -4,    39,    65,    -9,     9,     8,    -7,   -12,     7,    -9,   -29,   -28,   -24,   -15,   -64,  -144,  -197,  -145,  -136,  -244,   -20,   -15,   -70,     5,   -41,    55,    58,    43,   -57,   -15,    23,    19,    13,    -1,     8,   -17,    11,   -11,    -6,   -68,   -65,   -57,   -53,  -118,   -21,   -33,   -63,   -60,   -83,   -54,  -105,  -133,  -106,   -62,   -59,   -45,   -64,     8,     2,     3,   -11,     2,   -20,     7,    14,   -18,   -17,     6,    11,    -4,   -20,    -3,   -42,   -33,   -41,   -74,   -57,    15,    -1,   -34,   -18,   -18,   -26,   -56,   -51,    -4,    19,    -3,   -10,    19),
		    33 => (  -15,    -5,    -1,    17,    10,    15,     2,    16,    14,    -9,    14,    -1,     2,   -13,   -21,     2,     7,   -19,   -18,     8,    11,    17,   -16,     6,     3,   -13,     3,    -7,     0,    10,    -7,   -16,   -17,    -5,     3,     5,    15,   -19,   -22,    -5,   -16,   -25,   -17,   -18,    -8,   -36,   -12,    16,     1,     0,    -4,    13,    -9,    -9,    14,     1,   -20,     7,    -1,     4,     1,    15,   -14,    -4,   -50,   -65,   -26,   -27,   -77,   -70,  -118,    -2,   -40,   -23,   -40,   -33,   -68,   -29,   -33,   -41,     1,    12,   -19,   -17,     8,    20,    -3,   -12,     5,     6,    10,   -11,    -6,    -3,     8,     5,    -5,     1,     7,   -21,   -48,   -39,   -23,   -47,   -17,   -11,   -15,   -51,   -62,   -44,    -8,     0,   -11,    -6,     2,    61,   -19,   -16,    -7,    -7,   -18,    -4,    -2,     3,   -34,   -32,   -19,   -21,    -4,    -9,   -52,   -33,   -48,   -28,    -7,    -2,  -133,   -64,   -37,     8,     4,    -1,    -3,    25,    61,    -8,    20,   -14,   -43,   -69,   -56,   -63,   -77,   -27,   -68,   -24,     5,    52,    65,    42,     2,   -36,   -49,   -39,   -32,  -109,   -28,     4,    -5,   -11,    49,   -19,    48,    46,    17,    17,    -7,    12,    27,    13,    36,   -22,   -34,   -34,   -60,   -86,     9,    20,   -24,   -80,   -66,   -46,    -7,    -8,   -75,   -14,     2,    16,    84,     7,   -23,    45,     6,    50,    48,    53,    16,    46,    -4,   -56,   -41,   -74,   -67,   -30,   -61,  -137,   -76,   -55,   -57,   -55,   -43,   -22,  -112,   -26,   -19,    29,    75,    62,    44,    -8,    55,    63,    54,   -34,    18,   -38,   -61,    -9,    21,    28,    -5,    37,     7,    -1,   -67,   -39,   -21,   -13,   -21,   -57,   -92,     4,    15,   -83,   173,    40,    52,    -3,    92,    35,     1,    51,    40,   -78,   -55,     9,    58,    -8,  -112,    16,    45,   -12,     1,    39,   -47,     0,   -99,  -105,   -46,    -1,    18,   -70,   156,    46,   -20,   -46,    45,     0,   -52,   -95,   -71,   -63,     0,    11,    82,   -81,  -104,   -21,    21,   -22,    22,    33,   -12,   -13,   -87,   -40,   -10,   -10,     5,   -11,   -65,   -52,   -28,   -58,   -98,   -80,   -98,  -116,   -45,     2,    27,   -42,   -76,   -75,   -16,    -7,    22,     5,    19,    31,    30,   -20,   -42,   -89,   -30,     2,    18,     3,   -77,   -34,   -34,   -96,  -116,    -5,   -25,   -36,   -18,    -1,   -45,  -143,   -63,    -4,    -7,    43,    47,   -15,    -5,     8,    -1,   -29,   -34,    13,     2,   -15,     8,     9,   -50,   -30,    -9,   -49,   -69,     0,    16,    22,   -47,     6,   -41,    31,   -16,   -16,   -34,    46,   -28,   -31,   -66,    -1,    17,   -32,   -48,   -40,   -52,   -39,    -7,    53,   -23,   -38,     6,   -11,   -33,   -72,   -38,   -51,    -3,   -17,   -53,    18,    54,    36,    14,   -57,   -90,   -54,   -80,   -30,   -30,   -13,   -35,  -112,   -56,   -40,   -10,    24,   -19,   -46,    38,   -49,   -49,   -22,     3,   -35,    -3,    -2,    12,    25,    30,   -31,     8,    -6,   -53,   -81,   -41,   -40,    39,    -2,   -28,     0,   -16,     0,   -12,     1,   -25,   -34,     5,   -47,   -12,   -41,   -13,    75,    13,   -19,   -20,    10,     6,   -32,     3,   -77,    -9,     0,   -23,    -5,    38,     2,   -23,    13,   -79,   -53,   -17,    26,   -17,    65,     9,   -16,    -6,   -26,     3,    58,   -16,    30,    26,   -17,   -31,     6,   -21,   -90,   -80,   -47,   -26,    -4,    40,    -6,   -50,   -21,    -9,   -24,   -29,     7,     5,    50,    51,    38,    -2,   -60,    -3,    47,    97,   -16,    16,    76,   -12,   -30,   -37,   -85,   -85,   -43,   -16,    42,    66,    18,   -41,   -31,   -12,   -43,   -19,    -8,    16,    13,    64,    41,    13,   -27,   -16,    -7,    37,   -36,    33,     9,   -46,   -31,   -56,   -49,   -51,   -46,    27,    23,    88,    68,   -48,   -22,   -35,   -28,    -6,     5,   -18,    21,    24,    28,    39,   -25,   -51,    14,    -7,  -111,   -11,    53,    -2,   -55,   -14,   -31,   -49,    11,   -22,    31,    82,    68,   -69,   -57,     2,   -21,    -1,     1,     8,    35,    41,    11,   -10,   -68,   -99,   -20,   -51,  -104,  -103,   -67,   -90,   -20,    28,   -41,   -11,     8,    -5,     6,     3,    68,   -50,   -54,    -4,    14,   -27,     1,     7,    27,    74,    18,    -2,   -42,  -102,   -54,   -40,  -112,  -150,   -87,  -136,   -95,   -38,   -30,    74,    92,    38,   -36,    -7,    67,   -20,   -49,   -15,    15,     5,    12,    43,   -21,   -14,   -25,   -19,   -22,   -63,  -109,   -31,   -24,   -76,   -69,   -89,   -15,    61,    25,    42,   -36,     5,    18,    35,     6,   -38,   -55,    16,   -19,    -5,    -2,   -38,    -2,   -32,   -31,   -22,    29,   -61,   -77,  -100,   -16,  -115,   -40,    53,   126,    77,     2,   -38,   -23,     6,   -16,   -45,    29,   -78,   -40,   -22,   -10,    -2,     2,    30,   -34,   -88,   -96,   -31,    13,    54,     0,   -34,   -31,    22,   124,   178,    28,    55,   -44,    -7,     6,    46,    -3,   -73,  -187,   -13,    -1,     3,     5,     4,    12,    -9,   -66,   -71,   -70,  -115,   -82,   -77,  -120,   -64,   -55,    68,   121,    86,   -16,   -42,   -37,   -33,   -43,   -65,   -50,   -99,    16,    15,    -4,    -5,    16,     1,    17,    -4,    19,     4,     3,   -21,    17,    16,   -68,   -67,   -27,   -38,   -37,   -30,   -70,    -2,     7,   -25,   -16,   -36,   -40,    -5,    -4,     5,     4,    14,     0),
		    34 => (  -15,   -12,   -10,     7,     1,     4,   -17,    13,    -5,    17,   -19,   -11,    -4,   -13,     5,    14,     7,    16,    -3,     8,    -9,   -11,    -5,    -1,    13,   -14,   -12,    13,   -15,   -18,    19,    19,     9,     0,   -20,   -40,   -38,    10,   -18,     6,    11,   -76,   -61,   -17,   -12,   -32,     3,    10,    -6,   -17,   -27,   -16,     1,   -15,   -11,     1,    17,   -12,   -16,   -15,   -45,     6,   -34,   -63,   -28,   -12,   -34,   -35,   -14,   -47,   -60,   -27,   -16,   -52,   -12,    -5,   -59,   -22,   -22,   -13,    10,    -2,     3,    17,    13,   -12,    -5,   -18,   -25,   -21,   -91,   -46,   -72,   -38,   -15,   -27,   -35,   -70,  -114,  -114,   -71,    26,    -4,   -48,   -23,    -4,   -14,   -14,     4,   -22,    -2,    -6,     9,    -6,    -3,   -25,   -38,   -11,   -41,   -34,   -13,   -26,   -35,   -38,   -49,   -93,  -132,   -68,   -37,   -43,  -105,   -85,   -18,   -64,   -79,   -19,    22,    -9,   -18,   -23,     9,    19,    14,   -22,   -29,    -6,   -39,   -15,   -50,   -62,   -18,   -81,  -129,   -77,    -1,    52,   -27,  -164,  -146,     5,   -51,   -23,   -31,    59,    67,     8,   -59,   -14,   -11,    -3,    14,   -49,   -31,    65,   -51,   -10,   -52,   -48,   -76,   -52,   -24,     1,   119,     6,  -246,  -295,   -96,    16,   110,     4,    69,   -63,    26,   -25,    65,  -104,   -19,  -110,     2,   -15,   -22,    94,   -20,   -15,    13,   -47,  -128,   -75,    50,    43,    45,  -200,  -264,  -204,   -34,    55,    25,   -13,    64,    44,    28,    27,     4,   -55,   -37,   -97,    25,   -17,   -15,    13,    13,    53,    -7,   -38,  -135,    18,    62,    73,   -92,  -110,  -225,   -57,    15,     8,    28,   -10,    60,    20,    45,    -8,   -36,   -82,    14,   -81,    33,   -19,     8,   -38,   -63,   -25,   -66,   -92,   -78,    97,    11,    -4,   -58,  -199,  -151,   -17,    28,    52,    35,     7,    22,    12,    15,   -43,    -7,   -41,   -18,   -13,   -62,    -6,    -6,   -95,   -81,   -19,   -83,   -88,   -19,    98,    -2,   -67,  -131,   -63,   -44,   -31,   -20,     5,   -19,   -94,  -142,    10,   -94,    -6,   -35,   -36,   -14,    -9,   -66,   -39,   -63,   -71,   -43,   -86,   -18,   -31,    26,    49,     3,   -50,    -5,    58,   -32,     5,    -1,    74,   -38,   -42,   -79,  -100,   -65,   -29,   -72,   -96,    18,     1,  -115,   -79,  -117,   -59,   -87,   -49,   -57,     8,    42,   -27,     5,    -1,    25,   -25,     7,   -28,   -28,    14,   -21,    37,   -41,   -87,   -60,   -54,  -152,  -103,   -18,   -13,   -82,   -75,  -125,   -62,    -2,   -32,    -1,     7,   116,    31,   -35,    29,    50,    50,    59,   -23,   -71,    45,    50,    22,   -81,  -103,   -95,  -130,  -151,   -17,    -8,   -15,   -53,  -119,  -120,   -44,   -54,   -18,   -54,    12,    45,    -9,   -25,    24,   -15,    67,    58,   -67,     7,    43,   101,    36,   -79,   -27,   -60,   -63,   -71,   -10,    -7,     4,   -29,   -22,    19,   -52,   -78,    11,   -16,    19,   -17,   -30,   -19,   -12,    -4,    98,   -52,    -7,   -43,    84,   -66,    14,    -5,    28,   -62,   -42,   -23,    29,   -18,    15,   -32,     3,    -4,    28,   -54,     1,    41,    53,   -50,   -56,   -25,    27,     4,   -13,   -45,   -84,  -141,   -49,   -76,   -62,   -45,    20,    20,     3,   -28,   -17,    19,     8,   -66,   -13,   -41,   -49,     9,   -41,    42,   -17,   -77,   -23,   -50,   -66,   -44,   -12,    45,   -97,  -112,   -88,   -65,   -12,   -27,    31,   -11,     6,     2,   -32,   -23,    14,   -66,    24,    48,     3,   -22,    -7,  -107,  -116,   -87,    -8,   -41,   -38,   -14,   -22,     1,   -98,     0,   -11,    20,     3,   -28,     3,    -9,   -15,    10,   -18,     9,   -76,   -84,    24,    77,   -36,  -102,   -89,  -107,   -63,  -111,     3,    -2,   -33,   -24,   -15,     0,   -67,   -12,    31,     2,   -45,   -65,     2,   -12,    18,     8,   -25,     2,   -17,   -13,   -34,    16,   -61,  -150,   -91,  -147,   -51,   -39,    32,   -50,   -53,   -74,  -119,   -47,   -89,   -44,   -39,   -50,   -50,   -15,    24,    20,   -45,   -20,    12,     5,    15,   -41,   -66,    -5,   -54,  -188,  -117,   -12,    -2,     2,   -33,     0,   -36,   -65,   -77,  -140,   -76,    10,     8,   -44,   -68,    40,    28,    33,  -112,   -32,     5,   -20,    18,    14,   -48,   -59,    -2,   -70,   -99,    10,     7,    28,    69,    15,   -33,   -99,   -38,   -71,   -41,    27,   -61,   -42,    -5,    18,     7,    19,     3,     6,   -18,   -14,    20,   -40,   -31,   -30,   -83,   -56,   -64,    24,   -31,    20,    -1,   -67,  -117,   -72,   -21,   -37,   -25,    84,    55,   -91,    -6,    15,    57,    34,    19,     9,    -1,    13,    13,     1,   -22,   -85,   -45,   -12,   -20,    21,    28,    63,    29,   -91,   -10,   -19,    40,     1,   -39,   100,    89,    58,    33,    50,    41,   -12,    88,    -5,    20,    -3,     0,   -48,    10,   -74,   -18,   -88,   -46,   -86,   -72,    17,    11,    34,    23,    10,   -41,   -73,    -4,    75,    87,    26,    12,    72,    27,    32,   -13,   -17,    18,     4,     1,     7,   -16,   -69,   -15,   -48,   -58,   -60,   -81,    12,   -36,    32,   -26,  -100,   -42,   -12,   -43,  -100,   -47,   -50,  -152,  -139,    -6,   -29,     0,    -2,   -17,    15,    -9,    -6,    18,     9,    -3,   -32,    -9,    -7,   -30,  -123,  -120,   -86,   -74,   -93,   -12,   -51,  -106,   -34,   -70,   -52,   -42,   -33,   -24,   -18,     8,    13,    -7),
		    35 => (   18,    -6,    17,    13,     0,     4,   -11,     4,     5,    14,   -16,    -8,   -16,   -14,    19,    -4,    -3,     8,     8,     2,    -5,   -11,     3,     6,   -10,    16,    17,     5,   -11,     1,    10,    -8,    12,    -2,   -16,    -6,   -12,   -10,     8,   -31,   -26,   -20,   -18,   -37,   -62,   -55,   -21,   -42,    -8,   -26,   -17,   -13,    -3,    -7,   -19,   -10,    15,   -20,   -16,   -29,   -31,    16,   -52,   -45,   -42,   -85,   -99,   -79,  -111,  -102,  -238,  -160,   -94,   -50,   -36,    30,     5,  -111,   -46,    20,   -48,   -34,     5,     6,    15,    13,    -9,     8,   -17,   -99,   -80,   -67,  -157,  -169,  -131,   -33,   -39,   -11,   -34,   -40,   -71,    42,   110,    48,   -67,   -34,   -40,   -66,   -65,   -14,     9,   -16,    -3,     7,   -33,    28,   -62,   -33,  -104,     6,   -35,   -10,    56,   -34,  -106,   -37,    51,    68,   -21,   -50,     8,   -67,   -74,   -38,   -84,  -124,  -140,   -99,   -29,   -20,    -7,    -1,   -21,   -20,   -66,     8,   -58,  -138,  -103,   -56,   -58,   -23,  -103,   -91,   -46,   -94,   -90,  -165,  -178,   -28,    34,   -73,   -77,   -23,   -94,  -123,    40,    24,    -9,    -5,    63,   -92,  -101,    49,   -55,   -78,   -25,   -74,    19,   -32,   -89,   -39,     5,   -48,   -79,   -65,   -27,   -23,    -8,   -14,     2,   -20,    -1,  -114,   -17,     5,    13,   -26,    67,   -48,  -116,    46,  -108,   -49,   -20,   -17,   136,    30,   -41,    -7,    -9,    26,   -86,   -92,  -154,  -160,   -48,   -17,    13,    17,   -49,   -28,    -2,    75,   -17,    -3,   -80,    10,   -39,   -25,   -58,   -11,    -7,    13,    33,    46,   -34,   -33,    48,    40,    56,    43,    -3,    68,    68,    69,   102,   104,    95,    68,   -60,    48,    -4,    -7,   -86,   -60,   -42,  -142,    32,    49,   -12,   -16,   -22,   -74,   -39,   -13,    52,    47,   109,   176,   126,   144,    96,   116,   101,    73,   169,   135,   -97,    18,    -6,   -14,   -18,   -65,    -7,   -29,    39,    33,   -36,    -5,     8,    78,   -45,   -10,    19,    31,    15,    66,   146,   128,   126,   158,   109,    50,   183,   132,    66,    97,    17,   -23,    -9,   -19,    29,     1,   -37,   -90,   -35,   -63,    38,   -22,   -38,   -68,  -141,  -121,  -103,  -108,   -79,  -130,   -89,    24,    16,    63,    19,   154,   137,     9,    -1,   -21,    -9,    17,   -31,   -52,   -68,   -22,    -4,    49,    66,    92,    49,     0,   -69,   -93,  -155,  -134,  -274,  -442,  -280,  -187,  -189,  -112,   -91,    92,   141,   -45,     1,    -2,   -21,    30,   -30,   -95,  -110,    43,     6,   -22,   114,    38,    71,    16,    21,    -2,   -77,    -5,   -97,  -187,  -247,  -156,  -215,  -220,   -78,   -31,    95,   -45,    34,    10,   -25,   -31,    48,    -8,    41,    28,    78,    73,    -5,     7,   -15,   -16,   -22,    -5,   -41,    32,    -2,  -150,  -165,  -125,  -109,   -76,   -80,  -102,   -29,   -19,    22,     4,   -81,    76,   133,    59,    24,   100,    64,    77,   -16,    10,    28,   -11,   -63,   -73,  -122,   -32,    45,    -3,   -69,   -62,  -119,   -51,   -85,    41,   -28,   -60,     3,     6,   -74,    12,    49,   138,   -17,    73,    -3,    45,    -4,   -49,   -41,   -17,  -115,   -47,   -68,   -30,    35,    -1,    -8,   -57,   -46,   -64,   -39,    41,   -72,   -79,    14,   -16,  -138,    20,    36,    36,    25,   -55,   -29,    34,    15,   -22,   -90,   -90,   -83,    -7,   -42,    -7,   -55,    -5,   -45,   -83,   -28,   -26,  -136,  -149,  -141,  -141,   -35,   -21,   -77,  -145,   -68,   -43,     2,   -40,   -48,   -77,  -154,    63,    77,   -41,   -78,    19,   -61,    11,   -37,     5,    44,   -84,   -18,    72,    15,   -52,  -152,   -95,     4,     2,   -21,  -123,    56,    84,   -28,   -51,   -30,  -110,  -135,  -133,    -6,    55,   -88,   -69,   -30,    24,    17,    67,     7,   -96,    32,   126,   122,   141,  -133,  -105,    -4,     5,   -22,   -83,    67,    -2,   -59,   -14,   -59,   -54,   -73,     5,    27,    52,  -167,   -52,    20,    -1,     7,    52,    38,   -71,    24,    20,   145,   163,  -111,    -1,    -2,    15,   -25,   -58,   -30,    42,   -69,   -75,   -23,   -11,    17,    21,    35,    25,   -49,    87,   -26,    -9,   -17,   -11,    25,   -48,   -80,     2,   111,   189,    92,   -18,     1,    -8,   -60,   -12,   -30,    44,    47,   -65,  -102,    -9,    13,    28,    73,    20,    -3,    57,    28,    56,    -2,   -71,    15,   -15,   -68,   130,   219,   217,   215,    18,   -17,    -5,    67,   -15,     0,     3,   -37,   -94,   -87,    55,    88,   -43,    -1,   -57,    22,    31,   -35,   -10,    -6,   -73,     5,   -64,   -10,   206,   217,   195,   253,   -15,    19,   -17,   -15,     1,  -100,  -140,  -103,   -68,   -39,   -55,    12,    32,    69,   -29,    69,   -24,   -22,   -31,   -50,   -43,     8,    58,   141,    73,    55,  -152,   -49,    14,     6,    10,    -8,     8,  -138,  -154,   -92,  -132,  -100,   -55,   -73,    14,   143,    75,   -17,   -86,   -61,   -52,    24,    -3,   -77,    63,    81,   107,   113,   -16,   -24,   -16,    -8,    -1,    -8,     2,   -80,  -168,  -229,  -214,  -202,  -191,  -171,  -116,  -120,  -182,  -291,   -76,   -12,   -45,   -24,    23,    -4,    35,    -5,   -90,   -45,    11,    15,    -4,     9,     8,    16,     9,     1,   -38,   -17,   -47,   -43,   -24,   -13,   -38,   -45,   -33,  -157,   -83,   -34,   -63,   -88,   -58,   -38,   -68,  -148,  -106,   -14,    15,   -11,     1),
		    36 => (    1,    12,     4,    11,     0,    -7,    11,     2,   -16,   -13,   -12,    -6,    24,    12,    -1,    -8,    12,   -15,    -8,    16,    11,     9,    11,   -10,   -13,     3,   -14,    -3,   -15,   -13,    12,   -19,     8,    14,    60,    67,    63,    46,    93,    14,    -5,    42,   -60,     3,    11,    40,    87,    56,   171,    69,    67,    63,    19,     9,    -6,    15,   -13,     5,    54,    32,    86,    75,    85,   107,    62,   -34,   -49,   -64,   -89,   -88,    12,    47,    75,   147,    79,    37,    28,   158,   145,   108,    71,   103,   -19,    -8,    -7,    -4,  -118,    17,   -40,    56,   106,   101,     4,   -48,   -54,  -152,  -203,    -6,    91,    60,   -76,   -50,    26,   -49,   -47,    -7,   -79,    25,  -119,   -60,   -91,   -13,     6,    11,  -161,   -21,    52,   130,    95,   -42,  -104,   -87,  -115,  -199,  -261,  -109,  -138,   -73,    -5,   -55,   -28,   172,   112,    23,  -134,  -152,  -241,  -178,   -68,    49,     3,     1,   -74,   -93,    47,   100,    47,   -34,   -49,   -43,   -70,  -220,  -151,     6,    22,   -75,   -42,    -1,    49,    50,    91,    63,   -47,     6,  -114,  -171,     8,    14,   -18,   -12,    74,    25,    27,    95,    92,   -10,   -29,  -114,  -124,   -87,   -55,   -73,   -60,    88,    63,    19,     7,   -11,     6,     7,    34,   -65,   -52,  -136,   -65,   -19,    -1,   -11,   -11,   -34,   -32,    14,   -44,     4,   -74,  -136,  -232,  -172,   -57,   -68,    38,    60,   -63,   -90,   -31,  -160,    14,   -21,    71,   -87,  -199,  -186,   -38,   -76,     4,     2,   -79,   -62,   -37,    16,    63,   -73,  -114,  -220,  -217,   -35,    -7,   -18,   -25,    26,    -2,   -73,  -188,    -2,   -68,   -84,   -80,  -213,  -184,   -84,   -72,  -100,     5,     0,   -72,   -53,   109,   -33,   -17,   -14,  -120,  -113,   -60,   -10,   -32,    21,    64,    31,   -84,  -143,  -194,  -241,  -297,  -279,  -259,  -237,  -187,  -103,  -110,   -33,    16,    10,   -69,   -35,   -69,   -77,   -95,   -89,  -190,   -52,    23,    -3,    19,    31,     4,   -17,   -81,   -28,   -38,  -168,  -172,  -166,  -211,  -236,  -165,  -137,   -98,   -77,    -8,     4,    18,  -119,   -50,   -18,   -26,   -46,    23,     3,    23,    29,    55,    50,   -22,  -117,  -101,   -44,   -78,   -27,   -47,   -85,     1,  -202,  -209,  -190,  -124,  -106,    18,   -15,   -24,   -82,   -77,   -25,   -14,   -80,    -9,    20,    73,    53,    27,   122,   -42,    14,   -86,    54,   -18,    -3,   -36,   -70,    32,    24,   -84,  -191,  -195,   -98,   -14,     9,   -23,  -100,   -80,   -43,   -77,   -97,    20,    13,    36,   130,    29,    65,     4,    11,   -28,    39,   132,     0,    20,     6,   131,   112,  -111,  -220,  -105,    -4,    -8,     9,   -10,  -123,   -83,    20,  -110,     2,   -37,    48,    74,    24,     2,   -47,   -36,    -6,     3,  -166,    34,    63,    -8,   114,    82,     7,    29,   -78,   -99,     2,     6,    20,     4,  -105,   -13,    26,   -64,    -3,    48,    42,    46,   -89,   -33,   -39,    -2,  -116,   -95,  -120,    32,    89,    45,   138,    51,    22,  -102,  -143,  -173,  -100,     0,    12,    -1,   -39,   -33,    41,   -14,    74,   -22,    51,     7,    53,    88,    66,    54,     1,    30,    -2,     6,   -14,    58,   121,    68,   -13,  -136,  -158,  -165,  -131,     1,    -7,    -9,     6,    23,    39,    10,    24,    92,    -6,    32,    53,   -49,     5,   -31,   -53,   -49,   -19,    -7,     5,    48,   107,   -36,   -31,  -126,  -105,     0,  -134,    -3,   -20,     9,     2,    96,   -25,   -60,   -29,   -21,    97,    61,   -52,   -30,   -44,   -11,   106,   -19,    46,    73,    41,    25,   -23,  -194,  -151,  -114,   -97,   -20,   -55,     2,   -44,   -55,    22,    68,   -69,   -28,     0,   -58,    23,    46,    83,    -6,  -154,   -54,    40,   -14,   -18,    64,   -42,   -34,   -75,  -206,   -82,   -43,   -43,   -70,   -22,   -14,   -49,   -39,  -124,    83,    33,   -27,   -26,   -22,   -49,    21,    77,    75,   -42,   -13,   -26,  -113,   -76,  -110,   -31,    -6,   -13,   -30,   -99,   -53,   -65,   -85,    14,     7,   -14,   -61,   -59,   -55,   -74,    -2,   -21,   -12,    -1,   -34,    83,   -41,   -20,   -43,  -102,   -36,   -60,   -39,   -71,   -26,    15,   -83,   -68,   -66,   -68,   -63,   -16,   -14,    -5,   -23,   -43,   -83,  -111,  -123,   -62,   -77,   -40,     5,    13,    41,    59,    -5,    23,   -37,   -87,   -41,   -75,  -133,  -115,   -30,   -75,  -155,   -70,    15,   -20,    -3,    12,    14,   -22,   -48,   -70,   -79,  -133,   -90,  -115,    -1,    52,    39,    -9,    37,    65,   -79,  -154,    80,   118,    71,   -13,   -11,   -27,   -31,   -17,   -34,   -19,   -18,   -17,     9,    17,   -33,   -11,   -14,   -50,   -83,  -126,  -143,  -145,   -67,   -29,    27,    96,   120,     2,   -13,  -149,   -93,   -28,   -33,    -1,    -9,   -10,    19,    18,    10,    -5,    19,    19,    19,   -14,   -44,   -64,   -42,   -17,   -64,    36,    85,    17,   -14,    -1,   -22,   -18,    -3,   -27,   -65,   -17,    10,     2,   -20,    17,   -10,    18,     7,     1,   -17,   -17,     0,     1,     8,    -3,    -3,    -4,    -9,    -9,    12,   -17,    -2,   -26,   -27,     4,     3,    14,    -2,   -29,     0,   -22,     3,   -11,    15,     3,    10,   -10,    16,     3,     3,     6,    18,   -16,     7,    12,   -22,    -3,   -20,     2,   -21,    -1,     6,   -23,   -23,    10,     6,     5,    11,     2,    19,     3,    16,    -1),
		    37 => (    0,   -17,    -5,    10,     5,     9,    10,     4,    -1,     5,    -4,   -17,     0,   -11,    18,     2,     5,    -7,    -9,   -14,     8,     7,   -16,     5,    11,    16,   -19,   -17,     2,   -19,     6,    10,    -7,     2,    10,   -11,   -13,   -22,    -9,   -67,   -83,   -53,   -39,   -65,   -78,   -64,   -23,     6,    -6,    -3,    17,   -11,     8,    16,   -19,     9,   -16,     9,    -4,   -49,   -49,     2,   -16,   -56,   -98,   -37,   -10,   -85,   -36,    -8,     3,    -8,    -2,   -26,   -23,    12,    -6,     3,     6,   -16,    13,     0,    14,     6,   -18,    18,   -18,   -36,   -29,   -21,   -55,  -145,  -138,   -45,   -78,   -66,   -50,   -60,   -30,   -39,   -40,   -98,   -43,   -68,   -23,   -24,   -35,    -5,   -15,     7,   -19,    -6,   -17,    -3,    14,   -24,   -95,   -74,   -55,   -84,  -154,  -146,  -147,  -169,  -166,   -81,  -147,  -118,   -81,   -77,   -84,   -28,   -46,   -55,   -67,   -66,   -69,   -28,     6,    16,   -10,    15,    12,  -116,  -186,    27,   -58,    52,   168,    53,  -104,  -150,   -86,    62,   -49,   -28,  -180,  -214,  -149,  -224,  -185,   -96,   -97,   -97,   -28,   -87,   -13,   -15,     7,     5,    30,    35,   -17,     6,   -12,   -78,    -2,   -31,  -132,   -77,   -88,  -106,   -42,   -76,  -173,   -16,    46,   -15,     1,   103,     9,   -87,  -135,   -15,  -141,   -43,     7,    25,    27,    58,    52,    20,    48,    68,    10,     0,    17,  -102,   -58,   -32,   -52,  -121,  -101,   -18,     0,  -197,  -113,   -30,   -26,   -56,  -123,   -61,   -62,   -34,   -47,    25,   -71,    15,    62,    78,   128,    47,    14,   110,   -13,    19,    44,    10,   -92,   -54,   -57,   -48,    52,   -93,   -39,     4,   -42,    20,     2,   -63,  -112,   -33,     7,    36,     1,    28,   171,     3,    23,    -6,   -17,    20,   -80,    40,   108,    56,    82,    52,   -64,   -60,   -11,   -39,    12,    83,    69,   144,    27,   -90,   -68,    80,     3,    98,    54,    69,   182,    80,    83,   -68,     8,    59,    -1,    66,    17,    -1,    66,    79,   -17,    -4,   -21,    -5,   -30,   -27,   157,    60,  -115,   -11,   -59,    81,   -11,    60,   153,   130,   160,    27,   -58,   -11,   -48,    -6,    24,    60,    -7,    22,    26,    35,   -66,   -50,   -38,    13,   -78,    49,    51,   -46,  -178,  -150,   -36,   127,    17,    22,    21,   176,    76,    32,   -24,   -25,   -34,   -30,   -21,    16,    15,   -36,    30,    32,    15,   -60,    44,    25,   -16,    66,    89,  -102,   -91,    41,   -36,    95,    20,    64,    74,   160,    65,    43,   -56,   -46,   -90,   -68,    52,    42,   -24,  -111,    37,   -78,     8,   -27,   -33,   -42,   133,    87,    32,   -25,   -12,   105,   -49,   -48,   -27,    37,   165,   165,   -16,    69,   -50,   -90,   -65,   -14,    68,    53,   -73,  -202,   -37,   -42,    -5,    57,     2,    92,    68,    73,    41,   141,   137,   -61,   -74,   -22,   -10,    16,    96,    83,   -67,    11,    23,     3,   -37,    10,    79,     2,  -106,  -123,   -10,   -74,   -72,    23,    22,   140,    52,    25,    86,    63,    50,   -96,   -44,   -35,     2,     3,    40,    26,   113,    40,   -45,    45,    42,   113,    10,   -26,  -196,   -89,   -64,     6,   -30,    10,    13,    55,     5,   118,   168,   150,    64,  -240,  -102,     8,   -20,    -6,   -39,   -10,    66,    31,   -61,     5,    52,    47,   -74,  -103,  -164,  -143,    48,    37,    19,   -28,   -16,   -29,    42,    64,   166,    81,     0,  -231,   -65,  -149,    70,    15,    55,  -175,    -1,    11,   -58,    35,    52,    20,   -63,  -141,  -315,  -117,    90,    64,    16,    -1,   -13,   -68,    19,    46,    85,   -20,  -121,   -56,    -7,   -50,     3,    64,   -21,  -158,   -37,    19,    70,    23,     7,   -30,  -190,  -349,  -290,   -91,   109,     5,   -50,    22,   -68,   -34,   -53,  -150,  -226,  -112,   -89,  -100,    -6,    -9,    -9,    41,   -14,   -34,    33,   105,    78,    78,    11,  -189,  -264,  -360,   -99,   -40,     7,     4,   -22,   -46,   -63,   -78,   -96,  -112,  -163,  -152,   -18,   -79,     7,    11,    -2,   -16,   -19,   -36,   -85,    65,    23,    31,   -98,  -183,  -221,  -180,     1,   -80,    22,    48,    65,   -61,   -67,   -71,  -105,   -55,   -83,  -141,  -141,   -50,   -13,     5,    -2,     5,   -13,   -24,     0,    -6,    22,   -41,  -124,  -116,  -189,   -94,   -29,   -41,    41,     1,     0,    11,    18,    29,    28,   -48,   -77,   -90,   -64,   -56,   -88,    12,   -18,     6,   -40,   -38,    23,    33,   -20,   -51,  -123,  -113,  -164,   -97,    21,   -20,    83,    41,    -9,    11,   101,     4,    -9,   -73,   -85,  -127,    -3,   -38,   -64,   -16,   -12,    13,   -26,    -4,    15,   -15,    -8,   -58,   -99,  -108,  -141,   -65,    24,   -47,    -2,   -24,   -24,    33,    16,    60,    -8,   -14,   -32,  -132,    -5,    -2,   -18,    17,    -3,    10,   -36,    -3,    -8,   -19,    12,   -23,   -77,   -90,  -170,   -84,   -96,   -56,    61,   -20,    75,    70,    51,    74,    21,    15,    34,  -159,    -9,   -49,    10,   -14,    10,    -2,   -19,     3,     5,   -22,    -6,    21,    38,    23,   -32,  -168,  -107,   -54,  -155,   -62,    58,    44,    58,   112,    16,    32,    34,   -33,   -37,    17,    -2,   -12,    -3,   -20,   -19,    10,    10,    52,   -64,   -60,     7,    82,    70,    -1,   -24,  -103,  -125,   -56,    67,    81,    17,   -89,    13,    95,    59,    82,    14,    11,   -10,     5),
		    38 => (   -7,     0,     1,     9,    15,    13,    11,     3,    -6,   -14,    -5,     4,     7,     7,     2,    -8,     6,    17,   -17,     0,   -14,    -8,   -15,     5,    -5,    14,    14,    13,   -15,    16,     2,    19,   -16,    14,   -13,    20,   -17,    10,     9,   -15,    16,   -21,   -35,   -75,   -91,   -46,   -41,    -1,   -35,   -12,   -30,   -18,   -13,    -7,   -18,    10,     5,     9,   -30,   -10,    -1,   -20,    -5,     3,   -35,   -40,   -77,   -65,     9,   -20,     4,   -46,   -26,   -50,   -24,   -15,   -68,   -76,   -94,   -43,   -12,   -35,    -3,   -11,    11,    10,   -31,   -10,    -8,   -69,   -28,  -101,   -97,    10,   -11,   -65,   -61,   -72,     8,    65,    65,    52,    21,   -36,   -46,   -23,   -10,    14,   -14,    -8,   -52,   -12,   -14,   -18,    19,   -41,  -113,   -50,   -11,    -6,    11,   -17,   -33,   -17,   -50,   -69,   -20,    26,    36,    12,    22,    20,    78,    55,   -59,   -30,  -115,   -51,   -17,   -44,   -20,    -6,   -27,   -96,  -111,   -38,    -8,   -35,   -59,   -76,   -68,   -80,   -88,   -88,   -69,    34,   -25,   -20,    40,    52,    59,     8,    -6,   -75,   -42,     0,     4,   -61,    -6,     6,   -42,   -55,    -7,    25,   -47,   -26,   -38,   -83,  -123,  -126,  -101,   -64,    11,    21,     1,    -2,   -27,    56,   -40,    63,    16,     4,   -74,   -17,   -14,    -3,    15,   -73,   -52,   -33,    23,   -11,    -9,     7,    30,   -13,    22,   -27,   -25,    54,    17,    38,   -10,   -59,   -38,   -10,    -7,   -60,    -3,   -23,   -52,    43,    74,    28,   -31,   -46,   -28,    10,     8,    14,     7,    18,   -28,    48,    45,     0,     8,   -10,   112,   100,    24,    11,   -52,     3,   -56,   -31,   -63,   -17,    78,   144,   102,    44,    17,   -40,   -11,    15,   -25,   -36,   -39,   -19,   -85,   -80,   -12,   -55,   -24,    -6,    39,    73,    13,   -70,   -81,     4,   -47,   -15,    20,    90,    95,    93,    36,  -132,     9,   -19,    -1,    -6,   -36,   -48,   -57,   -49,   -48,    24,   -50,  -102,   -84,   -53,    11,   -19,   -27,   -41,  -104,   -54,   -14,    93,    85,    35,     1,  -134,   -71,  -122,    -3,    -8,   -21,   -10,   -30,   -46,   -66,   -40,   -74,   -19,   -21,   -92,   -46,   -49,    37,   -32,    25,   -61,   -21,    23,   -61,   -16,    93,     2,   -40,   -77,    41,   -80,    12,    11,   -11,   -61,   -25,   -61,   -44,   -91,  -119,   -12,    17,    -3,    19,    14,   -19,    41,   -27,    22,    40,    13,    62,    47,    -4,     1,    -7,  -112,   -64,  -125,     4,   -15,   -62,  -106,   -27,   -38,  -123,   -96,   -63,   -47,   -71,   -23,   -42,    27,     7,    12,    39,    74,   -36,   -26,   -75,   -66,    15,    -8,     6,   -55,   -19,    28,    -9,    -7,   -19,  -128,   -48,   -78,    63,    40,   -58,  -163,  -128,    16,    -7,    63,    44,    22,    51,   -62,   -68,  -141,   -40,    15,     9,    22,     0,    10,   -35,   -44,   -19,   -17,    -1,   -16,   -34,   -15,   116,    44,   -72,   -72,   -21,    38,    52,    38,     4,   -19,   -14,   -87,  -160,   -76,   -50,   -18,     9,   -68,   -80,     7,   -62,   -38,    13,    -8,   -27,   -37,   -25,    41,    58,    14,    35,    82,    51,    66,    28,   -69,  -109,   -82,    -7,  -117,  -176,  -112,   -75,   -29,   -54,   -94,   -73,    -2,  -117,   -55,    13,   -31,    -5,   -27,    -8,    36,   100,   167,   128,    95,    63,    -1,   -87,   -54,   -80,   -54,  -101,   -13,   -85,   -62,   -62,  -116,   -67,   -72,   -44,   -23,    11,   -25,     9,   -15,     4,   -13,   -12,    60,   107,    97,    90,    52,   -50,   -88,  -137,     4,    68,   -66,   -89,   -14,    10,   -22,   -67,  -103,   -99,   -36,   -19,   -36,     0,   -57,    -2,     6,   -16,   -73,    31,   124,    57,   -21,    15,   -62,  -143,   -83,   -48,    28,     6,   -22,   -65,    12,    30,   -92,   -55,  -103,   -85,   -54,   -15,     1,   -54,   -40,   -10,   -16,    -9,   -82,   -30,   109,   -24,    35,    22,   -82,   -99,   -75,   -89,   -44,   -47,   -34,   -45,   -43,   -49,   -97,  -117,   -95,   -91,   -22,   -29,   -11,   -54,    -7,   -53,   -41,   -32,   -70,   -11,    88,    12,    11,    49,   -61,   -28,    13,   -70,   -63,   -54,   -89,   -74,   -51,  -110,  -141,  -134,  -111,   -37,   -25,    -8,     2,   -56,    -6,   -52,   -38,   -15,   -46,    21,   -12,    11,    19,    57,   -33,   -14,    10,   -85,   -75,   -40,   -98,   -19,   -68,   -91,   -71,  -113,   -94,   -45,   -23,   -38,   -13,   -54,   -11,     3,     5,     8,   -67,   -32,   -59,   -70,    22,     2,    39,    15,    -5,   -38,   -16,   -55,     3,    21,   -58,  -129,   -93,  -101,   -63,    -8,   -25,   -18,   -27,   -96,     0,     0,     5,   -25,   -23,   -76,   -28,    65,    97,    83,   121,    46,    24,    23,   -19,   -77,    13,   -50,   -65,   -67,   -52,   -28,    -1,    -3,     3,   -42,   -31,   -30,    -1,     3,     1,   -27,   -23,   -38,   -83,   -10,    57,    47,    14,   -22,     6,    37,   -30,    51,    12,   -26,   -46,   -28,     4,     5,     8,    12,    -6,     0,   -20,   -47,     6,     0,    -2,     6,   -79,   -18,   -65,   -85,   -80,    24,     8,    17,     1,    20,   -36,   -54,   -61,   -12,   -26,   -13,   -12,   -80,   -38,   -52,     8,     4,    19,    18,   -19,   -16,    -9,    -9,   -11,    -1,   -39,   -18,   -19,   -19,   -14,    -7,    -8,     5,   -33,    -2,   -14,    -9,   -13,   -22,     5,    11,    -4,   -13,    16,   -15,    13,    -9,     6),
		    39 => (  -10,    -7,     4,    -3,    12,   -14,    -4,   -12,     6,     0,   -12,    12,   -20,    -4,     7,   -17,   -20,   -12,   -12,   -16,    -8,    17,     4,   -17,    -1,   -10,    -6,     6,   -20,    16,   -16,   -19,   -11,     7,    -8,   -17,   -11,    10,   -18,    -7,   -74,   -66,    -3,   -37,   -41,   -33,   -61,   -31,    -4,   -22,   -13,    -9,   -14,     3,    17,   -10,    17,     4,    16,   -18,    13,    12,     2,   -11,   -26,   -57,   -48,   -48,   -21,    10,   -53,     3,    -4,   -12,     5,    10,   -20,   -31,   -50,     5,   -10,    13,     4,    -4,   -13,     3,     6,   -43,   -32,   -14,   -24,   -37,   -89,  -127,   -75,  -128,   -57,   -79,   -49,   -70,   -40,   -27,   -36,   -32,  -100,   -76,   -28,     5,   -45,   -25,    12,   -13,    20,    14,    -2,   -33,   -70,   -96,  -175,   -28,   -76,   -77,     0,   -24,   -52,   -97,  -119,  -148,   -72,   -77,   -24,   -39,   -46,   -15,   -20,    -5,   -20,  -124,   -16,     5,    14,    12,    14,   -18,    -1,   -13,   -60,   -65,  -108,    20,    66,     5,   -11,    47,   -71,  -118,   -60,   -97,  -183,   -80,   -69,  -102,   -22,   -38,   -15,   -43,   -29,     2,   -13,    11,    -7,   -68,   -80,  -153,    20,   -51,    60,    65,    91,    29,    11,   121,    11,   -82,  -130,   -90,  -168,   -65,  -160,   -65,    43,    17,   -91,   -21,   -10,   -18,    19,   -28,   -86,   -76,  -115,  -132,   -95,   -53,    12,    99,    40,    13,     4,    32,   -33,  -131,   -47,  -127,   -56,  -105,  -180,   -65,    30,    -5,   -56,   -41,   -45,   -24,   -45,   -34,   -84,   -78,   -87,   -66,   -83,   -51,   -15,   -40,   -18,   -65,    12,    42,    64,   -43,  -100,   -55,  -111,   -53,   -88,  -101,     9,    -5,   -36,   -53,   -17,     0,    -2,   -19,  -110,   -27,   -11,   -35,    28,    93,    41,   -55,   -83,    39,    14,    50,    37,   -29,   -52,   -29,   -60,  -112,   -65,  -124,   -71,   -74,  -103,   -93,   -26,   -17,     2,   -51,   -80,     4,   101,   -42,    65,     1,    40,   -63,   -16,   -16,   -38,   -24,   -54,    30,    13,   -33,   -16,  -102,   -76,   -27,  -186,  -199,  -104,   -73,    -3,   -57,    -5,  -113,   -45,    68,   -24,   -15,   134,    85,   -53,  -108,   -53,   -83,   -34,    31,    32,    65,    27,    74,   -54,    11,   -34,   -68,  -153,  -116,   -88,  -171,   -12,   -66,   -15,  -102,   -61,    41,   -18,    80,    92,   -47,   -52,   -22,   -70,  -134,   -45,   -25,    56,    46,   -21,    50,     8,   -40,   -10,    41,   -79,   -61,   -15,  -115,   -90,   -41,   -15,   -99,   -43,    -5,   -68,    95,    -1,   -15,     9,   -20,    38,   -94,   -50,   -25,    13,   -67,   -33,    -6,    41,   -13,    50,    38,   -13,   -86,     5,   -84,   -50,   -26,   -31,   -24,   -28,    96,     5,    34,    16,   -12,   -20,    73,    81,    90,    15,    34,   -46,  -136,   -78,    20,    77,   -14,   -42,    46,    22,   -16,    40,  -119,   -49,     6,   -14,    -8,   -28,    87,    44,    61,    56,   -70,    28,    26,   -15,    38,    83,   -82,   -27,   -98,  -145,   -39,    44,    28,    31,   -17,   -20,    -3,    32,  -124,   -76,   -51,   -12,   -19,   -70,    23,   112,   -79,    53,   -27,   -14,   -36,   -28,   -24,    16,   -38,  -113,  -135,   -93,    10,    99,    86,   -28,   -26,   -82,   -13,    53,    -2,   -62,  -110,    18,   -13,   -64,    14,    28,   -44,    14,   -59,     2,   -34,   -13,     5,    37,    42,   -47,   -60,   -24,    38,    -5,    82,   -26,   -42,  -138,   -41,   -47,   -93,   -82,   -94,   -15,     8,   -67,    24,   -49,    50,    47,    31,   -43,    -3,    42,    69,   -11,   -10,    64,    77,    55,   -58,    16,    43,    43,  -136,   -88,   -56,   -41,   -91,  -108,   -71,    11,    -9,   -56,    -6,   -50,   -33,    26,    59,   -10,    58,    45,    48,   113,    61,    13,    -4,    -2,  -114,   -80,    23,    23,   -42,   -40,    27,     7,  -124,   -76,   -33,   -19,   -35,   -29,   -15,    24,   -14,   -99,  -106,    27,   -62,     5,   -71,   -91,   -71,   -67,  -118,  -112,  -118,   -34,    98,    21,   -30,   -40,    30,   148,    11,  -131,     1,    14,   -11,   -67,   -16,    14,   -14,   -27,  -111,  -188,  -191,   -74,   -54,  -100,   -97,  -140,  -141,  -176,   -97,   -56,    72,    12,     2,   -47,    10,    87,   -66,  -165,    -4,   -20,     2,   -73,    46,   -20,   -31,   -36,   -52,  -117,  -150,   -45,    59,   -23,    49,   -19,   -95,   -43,   -91,    -7,    19,    42,   -15,    17,     6,    62,  -112,   -76,   -18,    11,   -18,    -5,    75,    23,    14,   -35,   -49,   -72,   -76,   -52,   -56,     7,    33,     8,   -20,   -70,   -49,   -24,   -43,    36,    14,   -22,   102,   122,   -88,   -60,    -4,    11,     7,   -59,    -6,   -18,     6,   -32,   -43,   -54,  -106,   -69,   -83,     3,    -1,     6,   -53,   -28,    -6,    40,    84,   150,    29,   113,   178,    37,    41,     3,   -19,     5,    -6,    60,   -34,   -43,    26,   -16,   -55,   -75,   -67,   -17,    20,    -5,    26,  -111,  -133,  -139,  -109,   -23,    89,    52,    37,   -10,   -67,   -54,     8,   -27,    12,     6,    20,    13,    40,    -5,     8,    44,    19,    24,     8,     0,   -47,   -32,    36,    35,   -36,   -99,   -82,  -101,   -87,     6,    11,    43,    92,    65,   -13,    -4,     8,     2,   -17,   -18,   -13,   -24,   -38,    19,    -6,    11,   -10,   -14,    -6,    34,    40,    43,    -4,   -51,   -56,    44,    29,   -50,  -105,    -7,   -55,    12,    12,    -2,   -13),
		    40 => (  -20,    -3,     2,   -17,   -14,     8,     6,    -7,   -19,    -5,    12,   -12,    18,    -5,   -10,    -3,     1,    13,   -14,     5,    -9,     1,     7,    18,    10,     7,    -6,    -1,   -11,     3,     8,    -3,     7,    10,    19,    -3,    -4,   -16,   -31,    14,    42,    -6,   -12,    29,    54,    58,    -2,     2,    18,     9,    -3,    18,   -20,   -12,    -8,     0,    -8,     3,    19,    52,    39,    -9,     4,    11,   -57,  -113,   -97,   -62,  -102,  -155,  -122,  -154,   -34,   -71,   -62,   -95,   -94,   -19,   -86,   -49,   -32,   -14,    -8,    10,     7,   -14,   -18,    32,     4,   -29,   -71,   -29,   -39,    -2,   -13,   -51,   -45,     0,    -1,   -24,   -42,   -78,  -140,  -163,   -36,   -44,   -96,   -77,   -56,   -21,   -69,     2,    18,    -2,   -13,   -33,    -8,  -117,  -101,   -49,   -35,    58,   -10,   -42,  -103,    -7,     0,   -30,    28,   -74,   -91,   -54,   -66,   -45,    39,   -93,   -52,   -58,   -92,     0,    -2,    11,   -43,    46,   -12,   -52,   -15,     6,    61,   -45,   -14,   -56,   -56,    34,   -15,   -57,   -22,    29,    -5,   -73,  -103,   -74,   -18,   -67,   -41,   -51,   -79,   -70,    14,     6,   -30,   -33,    68,    54,    19,    13,  -119,  -104,    -8,   -39,   -49,    44,   -36,   -65,    21,    31,   -69,    52,   -12,    67,    24,  -126,   -64,  -139,   -72,   -37,    14,    -4,   -31,   -43,    68,    67,    15,   -47,  -143,    17,   -24,   -56,    -1,   -33,   -10,     4,    27,    70,   116,   109,    26,    32,    19,    48,   -93,   -53,  -145,    50,   118,   -64,    80,     6,    48,    37,   -35,    10,    -9,    -3,   -31,   -36,   100,     0,    48,    31,    52,    63,    90,   -68,     6,    48,    24,    71,  -122,  -163,  -133,   -21,    -8,   -22,    89,    -6,  -113,   -10,   -22,   -44,    28,     8,   -61,   -56,     3,   -38,    44,    -6,   -72,    24,    49,   -28,   114,   -37,    -6,   -19,     9,  -172,  -148,     0,    -7,    -9,    88,    -1,   -72,   -90,     2,   -46,   -14,   -19,   -68,  -104,    14,     3,    65,    -3,   -22,    29,    -7,   -44,    93,    56,   102,   -21,     0,  -114,  -138,     2,   -17,   186,   -63,   -18,   -84,  -104,    69,    96,    27,    38,   -24,   -21,    21,   -24,    21,   -53,   -61,    22,   -77,   -31,    53,    88,    70,   -68,   -70,  -116,  -114,    -9,    14,    27,   -24,   -27,   -81,   -70,   113,    78,    39,    44,    -8,    23,    11,   -49,   -81,   -68,  -141,   -92,   -31,   -27,    41,    96,    28,    14,   -11,   -29,  -124,     8,     4,    37,    45,    60,   -35,    32,    79,    83,   134,    54,   -22,    22,  -103,   -88,   -37,  -164,  -115,  -134,    39,    10,    21,    68,    85,    63,    17,    67,   -67,   -22,    -5,    18,   -13,    25,    23,   123,    99,   175,   103,    41,     7,    23,   -38,   -15,   -87,  -104,  -159,   -73,   -22,    59,    38,     3,     7,    97,   -25,   -14,   -99,    14,    -7,     5,   -39,   -48,   -10,    80,     5,    70,   154,    65,   -12,   -11,   -43,   -62,  -101,  -108,   -48,  -113,   -22,     1,    56,    99,    74,   138,    98,    20,  -156,   -41,    -8,   -15,   -35,   -70,    66,    -9,    81,   117,    44,    30,    38,   -51,   -86,   -84,  -119,  -104,    -9,   -25,    29,   -73,   -37,    88,    57,    -1,    51,   -55,  -173,   109,   -12,   -14,   -50,  -120,    26,   -49,   -12,    13,    69,    87,    -6,   -93,  -153,  -105,   -35,    55,    -6,   -28,   -74,   -60,    28,   -74,   104,   -37,    31,   -86,  -127,   123,    18,    14,   -37,  -121,   -32,   -98,   -25,    68,   160,    93,    31,   -75,  -151,   -77,    53,    24,    -2,   -28,     1,   -12,    32,     6,    58,   -65,   -10,    -5,   -77,   -52,    10,    55,   -55,   -48,   -30,   -71,   -52,   -28,   141,    57,    33,  -115,   -52,   -70,   -57,   -28,    10,   -50,   -17,   -78,   102,   -20,    47,   -16,    -9,  -148,   -13,   -12,    -5,    43,   -95,     5,   -21,    17,   -31,   -20,    55,    88,   165,   -62,    -5,   -46,   -35,   -71,   -54,   -45,   -64,   -29,   -90,   -65,   -39,  -121,  -108,   -79,    42,    14,    -5,   -18,  -131,   -59,   -31,     0,   -59,   -67,    31,   -26,    -6,   -55,   -67,   -86,   -65,    -1,    35,   -45,  -124,   -88,   -67,   -42,    75,   -38,   -66,   -60,    64,    31,     6,   -17,  -124,   -30,  -115,   -23,    10,    13,    86,    71,    55,   -66,   -27,   -27,   -34,   -15,   -81,  -103,   -79,   -10,   -64,    15,    24,   -40,   -45,    13,    64,    42,    -1,    19,   -13,  -142,  -108,   -74,     7,     9,   -11,    34,    44,    57,   -40,     3,   -43,   -43,   -54,   -64,  -128,   -66,  -125,   -33,   -81,   -74,   -86,   -27,   -60,   -10,   -19,   -18,   -19,    12,    12,    54,   -68,   -80,   -16,    80,    57,    58,    62,   -52,   -18,    27,   -71,  -126,   -81,   -85,   -73,   -85,  -110,   -90,   -18,    34,    -1,   -10,   -15,    17,   -20,   -12,  -106,  -158,  -137,  -109,  -110,   -99,  -147,  -146,  -175,   -85,   -75,  -199,  -200,  -181,  -220,  -149,  -118,   -91,   -84,   -44,   -27,     9,    -5,     3,     6,    14,    -8,    -5,   -42,   -60,  -148,   -74,   -71,  -125,  -140,  -161,  -108,  -103,   -87,  -112,   -83,  -155,  -150,   -98,  -126,  -108,   -47,   -61,     3,    -7,     9,   -19,   -13,    -8,    -8,   -11,    16,   -15,   -19,    14,     4,    -7,     2,     7,   -16,   -67,   -29,   -39,   -38,   -32,   -16,     9,     5,   -63,   -41,   -37,    -6,     4,     9,     7),
		    41 => (   18,    -5,     4,    18,   -18,     0,   -13,    -4,   -20,     5,     7,     7,    -4,     5,    -1,    19,    -7,    17,   -11,   -10,   -16,    20,    16,    10,   -19,    -6,    -7,   -17,    -2,   -14,    -4,    -7,    17,   -13,   -11,   -17,    14,    -2,   -22,   -19,   -41,   -51,    18,    45,     3,   -38,   -12,    11,    12,     4,    12,   -11,    -9,   -18,   -16,     1,     0,   -18,    17,   -15,    -2,   -14,     7,    -2,   -30,   -38,   -56,   -40,   -45,   102,   130,   171,   149,    86,    88,   172,   124,  -109,  -119,   -81,    10,    15,     0,    14,    17,   -12,    64,   120,    -9,   -57,   -90,    76,    52,   -19,  -163,  -162,     8,    15,    24,    70,   149,    68,    65,    79,   125,   113,   -65,   -77,   -39,   -30,    18,    18,    20,     9,    13,    76,     5,    25,   -34,   -97,   -76,   -42,    20,   -44,  -108,  -125,    22,   110,   110,    46,    83,    27,    30,    71,   -65,   -53,   -31,   -88,   -80,   -65,   -20,    -3,    55,    47,    11,    95,    35,  -105,   -71,   -78,   -36,   -39,  -118,   -60,   -19,    62,   106,    27,    -3,   -41,   -43,    64,   -68,   -16,   -37,   -74,   -71,   -37,   -12,    -7,   -79,     8,     9,    27,   -75,   -93,   -50,   -57,   -85,   -84,   -33,    20,    19,    65,    92,   -22,   -22,   -57,   -19,   -47,   -46,     7,    12,    -1,   -56,   -44,   -14,   -26,  -106,   -28,   -52,  -132,  -146,   -20,    53,    46,   -46,    11,     8,   -45,    89,    21,    13,    25,  -172,   -97,   -19,   -64,   -86,   -32,    -7,    -6,   -70,   -73,   -17,   -36,  -102,     3,   -55,  -145,   -75,   -62,    27,   188,   -15,   -51,   -36,   -32,    36,    57,   -13,   -41,   -24,   -95,   -11,   -55,   -53,   -38,   -30,   -17,   -69,   -37,    -3,     1,  -116,   -26,   -52,   -80,    -6,    25,    88,    63,    27,   -65,   -66,   -29,    37,    63,    52,  -141,   -59,  -151,   -76,   -83,   -36,   -49,   -30,   -33,   -24,   -51,    20,    -3,  -123,   -16,   -83,  -129,   -71,    70,   -60,   -64,   -33,   -13,     1,   -54,     1,   -12,     1,    -1,   -67,   -66,   -71,   -82,   -30,   -17,   -19,   -34,   -49,    59,    -4,    25,    10,   -13,   -48,   -68,     4,   -41,  -117,    18,    79,    -9,    -5,   -93,     2,   -12,   -23,   -68,  -147,   -79,   -85,   -40,   -57,   -10,   -53,   -26,   -77,    14,    -9,    15,    -7,   -16,   -10,   -34,   -38,   -68,   -84,    62,     0,    73,   -52,  -149,   -10,     4,    21,  -117,   -59,  -120,   -71,   -22,   -39,   -11,    -9,   -17,    10,    14,    -7,    11,    15,    -1,   -64,   -35,   -32,   -68,   -27,    89,    20,   -12,   -37,  -257,    11,    42,     5,   -54,  -187,  -115,   -69,   -89,   -57,  -119,   -94,    -6,    -7,   -11,     2,    14,    -5,   -14,   -62,   -77,   -98,  -121,    84,    54,    19,   -96,  -259,  -132,    68,     7,   -43,  -119,  -177,  -139,  -122,   -97,   -94,   -83,   -19,   -34,    37,     7,   -15,    -1,    22,    22,   -92,  -107,  -131,   -99,    98,    61,   -72,  -153,  -196,    19,    26,   -15,    -5,  -147,  -189,  -161,  -128,   -71,   -71,  -106,   -72,   -31,   -13,   -49,    -7,    10,     6,   -43,   -68,  -101,   -75,   -53,   -43,   -35,  -234,  -181,  -269,   -21,   -60,   -78,  -120,  -187,  -237,  -155,  -106,   -79,   -60,  -144,    37,   -72,   -90,   -34,    11,     7,   -14,   -68,   -12,    32,   116,   -27,   -77,   -60,   -24,  -148,  -188,   -65,   -13,   -88,   -61,  -104,    13,    81,    33,     7,   -16,  -126,     8,  -169,   -45,   -54,   -10,    -4,   -15,   -17,   -46,   111,    -7,   -30,    42,   -35,   -10,  -164,  -192,   -47,     8,   -19,    34,    -2,    16,    55,    97,    11,   -33,   -32,     4,   -55,  -100,   -14,     7,   -14,    20,   -32,   -77,   -29,     6,     4,    42,    45,   -26,   -38,  -104,   -28,     0,    17,    96,    11,   -38,    56,    85,   -24,    10,    47,   -14,   -75,   -89,   -63,     2,    -8,    18,    86,    84,  -205,   -32,   -77,   -16,   168,    32,   -14,     3,    50,    63,    47,    96,    40,   110,    86,    60,    34,   141,    73,     6,   -40,   -33,    20,    60,    57,   -25,   132,   115,    60,   -23,    53,    58,    71,   108,   -64,   -29,    57,   -20,    -6,    21,   -24,    46,    15,    68,    87,     5,   -36,    29,    46,   -54,    -3,    41,    36,   -55,    75,    47,   173,   113,    16,    39,    40,     1,   -12,    13,    -7,   -96,    -3,    -7,   -14,   -13,    -1,    42,    68,    61,    85,    96,    87,    36,    -9,    16,    -4,     7,   -23,    -2,    51,   128,   -60,  -102,    36,     7,   -49,     3,   -14,    16,    28,    -3,   -28,  -112,  -276,  -228,  -168,   -42,   -80,   -84,   -80,    47,    12,    -2,   -20,     5,   -30,   -26,   -61,   -39,   -52,   -30,    40,    26,   -28,    17,    -4,    30,     4,   -97,  -128,   -80,  -143,   -82,    -3,   -67,   -66,  -119,   -29,    22,    11,     7,     9,    -2,    -5,     6,    -4,   -22,     4,    30,    35,   -15,     1,   -20,  -129,    14,    32,   -76,  -241,     0,   -35,   -72,   -89,   -77,   -53,    -4,     6,    14,    14,    18,     2,     6,    11,   -40,   -63,   -23,   -15,   -52,   -59,    -8,     1,  -132,  -129,    17,    55,    65,   -74,   -17,    10,     5,   -23,   -19,    14,    17,     0,    -5,   -10,     9,    12,    12,    15,     3,    -8,    -2,     0,    20,   -16,   -50,   -46,   -17,   -38,    13,   -38,   -60,    -7,   -11,    -1,    -3,    17,     9,    20,   -19,   -11,     0,    19),
		    42 => (  -18,   -16,    14,     9,   -13,   -10,     8,   -17,    18,     6,    -7,     7,   -20,   -26,    20,    31,     2,    12,    -3,   -19,    -8,     5,     0,    -8,   -17,    -3,    -6,   -11,    10,   -12,    -6,    18,    -6,   -10,     1,     0,    19,    -2,   -48,   -41,   -36,     7,   -45,   -50,    16,     5,   -19,  -134,   -45,   -38,   -31,     5,   -20,   -14,     1,     1,    19,    -4,   -13,   -49,   -30,    -4,    -6,   -24,   -15,    -4,    91,   103,     8,    27,    53,    55,    94,   110,    35,   -11,    -4,   -31,   -49,   -29,    11,    13,   -15,     3,   -16,    10,    -6,   -74,   -87,   -43,   -17,   -51,    46,    51,   120,     6,   -30,   -14,   -38,   -18,    21,   100,   -74,   -11,   -15,    55,    -6,   -51,   -22,   -34,    -6,    13,     0,   -18,   -37,   -63,     0,   -24,   -37,   -10,    86,   169,    74,    -6,    81,   -30,   -36,   -11,    57,    28,    30,   -24,   -95,   -64,   -22,   -70,   -82,   -55,  -131,   -69,   -14,    -1,   -23,    -4,   -20,     6,    24,    46,     7,    17,    54,   126,    41,    96,    91,    50,    93,   -26,   -25,    58,    35,    -3,   -83,   -76,   -69,   -23,  -173,   -64,    13,    10,    31,   -52,   -25,    57,    62,   109,    48,    27,    49,    29,   -16,   -40,    26,    61,    79,    33,    82,    -1,    37,    82,   -49,  -184,  -188,   -14,  -141,   -25,    14,    -5,    62,   -34,   -21,    44,    61,    83,    40,    15,   -41,   -27,    73,    57,    -9,    63,    60,    29,    -1,   -45,   -27,    21,   -88,  -108,    12,    82,  -214,   -90,   -51,    74,    78,   -26,   -10,    17,    35,    15,   -38,   -10,   -48,    32,   -41,   -42,   -33,   -75,    20,   -44,   -61,   -32,  -103,   -49,   -19,   117,    59,   -29,  -146,   -86,    11,   -89,    89,    26,     8,    11,    22,     3,     9,    47,    62,     5,   -51,   -63,   -81,   -33,   -35,   -17,  -105,   -82,   -36,    20,   -33,    73,   -15,  -115,   -51,   -35,   -20,   -37,   100,     1,    33,     9,    -6,   -11,   -49,   -11,    17,    30,   112,   -12,   -28,   -10,   -11,    30,   -74,   -64,   -52,   -41,   -97,   -88,   -41,   -67,   -32,   -70,    -1,   -49,   -30,   -62,    -3,    30,     7,   -26,   -20,   -81,     4,    26,    59,   -72,     0,    41,     5,   -32,  -107,   -18,    28,     1,   -55,    21,   -43,    53,   -87,  -111,    10,   -47,  -121,   -36,     3,   -12,    11,   -45,    52,   120,    66,    36,    77,   -69,    17,    12,   -25,   -17,    -2,    90,   -34,    55,   102,    71,   -12,   -10,    -4,     2,     1,   -24,   -61,   -74,   -16,    -4,    63,    61,    86,    39,    -1,   -39,    -3,    -8,     2,   -37,     9,    37,    84,   108,    69,    72,    75,    38,   -37,   -57,   103,     8,    -8,   -62,   -18,   -11,   -88,  -101,    20,   140,    99,    19,   -51,   -24,   -57,   -69,   -95,   -48,   -41,     2,   133,    99,    62,   107,   124,   148,   122,    25,    78,    78,    17,   -44,    75,    26,   -76,   -43,    -2,    32,   106,    44,   -60,    31,   -31,  -146,  -121,   -42,   -33,    20,    16,   107,   122,    92,    58,    94,    14,    16,     8,    69,     6,    -6,    84,   -56,   -78,   -81,   -29,    73,    51,    48,    28,    47,   -70,   -99,   -84,    75,    15,    40,   139,   143,   124,   161,    85,   193,    60,    77,   111,    55,    -4,    -7,    82,   -19,   -93,   -44,   -50,   -24,    73,   116,   106,    71,    43,   -27,     5,    42,   -61,    -3,   106,   174,    98,    35,    30,    28,   -33,   -62,    83,    61,    -5,    -3,    11,   -38,   -46,   -28,    -8,    11,    40,    91,   159,    72,   -11,   -30,   -61,   -28,    -7,    91,   153,   193,   147,    51,    26,    42,    47,   -86,   -39,    96,    12,   -29,   -59,    -9,   -24,    -6,   -17,    21,    42,   111,    85,    48,    38,  -109,    -9,    15,     8,   245,   265,   229,    90,    54,    70,    27,    24,   -91,    -5,    66,     0,   -42,    19,    29,    12,   -80,   -98,     8,    56,    17,    79,    62,    71,   -25,   -65,    38,   188,   169,   182,   124,    64,    -7,   -72,    11,   -23,   -19,   -47,     3,   -11,    -9,    61,     0,    96,   -30,  -100,     9,     1,   -46,   -39,     4,     2,    26,   -19,   130,   209,   188,   144,   147,    38,   -21,   -21,   -44,   -87,   -37,     8,     9,    -9,   -19,   -26,     9,   -43,     4,   -78,   -49,    -5,   -49,   -39,    -6,    85,   -14,   -23,   129,   276,   178,   235,    82,    53,   -20,   -20,   -35,     4,    64,    -4,   -11,     2,    14,   -13,   -11,   -46,    -6,   -39,     4,    54,   -53,  -156,  -102,    -5,    19,   105,   219,   298,   241,   187,    89,    -3,    58,   -69,    -7,    42,    47,   -70,    13,   -16,    13,   -52,   -71,  -216,  -214,   -64,   -47,   -13,  -144,  -116,   -74,   -58,    95,   138,   104,   214,   207,   151,    42,    -7,     2,   -49,   -29,    46,     3,    32,    15,    16,    17,    -7,   -38,   -84,  -140,    90,    28,   -24,   -56,    -2,   102,   162,   196,   216,   200,   142,    67,    73,    39,   -26,   -43,  -130,   -13,    18,    49,    33,     1,   -11,    20,    -8,     1,   -37,  -103,  -153,  -142,  -141,  -153,  -166,   -84,  -119,  -108,  -146,  -107,  -107,  -105,   -93,  -129,   -53,   -50,  -154,    -3,   -12,    -6,    15,    13,   -14,     0,    11,    18,   -29,   -17,   -14,   -24,   -27,   -16,   -30,   -33,   -13,   -34,   -39,   -14,   -23,   -25,   -34,   -11,   -85,  -122,   -20,   -26,   -20,    11,   -16,   -11),
		    43 => (  -15,   -11,   -14,     4,    -7,    -8,    -4,    16,    18,     9,    -5,     6,    -2,     1,   -26,    -4,    10,    -2,   -15,     6,     9,     4,    12,    12,   -10,    -1,   -14,    -2,     7,    -4,    -7,    -2,   -19,   -13,     5,     5,   -17,   -12,   -36,   -44,   -32,   -71,   -56,  -127,  -173,  -191,   -71,   -20,    -3,   -16,     1,   -13,    18,    -4,    -3,     5,    -9,    11,    -1,   -15,   -31,     9,   -41,   -69,  -130,  -130,   -28,     1,   -15,   -13,     0,    -4,    32,   -12,   -69,   -54,   -78,   -92,   -95,  -119,   -42,     2,     1,    -1,     1,    -1,    -2,   -49,   -28,    24,    -8,    33,    79,   -28,    -1,    32,   114,   -15,    -7,   117,   129,    93,    40,   -71,    11,   -56,   -93,  -211,  -174,   -70,    15,    -1,     4,    90,  -139,    33,    40,   -44,   -94,  -104,    34,    67,    99,   -26,     5,    -1,   -15,    18,    68,   -36,   -53,   -93,   -78,   -20,   104,  -101,  -208,  -189,   -48,    -3,    -3,     7,   -36,    27,   -39,    -7,    29,    39,   -16,    11,   -14,    10,   -12,    41,    14,    37,    58,   -33,  -121,   -14,    55,   -37,   -57,   104,   -25,  -219,   -78,   -10,   -11,    20,   -87,   -38,   -88,     9,    81,    61,    14,    17,   -20,   -92,   -98,     3,    47,    74,    54,   106,    64,    49,    43,    86,    32,    37,   132,  -199,  -167,   -79,     7,   -11,   -20,    15,    14,     3,    10,    30,    -3,   -11,   -57,   -31,   -16,    27,    38,     9,   -42,    66,    75,    27,   -38,    25,   -25,   165,    74,  -269,  -156,   -90,   -62,   -23,    42,    66,    19,    -2,   -40,    20,   -16,   -40,    36,   -15,    78,    71,   -55,   -90,   -22,    29,    47,   101,    14,   -72,    76,    73,    12,  -296,  -192,   -11,    -1,  -111,    -1,   -34,    56,   -12,   -78,  -107,   -97,    -5,  -106,   -16,   183,   128,    49,    22,    63,    22,   -15,    26,    79,    -7,   120,    86,  -151,  -234,  -204,   -80,     9,  -111,    24,    41,   -56,   -66,  -125,  -132,  -150,  -156,  -181,   -41,   110,   166,   208,    67,   -56,   -34,   -63,   -45,     7,    44,    15,    39,  -150,   -96,  -152,   -82,    -9,   -61,   -19,    86,    12,   -72,  -179,  -164,   -73,  -121,  -229,   -49,    30,   168,   104,    92,    34,    12,   -11,   -60,   -35,   -58,   -80,  -151,  -384,  -194,  -124,   -19,     6,   -30,    11,     8,   -30,    -3,   -73,  -132,   -45,  -211,   -43,   -89,    39,    94,   238,   118,   -23,    47,    51,   -56,    -2,   -36,  -230,  -268,  -282,  -140,  -102,   -19,    -1,   -17,  -237,   -51,   -64,   -72,   -32,   -67,   -20,   -85,  -102,   -54,    17,    75,   164,    61,   148,    33,    42,    36,    18,   -69,  -158,   -67,  -166,  -167,  -112,   -19,   -24,    60,     8,  -137,  -148,   -98,   -63,   -79,   -66,   -29,  -115,   -33,    -4,    83,    65,    99,    39,    -2,   -88,   -71,   -78,  -109,   -55,    14,  -132,  -152,   -86,   -25,    -6,    33,    -1,   -89,   -22,   -22,    27,   -14,    28,  -134,  -129,    33,   125,   126,    97,   123,   -33,  -129,  -147,   -67,   -42,   -17,    72,    72,    57,  -115,    21,   -59,     2,    12,    37,    70,    13,   -40,     0,    10,     0,   -60,   -21,    68,    46,    24,    97,   -38,  -154,   -87,   -42,   -21,   -75,   -69,    91,    17,    58,  -213,  -140,   -67,     3,    27,    50,    60,    39,   -79,   -33,   -32,  -102,   -69,   -14,    95,    13,    51,    -8,  -103,  -132,   -77,   -76,   -25,  -105,   -26,    10,    11,     7,  -166,   -37,   -57,   -42,    16,    65,    90,    -1,   -24,    27,    66,   -53,   -30,    73,   120,     0,     5,   -49,   -60,   -38,     9,   -51,    16,    31,    54,   -45,   -49,   -88,  -144,   -30,   -80,    -3,   -61,    51,   149,    70,   105,   -55,    68,    -4,    37,    95,    27,   -85,   -57,  -116,    23,    19,    51,    51,     9,    34,    31,   -71,   -37,   -54,  -115,  -143,   -80,     4,   -60,  -102,    33,    -5,   -73,   -75,    43,    64,    19,    63,    30,  -105,   -33,   -35,    63,    70,    29,    -9,   -25,   -16,    32,   -45,    -7,   -73,   -94,   -23,    -2,   -14,   -23,   -63,    31,     7,  -114,     3,    77,    79,   -27,   -60,   -58,   -50,    15,   -26,     8,   -19,     5,    -8,     7,   -53,   -45,    -4,   -74,  -179,  -116,   -48,   -14,     4,     1,   -30,    40,   -77,   -48,    84,     6,   -71,   -39,   -27,   -31,   -12,    10,     0,    -6,   -20,    24,   -34,   -35,   -21,    16,    -3,  -129,  -157,  -211,   -18,    -4,     1,     6,    41,   121,   -29,    10,   102,    32,    63,    19,    90,    49,   -59,    52,   -71,    -2,    66,    -6,    61,   -20,   -49,   -72,   -83,  -106,   107,    20,   -66,    15,     8,   -14,    47,   121,   -24,    -3,    34,    11,   -52,   -66,    10,   168,   -92,   -10,   116,   -30,   -27,   -56,     4,     7,   -11,   -19,   -53,   -54,  -112,   -99,   -41,    17,    14,    -2,    16,   -62,   -74,   -61,   -95,    27,    43,     6,   141,   134,   209,    63,    -9,   -67,    56,     3,    25,    74,   -84,  -173,  -202,  -226,  -104,   -21,   -36,     8,    -8,    19,     5,   -63,  -141,   -67,   -76,   -35,   -15,   -40,    64,    39,    77,    18,  -121,   -70,   -11,    18,    34,   -63,   -55,  -119,  -161,  -106,    -5,     3,   -18,   -11,   -18,    -8,    10,    19,   -35,   -55,   -44,   -36,   -36,  -111,  -118,  -131,  -103,  -193,   -81,   -87,   -57,   -30,   -32,  -116,  -130,   -58,    -7,    19,    -8,     5,    -7,   -12),
		    44 => (   11,    13,    19,    16,   -18,   -11,    16,    20,    12,    19,     8,     6,     1,    -2,   -16,   -13,     2,     1,    -8,    17,    -1,     7,   -10,   -10,    18,    19,     7,    17,    -5,     9,    16,   -17,    -2,   -19,   -20,   -30,    -2,   -16,   -96,   -37,  -134,  -105,   -10,   -64,   -49,    -5,   -16,   -11,   -60,    -9,   -22,   -38,   -18,   -13,    -2,    15,   -12,   -19,   -18,  -101,  -108,  -121,   -50,   -89,   -73,   -67,   -28,  -123,    30,    12,   -62,  -147,   -94,   -77,   -78,   -29,   -34,   -44,   -63,   -13,    -9,   -16,    15,   -14,   -18,   -19,    -2,  -130,  -200,  -109,  -115,  -107,  -129,   -79,    62,   -48,  -121,  -246,  -148,   -16,   -34,   -12,  -103,  -110,   -23,   -33,   -81,   -43,     2,   -45,    -5,    18,   -19,    11,   -21,   -82,   -40,    28,    34,     7,   -23,    -3,  -107,  -182,   -19,    28,  -162,  -209,  -228,  -204,  -111,   -36,   -16,     4,    37,    62,    89,    26,   -57,   -30,    -3,    13,   -24,   -18,   -21,     3,   -38,   -33,  -111,  -177,  -141,    10,   113,   -40,   -80,   -30,   -95,  -383,  -203,    22,    90,    33,     9,     6,     5,    -5,   -52,   -35,   -16,    -5,    -3,   -75,    58,   196,   -26,  -125,   -73,   -56,   -93,    32,    88,    28,   -67,   -72,  -277,  -299,  -123,    90,    62,    26,     2,    63,    83,  -186,    59,  -160,    -4,  -137,   -14,   -64,    25,   166,   -85,   -48,   -37,   -16,    29,    53,    -6,    56,   -25,  -148,  -325,  -305,   -19,   102,    48,   -32,     7,    45,   -35,   -48,    63,  -168,   -56,  -118,    27,   -39,    -1,    39,   -62,    34,   -68,    -1,   -55,   -12,    58,    46,    17,  -154,  -394,  -119,    52,    51,    27,   -29,    76,   -76,     4,   108,    47,  -106,    10,  -100,    12,   -55,   -23,    29,   -54,   -38,   -44,    17,    -9,    11,    95,   100,    67,  -197,  -202,    54,   100,    36,    50,    29,    43,    33,   107,  -101,   -97,   -66,    15,   -65,   -93,    27,    58,    98,     5,   -52,   -10,    31,   -35,   -30,   -14,   129,   -48,  -217,  -146,    32,   101,    84,    11,   -16,    40,    67,    32,  -183,   -59,   -13,   -19,   -41,   -51,  -126,   -55,    41,   100,   -19,    46,   -41,    25,    -9,    96,   -45,  -147,  -216,  -128,   -49,    17,    19,   -93,    69,     2,   -21,    71,   -90,   -89,   -71,   -12,    -3,   -94,  -118,  -165,   -51,    25,    80,    65,   -63,   -24,    65,    86,    50,  -181,  -101,   -25,   -19,   -30,    64,     0,    91,    22,    70,  -110,   -95,  -186,  -107,    11,   -29,  -106,  -117,  -138,   -76,   -21,   -22,    41,    41,    67,    91,    22,    29,     8,    26,    31,    63,   -51,    64,    56,    36,   -12,   -42,  -187,  -154,  -147,    -2,   -13,   -18,   -24,  -125,   -97,   -10,   -14,     3,   -21,    55,    15,    61,    13,   -27,    63,    16,    -7,     6,   -31,    57,    24,   -42,   -51,   -27,   -90,  -104,  -119,     0,    -4,    -4,   -15,    37,    -5,     0,     3,   -20,    51,    18,    58,    46,    -1,    23,    42,     7,   -32,   -17,     4,   105,  -195,   -58,   -33,   -22,   -93,  -142,  -100,    -4,    -7,   -16,   -49,    32,    -3,   -32,  -133,   -11,    14,    10,     3,    -4,   -20,     1,   -53,     9,   -23,   -38,   -33,   -43,  -142,   -78,   -46,   -77,  -113,  -157,  -155,   -32,    -8,     3,   -64,    30,    84,   -13,   -96,   -45,   -63,   -32,   -31,   -28,    -4,     2,   -26,     9,   -53,    27,   -23,  -102,  -158,    27,   -30,   -32,  -119,    11,   -27,   -41,   -72,    14,   -83,   135,   178,   -78,   -50,   -99,   -75,   -90,  -178,    -5,   -65,    10,    19,   -15,    20,   -83,    -2,   -38,    13,    74,    35,    36,    -1,    68,    -8,   -18,    -6,   -88,   -41,   112,    57,   -83,  -109,   -67,   -36,   -97,  -104,   -24,   -85,     9,   -18,   -50,   -10,    16,   -35,   -39,   -25,    32,    21,    33,    73,    45,   -20,   -37,    19,     4,   -30,  -138,  -125,  -149,  -131,   -79,  -102,     0,   -56,   -59,   -79,    -3,   -26,   -46,    23,   -14,   -48,   -50,  -132,  -115,   -77,   -41,  -123,  -181,   -33,     9,     9,     2,   -33,   -82,  -135,   161,   -13,    26,   103,   130,   -36,   -15,     8,   -13,   -40,   -28,   -19,  -136,  -116,    15,    16,   -17,    17,    50,   -68,  -240,   -81,   -20,   -16,    20,     8,   -90,  -153,    89,   100,    64,    57,     3,    63,     5,    -1,    -6,   -52,   -28,     7,   -58,  -105,   -46,     0,    17,    -7,    65,   -78,   -73,    36,    17,    14,     8,    -3,   -85,  -130,  -253,    41,    62,    51,    45,    32,    -6,    40,   -24,    26,    29,    79,   -55,   -51,   -29,   -19,    41,    18,    42,   -49,    14,    47,    15,     9,    10,   -10,   -29,  -197,  -166,   -28,   -83,     2,    28,    46,   -27,    17,    -1,    -8,    74,    34,   -90,  -213,   -50,   -38,    57,    30,    58,   -79,    84,   -61,   -17,    18,   -18,   -33,   -12,    -3,  -119,  -104,     2,   -15,   -64,     4,    16,    33,    56,     5,   -75,   -83,  -180,  -109,   -78,   -19,   -34,    50,   114,   -23,   -52,   -11,     2,     7,   -11,    -5,  -100,    10,  -110,  -104,  -174,   -86,  -108,  -113,   -79,  -147,  -207,  -236,  -317,   -66,   -87,  -133,   -64,   -80,   -84,   -62,    45,     3,   -17,    -8,    -9,    -3,    -7,     0,    10,    16,    -1,   -56,   -80,   -70,   -52,  -111,  -131,   -17,   -72,  -113,    -8,   -90,  -120,   -64,   -57,     8,   -18,    12,    -1,    -9,    20,    12,     8),
		    45 => (   -3,   -17,    -7,     0,   -14,   -18,    -3,   -18,    18,   -18,     8,    14,    11,   -10,   -20,     7,   -19,   -14,    13,    11,     2,   -12,    -8,    -1,    -9,    -8,    16,   -12,     0,    -1,     8,     0,    -3,   -13,   -14,    -3,    13,     4,   -16,   -37,   -34,   -36,   -52,   -79,   -90,   -69,  -100,   -97,   -96,   -77,   -11,     3,     7,    -4,   -19,    18,   -11,   -10,   -35,   -39,   -43,   -11,   -20,   -17,  -105,   -25,   -55,   -38,   -75,   -98,  -103,   -94,   -27,   -53,   -63,   -67,   -54,   -82,   -78,    48,  -135,   -19,    -6,   -17,    19,    -3,   -19,    85,   185,   -32,   -78,   -89,   -28,    40,   -29,  -123,  -101,  -163,  -135,   -66,    46,     8,    13,   -13,     7,    33,  -130,  -107,     3,   156,   140,     8,     7,    16,   -56,   149,    -7,    -7,   -88,   -77,   -70,   -18,    -9,  -145,  -158,  -110,   -82,   -57,  -107,   -97,    -7,    99,    -9,     1,   -95,     7,   123,   103,    10,   -44,    13,     2,  -103,   162,   -40,   -34,   -51,   -98,   -86,   -44,     7,     3,  -128,   -52,   -43,   -28,   -59,   -21,   -18,    68,    16,   -20,   -50,   -32,   -48,    36,    -7,   -41,    -9,    -3,   -80,   -28,   -52,   -38,   -59,  -104,   -53,   -13,   -19,   -90,    -8,    12,   -22,     5,   -13,   -75,    -6,   -39,   -44,   -80,   127,    96,    62,   128,   140,     7,     5,   -22,    16,   -43,   -32,   -76,   -58,   -73,    14,   -30,    -5,   -11,    46,    57,    59,    30,    68,    87,   -17,   -67,    -4,    49,    43,    52,    35,    -9,   164,    38,   -50,   -15,   -84,   -25,   -44,   -67,   -41,   -33,   -30,     3,     6,   -22,   -26,     6,    53,   -15,   -24,    19,    16,   147,   168,    79,   117,    94,    33,   -24,    58,    79,    19,   -36,  -163,  -116,   -54,   -57,   -81,   -44,   -26,   -50,   -56,    -8,    39,    -2,    34,     1,   -11,    26,   -39,   -89,    53,    21,    48,    81,   211,   166,    35,    39,     2,   -14,   -73,   -84,   -89,    46,   -42,    -4,    16,   -52,   -62,    -6,    67,   -11,    -7,    28,    68,   -93,  -326,  -347,  -189,  -165,  -176,   -60,    -3,    42,    20,    65,    -1,    12,     1,    69,    35,    42,   -33,   -38,   -74,  -141,   -29,   -91,  -105,   -69,     6,   -17,    17,   -22,  -172,  -202,  -300,  -276,  -278,  -219,  -177,   -38,    -6,   -40,    11,     1,    -6,    89,    41,   -18,  -104,  -139,  -120,   -90,   -27,   -89,  -121,    -6,    56,   -25,   -43,    33,     3,   -33,  -129,  -230,  -204,  -362,  -234,  -115,   -19,   -67,    -9,   -18,     1,   112,   -14,   -51,   -31,   -49,   -69,    -6,   -39,    -2,    80,    18,    34,    36,   -18,    24,    53,   104,    62,    69,    -8,  -133,  -189,   -55,    10,   -75,    23,     1,   -28,    67,   -81,  -116,   -12,   -78,   -96,   -23,    -4,    45,   -18,    10,    16,    72,    60,   -64,     0,    36,    94,   -27,     0,    86,    43,   -56,   -34,   -65,    19,    -8,   -72,    12,   -64,    -1,    46,   -17,   -40,  -108,   -32,   -48,   -46,    56,     7,   -80,   -47,   -10,   -43,   -30,    97,   -10,   -26,    73,   127,    -3,   -10,   -13,   -16,   -54,  -149,     7,    20,  -101,   104,    24,    11,  -153,  -128,  -140,   -86,   -28,   -13,   -55,    48,    34,    -3,    -4,   115,    84,     3,   -60,    15,    51,   -29,   -32,   -16,   -62,  -181,   -62,    78,   -22,    89,   171,    69,    10,    14,   -95,  -177,   -79,   -93,   -79,     2,    -1,   -14,   -52,    67,    -1,  -144,  -110,   -24,   -23,   -58,   -36,   -14,    -8,  -141,   -12,    19,    31,    51,   133,    78,    15,    30,   -45,    -5,   -52,    -3,    -4,   -12,    10,   -51,   -66,   -50,   -33,   -75,  -147,   -94,   -43,  -113,  -100,    11,   -28,   116,  -128,   -45,   -24,    58,   108,    75,   112,    51,    84,    81,    61,    28,   -11,   -30,   -50,    29,    47,   -34,   -59,   -70,  -100,   -61,   -47,   -64,   -76,    16,   -22,    96,  -166,  -114,   -10,    -3,   -71,    27,    42,    58,    42,    41,    -9,    16,     0,   -17,   -10,    -8,   -40,   -30,   -61,   -31,   -33,   -33,   -30,   -19,   -15,   -14,     6,   -55,     3,   -73,    46,   -41,   -12,  -105,   -71,   -50,    41,   -44,   -23,    32,     0,    29,    26,    24,   -45,   -76,    -3,   -13,   -26,   -30,   -29,   -18,   -15,    -9,    -9,  -160,    49,    63,    -7,   -83,     6,  -103,   -50,   -40,   -17,    -1,   -31,    22,    17,     3,     2,    -5,   -65,    -4,    46,    17,   -11,   -24,   -18,   -11,    13,     9,   -14,    19,    28,    95,   122,    14,   -65,   -85,   -78,    -8,   -11,   -74,   -98,   -12,   -44,    -2,    55,    68,     6,    -3,    46,    29,    -7,   -70,   -33,   -23,   -19,   -12,     6,   -76,     0,   -24,   -28,   -91,  -168,  -146,   -57,  -168,  -202,   -71,   -20,   -56,   -82,  -107,   -68,    12,    60,    49,    -5,    40,     9,    25,   -96,   -37,    -6,     9,    18,     2,    35,   -66,   -43,     5,   -39,  -105,   -27,  -184,  -175,    14,   -47,   -54,   -24,    -5,   -28,   -15,   -17,   -22,   -66,    27,     5,    19,    11,   -20,   -13,    15,    16,    18,   -22,   -34,   -43,   -68,   -38,   -52,   -43,   -29,   -43,   -33,    67,   145,   135,   112,    56,    -9,    81,     6,   -36,     3,   -16,   -15,    15,    12,    -2,    -5,   -17,    15,    15,    -6,   -26,   -11,     4,   -11,     3,    12,    -4,    -6,     3,   -14,    -2,     0,     5,   -38,   -37,   -32,   -33,  -104,   -19,    -2,    -3,    13,   -15),
		    46 => (  -11,     9,   -16,    -6,   -20,   -12,    -1,   -11,   -20,     0,    17,    -5,     6,    10,   -18,    14,     3,     4,   -13,    18,    -7,   -16,   -15,   -17,    15,     1,    13,    10,   -10,    10,    -3,   -11,    -4,    -3,    53,    76,   105,   113,    56,    38,    14,    36,    35,    13,     3,   -11,    24,    27,   137,    43,    24,    39,    -8,     6,   -10,     3,     1,    -8,    18,    13,    23,     7,    82,   114,   117,    58,   -36,   -33,   -34,    -3,   -15,   -12,   -21,   -51,   -17,    70,    63,    21,    24,    70,    64,    20,   -15,    -1,     8,    -9,   -92,   -62,     5,    15,    51,    85,    34,    62,     6,   -83,   -97,   -32,   -13,   -13,    -8,   -19,   -19,    28,     4,    63,    -5,    74,    90,    -3,   -37,    -7,    -4,   -19,   -48,   -22,     8,    23,    21,    12,    17,    21,   -60,   -53,    -1,   -51,   -26,    53,    40,     1,   -20,     1,   -14,    37,    -3,    32,    23,     8,    44,    58,   -15,    12,    14,   -34,    19,   -37,   -14,    19,    16,   -46,   -81,    13,    -7,   -46,    31,   -33,   -63,    18,    18,    14,    34,     0,    14,    43,    45,    12,    98,    62,     8,     0,     4,   -10,   -20,   -10,   -37,    16,     3,   -35,    16,   -15,    13,   -54,   -58,   -81,  -101,   -11,    22,    37,    51,    77,    52,    36,     2,   -59,    31,    40,    -9,    -2,    15,   -30,    -7,   -23,   -50,   -56,    26,    14,     6,   -26,   -91,   -43,    34,     5,   -46,   -26,   -53,   -12,    -5,   -17,   -25,   -20,    40,   -34,    14,    25,    11,    13,   -10,   -66,   -22,     0,   -30,   -66,    26,    25,   -12,   -89,   -58,   -20,   -22,   -60,    29,    44,   -45,   -47,   -81,   -30,  -119,  -100,   -70,   -75,   -26,   -82,     6,    14,   -11,   -20,   -37,   -77,     4,     0,    56,     9,   -35,   -62,   -64,   -66,   -21,    30,     5,   -18,   -59,  -106,  -113,   -91,  -146,  -106,   -36,   -56,    12,   -21,    -4,    -5,     1,   -38,   -17,   -57,     1,   -28,    47,   -64,   -61,   -98,   -46,   -67,    -8,    37,    -9,   -85,   -96,   -51,   -91,   -69,   -97,  -102,   -37,   -35,   -29,   -48,    -1,     2,   -12,   -14,    -6,    24,    58,    -5,    12,   -53,  -105,   -64,   -25,     0,    45,    -7,   -96,  -107,   -83,     1,    11,     0,   -22,   -29,    15,   -59,   -40,    -3,    13,    -9,    -3,    -9,   -55,    33,    13,   -30,   -16,   -43,   -96,   -40,   -37,    26,   -23,   -61,   -60,    45,    32,   -10,    22,    41,    31,    24,    29,   -77,   -91,   -18,   -13,     8,   -24,   -16,   -32,    52,   -19,    17,    46,   -74,   -91,   -52,    24,    25,   -71,   -26,     2,    -7,    29,    36,   -17,   -18,     1,    40,    58,   -57,   -54,     9,   -17,   -16,    12,   -10,   -24,    80,   -23,    21,    19,   -63,   -65,    66,    39,   -21,   -64,    -6,    15,    72,    70,    64,    -6,   -62,   -17,    44,    50,   -20,   -37,   -45,     4,    18,   -28,   -23,   -13,    46,   -15,    -3,    -3,   -26,   -70,   -18,   -37,   -83,   -32,    32,    64,    52,    64,    81,   -15,   -33,   -26,    58,    66,   -39,   -47,   -87,   -19,    13,   -19,   -39,   -10,    25,   -21,   -70,    19,   -41,   -40,   -29,   -73,   -19,    21,    15,    30,    66,     6,   -49,    -9,   -22,    -6,     5,    -2,   -21,   -40,   -74,    -4,    10,   -38,    -6,    -5,   -59,    -1,   -81,    23,    -7,   -25,  -114,  -100,   -11,    38,     9,    -9,     7,   -13,   -37,    51,    39,   -11,   -19,    -2,     7,   -28,   -81,    -3,    -9,   -36,    -4,   -21,   -54,   -85,   -43,    44,    33,   -22,   -60,   -32,    29,     0,    21,    -7,   -44,   -32,   -34,    57,    -6,     1,   -52,   -38,    -2,   -85,   -62,    -6,   -17,     4,     1,    -9,   -57,    -7,   -16,   -17,     8,   -48,    23,    -4,   -33,    19,   -49,    -5,   -40,    -7,   -33,    38,   -17,   -19,   -14,   -20,   -33,   -34,     1,    11,    -4,     8,   -44,    16,   -30,   -38,   -18,    -5,   -40,    38,   -10,   -61,   -43,    14,   -21,   -72,   -29,   -15,    13,    51,    28,   -39,   -60,   -20,    24,   -30,    -6,   -18,    19,    -6,   -27,     4,   -41,   -48,    13,   -19,    28,   -15,    -3,   -54,   -67,   -26,   -41,   -26,   -37,    -8,    19,    37,   -28,   -74,   -34,   -50,    12,   -16,     3,     0,    -8,     9,   -11,    -1,    -7,    29,    -7,     4,   -26,    -3,   -42,   -18,   -34,   -54,    -3,     8,   -16,   -59,   -34,   -49,   -25,   -82,   -47,   -31,   -40,    22,   -11,   -13,     7,    -4,   -30,    11,    -2,   -36,   -30,    26,    27,    15,    28,    53,   -49,   -27,   -47,    35,   -18,   -56,   -85,   -50,   -75,   -31,   -21,   -39,     7,   -29,    12,   -15,    -4,   -18,     4,   -25,     1,   -29,   -47,   -36,   -46,   -36,    -5,    -5,   -41,   -36,   -56,     3,     8,   -14,   -82,   -85,   -17,   -18,   -21,    -7,   -16,   -10,    18,     3,     4,    -1,   -17,    12,    -8,   -38,   -24,   -18,     7,     6,    -3,    -1,    -4,     1,    -5,   -20,   -27,     2,    -3,   -57,   -15,   -27,   -63,   -15,   -14,    11,     4,   -11,    14,    -9,    -5,    -4,   -17,   -13,   -22,     1,     7,     6,     0,    14,   -19,     8,     2,   -16,   -10,   -12,    -7,   -15,   -44,    -9,     6,    15,    12,    13,     8,    18,    14,     6,    14,     1,     8,     8,     4,     4,    -9,     4,   -20,    11,     9,   -17,   -15,    -4,    12,    13,    13,    -7,   -18,     2,     3,   -20,     7,    11,    12),
		    47 => (   -5,    -5,    10,   -19,    11,     4,   -12,    16,     5,     2,     1,    14,    -8,     8,   -18,    -3,     7,     3,     0,   -19,    -5,   -15,   -11,    13,   -11,    -4,    19,   -11,   -17,    -1,     4,   -15,    15,    18,    18,     1,   -17,    16,   -14,  -107,   -75,   -91,   -26,   -18,   -42,   -32,    11,    10,    17,     7,    12,   -16,    -2,   -15,     5,    -8,    14,   -20,    -5,   -11,    -6,   -19,    -8,    -4,     5,   -15,   -23,   -77,  -112,   -74,   -58,   -47,   -21,    10,     1,   -20,   -23,     3,   -25,    -6,   -19,     0,   -18,    16,     2,    -4,    19,   -38,   -41,   -19,   -30,   -66,   -54,   -37,     2,   -29,   -58,   -30,     6,   -85,   -86,   -53,   -37,   -14,   -33,    -6,   -72,   -18,   -24,    10,   -11,   -14,    13,   -13,    20,   -17,   -11,   -64,   -72,   -67,   -95,   -44,   -61,   -96,  -111,   -88,   -57,   -73,   -66,   -77,   -46,    -9,   -43,   -30,  -103,   -59,   -40,   -36,   -21,    -3,   -11,    14,   -11,   -54,   -40,  -102,  -129,   -82,   -22,   -26,   -98,   -16,    25,    -2,   -72,  -162,  -174,  -115,  -160,  -201,  -182,  -116,  -104,  -101,   -83,   -30,    -4,    18,   -15,     1,    13,    23,   -51,  -114,  -145,  -181,  -153,  -229,  -192,   -52,    67,    72,    24,   -59,  -113,    35,    55,     4,    38,   150,    40,    81,   -91,   -33,   -92,   -24,   -17,    84,    53,    79,    38,   -28,    79,    -6,   -74,  -198,  -179,  -170,  -130,   -34,   -22,  -102,    -3,     0,    41,   -63,  -125,   -62,   -51,   -30,   -24,    14,   -50,   -39,   -51,    97,   -41,    -6,   -15,     5,    82,    84,   -63,  -155,  -154,  -151,   -76,  -123,  -133,  -146,   -94,   -67,    28,   -69,   -80,  -128,   -48,    74,    38,     3,  -146,   -51,   -37,    87,   -48,   -42,    -3,    26,   133,   -12,    21,   -47,  -117,   -47,   -70,  -122,   -15,   -23,   -13,     7,    15,   -67,   -54,   113,    75,   155,    97,    31,   -97,     9,   -22,    50,    20,   -23,  -119,   -40,    55,     5,   -70,   -37,    -2,   -10,     9,    59,    25,     1,   -30,    83,    53,    50,   -12,    76,    68,    -9,   -69,   -22,  -109,    31,    -9,    25,    16,     8,    -2,    20,   -35,    94,   -30,     0,   -11,   134,    93,    64,    68,     0,   -54,   -46,    10,    45,    27,    44,    28,    47,   -27,   -59,   -21,   125,    -1,    -4,    35,    83,    67,    69,   -69,    74,    89,     2,    20,    88,   121,    25,   -64,   -67,    56,    88,    20,   -27,    -6,   -30,    64,    -9,   108,    80,   149,   150,     9,    28,    69,    89,    68,    29,    30,   -96,   -30,    12,    61,    21,     5,   -64,   -72,   -72,    42,   -23,   -20,   -12,    89,    51,    70,  -112,   108,   103,    59,   -26,   -29,    73,   125,    93,    25,   158,    10,  -107,    42,    52,    79,   -21,  -154,  -206,   -58,   -59,   -32,   -58,    75,    23,    50,    47,    33,    16,     8,   -36,   -89,   -17,    14,   -17,     4,   130,   -89,    43,   -21,    62,    -1,    84,    79,   -81,  -252,  -216,  -118,   -18,   -10,    39,    -1,    91,    73,   -10,   -25,  -123,  -105,   -26,    -7,    -2,    10,   -21,   -11,    62,   148,    11,    23,    33,    -8,    -4,   -75,  -308,  -355,   -71,   -40,    -2,   -15,     7,   -81,    27,    75,    53,    22,   -78,  -135,  -170,     9,   -73,    15,    -5,    77,    -5,    89,    -7,   -23,   -23,    -4,   -84,  -205,  -253,  -205,    -8,   -37,    19,   -65,   -23,   -44,   -63,    86,    59,    26,   -65,  -106,  -119,    17,  -104,    38,    11,    72,  -118,     4,   -27,     1,    62,   -17,  -174,  -257,  -115,   -68,     6,    28,    12,  -108,     1,   -39,   -39,    89,    43,    10,   -97,  -102,     4,    19,     1,    -4,    89,    15,  -127,   -28,    -7,    65,    19,   -62,  -188,  -218,   -77,   -41,    91,     5,   -26,   -13,    50,   -55,    41,   -22,   -52,   -41,  -101,   -91,    22,   -17,     7,   -10,    19,    -9,   -52,   -24,   -30,   -26,   -63,   -86,  -147,  -104,   -20,    24,     6,    20,   -45,   -81,    38,   -28,    -7,   -43,   -18,   -38,   -75,   -67,   -13,    -2,    -6,    17,    20,    -4,   -91,  -110,   -73,  -121,  -174,   -92,   -74,    15,    36,   -15,     7,    -8,   -56,   -64,   -14,    36,    32,     2,    28,   -32,   -92,   126,    -2,   -20,    14,     4,    -7,   -22,  -132,   -57,   -67,   -89,  -124,   -84,     9,   -29,     4,    28,    48,   -22,    38,   -35,   -68,    34,   -61,    94,   -35,    -2,   -96,    19,    15,   -10,    -4,   -17,    -5,   -25,   -93,     0,    17,  -113,   -55,   -21,   -62,    49,    16,    20,    -3,    -2,   -63,   -14,     9,   -35,     0,    45,   -75,   -16,   -91,    40,    -3,   -20,    15,    -2,     1,     2,    24,    50,     5,   -66,     6,   -11,    74,     1,    56,    33,  -101,    50,   -14,   -27,     1,   -56,  -109,    50,    19,   -31,  -118,    19,   -62,    13,     5,     5,    -1,    -8,    10,   -29,    38,    35,    26,   -14,    -5,    44,    92,    63,    13,   108,    39,    70,    -3,   -29,    25,   -30,    24,    -2,  -117,    39,   -23,    18,   -12,    -1,    12,    -4,   -27,   -16,   -53,    12,   -60,     1,    -4,   -85,    -3,   120,    81,   -24,   -46,     8,    27,   -48,   -79,     8,    45,    27,    23,   -23,   -14,   -15,     9,   -17,   -17,    -2,     4,    22,    49,   -23,    29,    77,    68,   -23,     5,    25,    64,   -27,   -49,    30,    83,  -100,   -18,    -4,   117,   114,   107,   -19,    -3,   -16,    13),
		    48 => (  -16,   -14,    -3,    -5,     5,    18,     9,   -14,   -13,   -10,    -4,    14,   -11,    -8,    -4,   -18,    14,   -19,     3,   -15,    12,     5,   -13,     9,     3,     7,    12,    16,    17,     2,    -2,    19,   -16,    -7,    -3,   -16,    -1,   -15,     3,   -12,    -4,   -12,   -29,   -14,   -51,   -24,   -30,    -1,    17,    -1,   -19,   -12,    15,    -8,     7,    -8,    16,    15,     0,     8,     2,     0,    -9,   -20,   -63,   -74,  -109,   -85,    15,     6,    12,   -54,   -54,    -4,   -26,    14,   -78,   -69,   -65,   -30,   -42,   -15,    17,   -10,   -20,   -16,   -18,     4,   -33,   -57,   -86,   -77,   -53,   -57,   -65,    21,    59,    43,    14,   -42,    -3,   -22,    71,    24,     9,   -14,   -16,   132,    13,    18,   -33,    19,    15,   -11,    17,   -48,   -82,  -122,   -88,   -93,   -42,    18,   -34,   -21,   -51,   -74,     1,   -62,   -21,   -31,   -54,    66,   159,   182,    45,  -116,  -122,   -43,    54,   -14,     0,     3,   -44,   -29,  -103,   -57,   -47,   -18,   -15,   -51,   -36,    14,     3,   -63,    -5,  -157,  -114,   -81,  -109,    22,    95,   127,    61,   -50,   -82,   -32,    13,   -16,   -12,     0,   -40,  -135,   -21,   -50,   -16,    11,   -78,   -27,   -25,   -21,   -35,   -30,   -43,   -76,   -32,   -23,    11,   -33,   -27,    -9,   -18,   -41,   -97,   -61,     3,    24,    -2,   -32,   -24,   -82,    -5,    -2,     1,   -19,    -6,   -47,   -52,   -73,   -97,     2,     7,    27,    14,   -52,    -5,   111,    14,     2,    33,   -25,   -95,   -49,    31,    50,     1,   -72,   -27,    35,    27,    26,    24,    -7,   -14,   -56,   -77,  -120,  -107,   -96,   -30,    29,   -44,    44,   -19,   -52,    17,   106,    89,   -12,   -69,    16,    42,    95,    -1,   -46,   -63,   -36,    36,    -1,    27,    41,   -20,    20,   -12,   -78,  -115,  -175,   -78,   -46,   -42,   -20,    -4,   -18,     9,    45,   -16,   -28,   -25,   -41,   -22,   -10,    18,   -44,   -81,   -80,     7,    46,     3,    -6,   -40,    47,   -25,   -33,   -99,  -120,   -58,   -20,    44,    34,   -26,    66,    81,     7,   -19,   -25,   -30,  -102,    -5,   -41,    -7,     4,   -47,    60,   -43,     5,    30,   -29,    13,    43,    46,   -26,   -21,     2,   -35,  -121,   -26,    79,   -21,    10,    38,   -22,   -74,   -67,   -97,   -60,   -10,   -35,     4,    15,   -50,   -48,   -32,   -13,   -42,   -52,   -97,   -25,    37,    99,    17,   -71,  -101,   -98,   -10,    46,   -45,   -32,    13,     0,   -48,     5,    13,   -34,   -56,   -48,    -1,    -1,   -60,   -56,   -96,   -33,   -29,   -12,    -1,    45,    23,    98,    49,    28,   -88,   -76,    12,   -33,  -147,   -47,   -49,   -35,    -8,   -19,   -73,   -60,    11,   -15,   -17,   -22,   -40,   -81,   -58,   -74,  -134,   -89,    26,   -65,   -23,    34,    24,    45,   -36,   -60,    19,   -81,  -102,  -113,  -101,   -36,   -78,   -53,  -102,   -36,  -121,   -48,   -23,    -7,   -31,    33,    -3,    -7,  -105,   -91,   -79,   -63,  -121,   -22,   -30,    60,    50,    52,    34,     2,  -106,  -125,   -94,   -22,   -65,   -44,   -36,   -19,   -88,   -80,   -19,   -25,   -37,    48,    -8,   -45,   -65,   -83,   -16,   -73,   -50,   -19,   -50,    37,   -66,   -24,   -24,    -3,   -96,   -45,   -70,    31,   -71,   -59,   -42,   -48,  -103,   -82,   -12,   -26,   -59,    53,   -12,   -59,   -92,   -83,  -159,  -163,   -29,     3,    45,    58,   -71,   -47,   -97,     8,     7,   -64,    41,    47,    93,   -20,   -60,    -9,   -11,   -49,   -34,   -18,   -28,   -24,   -24,   -51,  -115,  -105,  -106,   -66,   -14,    37,   104,   -35,     4,    42,   -39,    65,    19,    16,   -22,     3,    40,   -27,   -47,   -30,   -29,   -29,    10,    15,   -20,   -31,   -17,   -43,  -104,   -87,   -80,   -40,   -39,     5,    97,   -60,    -9,    50,   -84,    84,    82,    22,   -33,   -33,    13,    29,   -66,   -25,   -75,   -28,    17,    18,   -34,   -19,   -60,   -46,  -132,  -108,   -56,    -7,    56,    79,    64,   -45,   -54,    15,  -123,    94,   -51,    56,    20,    -5,   -10,    12,   -30,   -35,   -90,    -1,   -34,    -9,   -21,   -18,   -59,   -74,  -149,  -134,   -72,   -31,    47,    59,    19,   -75,   -31,   -12,     2,     1,    -1,    53,   -12,    19,    31,    19,  -111,   -23,   -74,    15,   -23,     5,   -36,   -14,   -28,   -73,  -189,  -149,  -136,  -104,     7,    10,   -25,    28,   -45,    16,   -37,   -95,   -40,    -9,    12,    82,    18,   -75,   -66,    -6,   -55,   -24,    12,    16,   -43,   -50,   -16,   -48,   -77,   -65,  -115,   -81,   -22,   -77,    -5,   -24,    -8,    21,   -10,    36,   -52,   -10,    89,    24,    75,   -15,    10,   -18,   -44,     3,    -6,     7,    -9,     1,   -18,   -45,  -114,  -114,  -119,   -53,   -15,   -41,   -80,  -118,   -79,   -40,    79,   -64,    19,    12,   107,   -19,   -41,   -37,   -71,   -32,   -13,   -13,   -18,     1,   -51,   -12,   -49,   -57,   -44,  -113,  -103,   -95,   -66,   -83,   -66,   -73,   -14,    91,   112,    58,    67,    33,    33,   -41,   -16,   -16,   -14,    -9,    -4,    13,     0,   -17,     6,   -71,    -3,   -38,   -63,   -26,   -16,   -61,  -119,   -67,   -60,   -82,  -137,  -107,   -73,   -35,   -20,  -124,  -141,   -49,   -65,   -21,   -15,    -6,    11,   -20,   -12,   -10,    10,     3,   -16,    -7,   -17,   -15,   -25,   -27,   -25,   -37,    10,     5,   -46,   -28,   -57,   -62,    -1,     3,    -8,   -19,    -2,   -18,    17,    12,    20,    -8),
		    49 => (  -11,   -10,     5,     4,     6,     5,    13,   -15,    -7,     8,     0,    10,     3,    -4,    -2,    -7,     6,    14,     8,     7,    15,   -19,    -4,    11,   -16,    16,    -3,    12,    10,     2,     7,     8,    -1,    -1,    14,    -4,   -20,   -14,   -25,   -53,   -52,   -45,    -5,  -145,  -132,  -114,   -43,   -18,    13,   -25,    -2,   -19,    19,    -4,    -8,   -17,   -19,    10,   -11,   -34,   -25,     4,   -21,   -60,   -57,   -33,   -35,   -88,   -41,   -46,  -113,   -49,  -104,   -27,    -7,   -26,   -75,   -18,   -19,   -48,   -13,    17,     5,    -1,   -10,    20,    -9,  -162,   -48,   -46,   -21,   -84,  -100,  -128,  -118,  -117,  -229,  -159,  -187,  -179,  -170,   -82,    23,   -87,   -90,   -67,   -40,   -18,   -31,   -30,   -17,    13,     3,    11,   -48,   -53,   -52,  -119,  -164,  -117,   -91,  -159,  -120,  -219,  -258,   -59,  -148,  -104,   -62,    15,    51,  -269,  -141,  -179,  -102,   -25,   -21,  -111,   -99,   -25,   -13,    13,   -31,   -52,   -12,   -60,  -122,  -102,  -112,  -105,   -63,    17,   -39,    57,   -65,   -25,   -96,   -88,   -83,   -76,   -44,   -53,  -169,  -144,   -92,   -85,   -75,     7,   -16,   -28,   -38,  -146,  -172,  -355,  -179,   -23,     3,   144,    31,    60,   -19,   112,   -15,    14,    24,    52,    72,     1,    48,    40,  -107,  -110,  -168,  -153,   -96,   -64,    19,   -89,  -121,  -155,  -273,  -342,   -23,  -106,   -41,    21,    54,    64,   107,    25,   -30,    83,   -13,    49,    28,     4,   -17,     3,   -58,  -152,  -155,  -130,   -99,   -37,  -148,  -107,   -94,   -93,  -170,    -5,   -15,  -104,    16,   -44,   -27,    -2,     2,   -71,    -4,   -54,    -7,   -18,    46,   -46,    -5,    55,   -60,   -64,   -96,  -149,  -136,   -64,   -29,   -56,   -11,   -50,  -161,   -13,   -21,    -2,   -40,   -72,    -5,    31,    -7,   -27,   -50,    95,   -35,   -46,   -52,    21,     1,    51,     1,   -27,   -56,  -143,  -148,   -54,   -18,  -106,  -162,   -11,    34,    17,   -63,   -56,   -32,    37,   -27,    37,    30,   -56,   -74,   -77,   -31,    45,   -26,    34,    59,    21,    44,   -29,   -76,   189,  -150,  -103,    12,  -245,    75,   -27,    83,   -24,   -46,   -31,    44,   -23,    94,    15,    16,    23,   -63,   -32,    11,    98,    25,    29,    64,    69,   139,   -70,    17,   194,  -118,  -117,   -21,   -58,    40,    41,   149,    34,    19,    54,    10,   101,    -4,    49,  -104,  -123,    20,     5,    35,    99,   121,   135,    47,    89,   101,   145,  -156,  -298,  -178,   -33,    11,  -115,   -88,    16,   196,   152,    53,   116,   106,    64,    74,     8,    30,    31,    63,    49,   118,     0,    51,    81,   110,    80,   218,    43,  -255,  -159,  -110,    -1,   -43,   -93,   -55,    34,   151,   124,    33,    50,   129,    36,    88,   -42,   -52,    33,   -26,     2,    81,    15,    57,    99,   -14,    44,   240,   -15,  -359,  -239,   -21,   -13,   -16,   -15,  -197,    42,   139,    14,   -64,    57,   153,    81,     9,   -87,   -66,    25,   -49,    78,    74,   128,    91,    82,   -44,   -85,    -8,   -85,  -319,  -184,    75,   -35,    14,   -17,  -175,  -107,    27,   -89,   -12,   -12,   -19,   -81,    96,   -81,   -40,   -43,   -41,    -7,   -19,    10,   -15,   -49,   -32,  -149,   -42,   -78,  -269,  -144,   -29,   -99,    13,     0,  -202,    -6,   -71,   -79,   -74,    17,   -10,   -45,   -43,  -121,   -28,   -57,   -60,    33,    17,    38,   -64,   -84,   -82,   -78,   -77,   -65,  -215,    -9,   -35,   -69,    88,    -5,  -189,    23,   -72,  -116,   -52,   -21,    11,   -18,    19,   -26,   -71,  -133,     0,   -29,   -22,    -7,    33,   -13,  -101,    20,   -13,  -170,  -369,   -37,   -96,   -59,    13,   -24,  -101,   130,   -59,  -138,  -116,  -126,   -85,   -99,   -89,   -69,  -105,  -225,   -39,   -14,   -61,   -52,   -28,    43,   -12,   -60,    64,   -86,  -167,   -18,   -79,   -29,    20,    -2,  -181,    97,   -54,   109,   -62,  -266,  -205,  -123,  -152,   -29,  -126,  -141,    29,   -50,    18,    19,   -57,    39,  -111,   -75,   -40,   -30,    23,    67,   -45,   -14,    -8,     3,  -181,   121,    32,   114,   -59,  -110,  -117,  -105,  -155,  -124,  -125,    -6,  -158,   -65,    19,   -60,   -99,   -58,  -126,   -35,   -59,  -132,   -64,    51,  -311,   -13,    18,   -20,  -166,   105,   -92,   -40,    27,    81,    85,    -7,    37,   -61,   -27,     0,     6,    31,   -44,   -70,   -95,  -144,   -50,   -21,   -24,  -140,    13,   -45,  -186,   -39,     7,     7,  -131,    89,   -26,   -64,   -53,    21,    -4,   -65,     7,   -76,   -56,    -3,    -5,   -88,   -72,   -55,   -51,   -33,    -9,    59,    63,   -37,    -3,    -7,   -29,    17,     2,    12,  -127,  -132,   -21,    65,   -87,    47,   -33,   -17,    29,    71,   -30,   -56,  -125,   -16,    18,   -80,    13,    38,   -58,    14,    92,   114,    -3,   -45,   -64,    -3,   -16,    12,    90,   -88,   115,    48,  -149,  -177,   -58,   -35,  -117,   -92,    32,   -14,   121,    -3,    55,    92,    89,    58,   134,   162,    30,   -24,   -48,    -5,   -74,    19,    -4,     4,     1,    69,    85,    -1,    29,     6,    27,    29,   -74,   -19,    90,    25,   126,    26,    56,   137,   178,    48,   129,   124,    71,    75,    73,    19,    19,   -10,   -14,    -5,    -6,    -3,   -92,  -114,    43,    27,    57,    38,   -18,    36,    13,   -57,    86,    69,    46,  -158,   -53,    85,    10,   -97,    33,   -93,    13,   -13,     0,     6),
		    50 => (   -3,   -11,     9,    13,    15,    -7,    -1,     3,    13,    12,    -5,    11,   -11,    18,   -19,     8,     1,   -10,   -12,   -11,   -15,   -15,    19,   -20,    12,    20,     4,   -14,    -4,   -17,    18,    16,    19,    10,     9,    16,    17,   -13,    -6,     6,    12,    20,   -11,    12,   -14,   -16,     1,    12,   -14,   -17,    19,   -13,   -16,    -7,    16,     4,     5,    -7,    -4,    32,    52,   -32,   -30,   -22,   -39,   -50,   -70,  -118,  -131,  -134,   -69,   -97,   -75,   -77,   -34,    14,    17,    -3,   -84,   -18,     7,     6,   -19,     2,    15,   -19,     8,    12,    -4,    28,   -47,   -31,  -134,  -131,   -44,     2,     0,    48,    -7,  -105,  -133,   -61,   -37,   -10,   -30,   -12,   -35,   -20,    -9,   -17,   -17,    17,   -14,   -14,    -5,    15,   -35,  -113,    71,   -13,    78,    84,    45,    60,   -27,    -9,   -14,   -85,   -17,    39,    46,     9,   -92,  -131,   -31,    -7,   -18,   -10,   -38,    -4,     4,    12,     3,    34,    18,   -70,     1,   -36,  -115,   -21,    25,    54,    21,    56,    31,    -9,    49,    14,    34,   -23,   -29,   -30,    -4,   -19,   -62,   -84,   -67,   -83,     8,    10,   -55,   -27,    40,   -32,     1,   -49,   -51,   -20,    23,    27,     4,    -4,    11,    23,    82,    35,    45,   -29,   -22,   -87,   -36,   128,    79,   -99,  -106,   -23,    12,   -26,   -50,   -29,   -43,    57,    46,    29,   -22,    42,    85,    21,    21,     0,    39,     6,     3,    55,    -8,   -32,   -91,   -74,   -50,    49,    61,   -73,   -82,    35,    24,    -1,    15,   -52,   -49,    -3,   -11,     7,    73,    80,   -21,   -13,   107,    55,    68,   -40,    12,   -55,    -6,   -50,   -10,   -39,    27,     8,    18,   -79,  -112,   -47,   -10,     0,     1,   -33,   -89,    81,   -74,    -6,   -14,    31,    -6,    -2,   -32,    -9,    10,    13,   -59,   -88,    92,    89,    96,    41,    68,    -4,   109,  -124,  -106,   -15,    15,   -13,     3,   -35,  -128,    15,     1,   -13,    38,    21,    60,   -13,  -117,   -48,   -15,   -18,   -66,    41,    58,   -29,   -78,   -41,   112,    25,    98,   -81,   -71,   -15,    -1,    44,   -59,   -71,  -101,    -9,    16,   -11,     8,    17,    54,  -106,  -115,  -115,   -94,  -117,   -36,   -14,    -1,   -86,   -59,   -83,   -52,    17,    66,   -43,   -12,   -19,    20,    10,     7,   -47,    -4,   -74,    25,   -33,     4,   -22,   -75,   -27,   -84,   -77,   -77,   -99,   -68,   -38,   -79,    16,   -21,   -41,   -15,  -114,    14,   -38,   -80,   -36,    -2,    40,    12,    18,    92,    -9,     4,    -4,    96,    24,   -67,  -173,  -164,  -235,  -191,  -129,   -96,   -86,   -17,   -67,     2,   -13,    17,   -76,    -7,   -21,   -40,   -34,   -13,     5,   -12,   -53,   -49,   109,    53,    88,    37,    27,   -63,  -231,  -166,  -196,   -77,  -114,  -164,  -128,   -34,    11,   -53,    13,   -41,    50,   101,    -7,   -79,     4,    20,    10,    -4,  -130,    32,    96,   105,   -30,    15,    56,    53,  -140,  -259,  -152,   -50,   -71,  -102,  -100,   -69,   -10,   -24,    32,    13,   -34,    28,     1,    -9,   -62,    20,    -1,   -16,  -154,    80,    94,    11,   129,   -61,   -22,    21,   -73,   -62,  -134,    -8,   -80,  -189,  -157,  -130,  -109,    37,   100,    18,    -4,   -16,   -42,   -56,   -12,   -10,     7,   -38,   -27,    52,    77,    45,    10,   -31,   -46,    51,   100,    46,    36,   -46,  -208,  -262,  -143,  -183,   -89,   -34,   -19,   -29,    14,   -60,   -62,  -105,    14,    -1,     4,   -22,    47,   -68,    74,   119,    76,    23,    25,   -36,   -29,     7,   -74,  -118,  -168,  -206,   -90,   -39,   -16,    94,    51,    46,    24,    24,   -52,   -73,   -31,    -1,     0,    12,    20,     8,    66,   -18,    20,    19,   -36,   -27,   -21,    46,   -31,   -32,   -81,    -4,    63,   -85,     4,    47,    73,    79,     4,     8,   -55,    -9,   -25,    -4,    11,   -12,    22,   108,   133,   -52,    -6,   -49,   -95,   -75,    18,    39,   -20,    -9,    -1,    26,    40,    18,   -14,    38,    50,   -44,   -15,    21,   -67,   -18,   -15,    12,   -31,     0,    96,   142,    29,    84,    24,   -82,   -27,   -59,   -12,   -60,   -27,    66,    65,   -49,    -7,    -4,   -10,    -3,    60,    85,   -23,   -26,   -21,     1,    44,     0,    -5,   -17,   -22,    23,    68,    70,   105,    74,   -21,    20,   -31,   -10,     0,    28,    24,    29,    33,    -2,   -35,    12,   -20,    36,    22,   -63,     5,    -3,    26,     1,   -19,   -16,   -95,   -96,    20,   -40,   -66,     4,    -6,    27,     9,    69,     3,   -25,    53,    -1,    73,    12,     1,   -86,   -85,   -37,   -35,  -147,     5,   -33,     3,    11,   -20,    -7,   -26,   -53,     6,    40,    34,   -18,    77,    98,    20,    35,    69,   -57,    37,   -20,    77,    47,    74,   -83,   -98,   -97,   -45,    35,    36,     3,   -16,   -15,   -11,     8,    -9,    -7,   -33,   -23,   -22,   -36,    -5,   -24,   -96,   -72,   -66,  -100,  -157,  -176,  -179,  -228,  -149,  -114,  -138,   -77,   -10,   -40,   -16,    17,    13,    15,   -18,   -14,   -12,   -21,   -38,   -49,   -36,    12,   -50,   -40,   -52,   -23,  -105,   -89,  -160,  -113,   -93,  -132,  -138,  -105,  -122,   -73,   -84,    18,   -20,   -13,   -16,     6,     1,    10,   -13,   -18,   -14,   -12,    11,   -16,    -7,    -9,    -4,   -25,    13,    -8,    -9,     0,   -25,   -18,   -21,   -20,   -81,   -68,   -89,   -17,    19,    16,   -19),
		    51 => (  -18,   -20,    -7,   -11,    -7,    20,     8,    -4,     7,    11,     8,     2,     9,   -15,     1,     1,    -2,    -7,     2,     4,    15,     5,    13,    -9,    17,   -12,   -19,    -6,   -18,     1,    18,   -12,   -12,     3,    14,   -19,   -18,   -20,   -14,   -10,     3,   -17,    29,    16,   -16,   -10,   -26,    11,     0,    -7,    10,     3,    11,    -5,   -12,    -8,     2,    -8,    -6,     3,     5,   -12,   -15,   -11,   -34,   -59,  -120,  -108,   -77,    23,   -84,   -28,   113,    29,  -113,  -114,   -32,   -69,   -59,   -35,   -16,    17,     2,   -17,    -5,    -6,   182,   103,     3,   -81,   -50,   -16,   -48,   -60,  -105,  -157,   -86,   -15,   -69,   -98,   -37,   -52,   -23,   144,   120,  -108,   -21,   -59,   -23,   -14,    20,   -16,     5,     7,   160,   166,   -11,   -87,   -51,   -38,   -45,  -112,  -140,   -53,   -14,    87,    79,     0,   -92,  -142,    76,    30,    45,   -44,   -21,   -37,     1,   -22,   -69,   -64,   -13,     2,   155,    83,    27,   -13,    -8,   -68,  -178,  -199,   -44,    14,   -52,    39,    12,    12,    53,  -113,   -57,   -33,   -91,   -62,   -38,   -12,   -20,   -17,   -61,   -64,     0,    -6,   -61,    18,     7,   -32,   -68,   -11,  -167,  -215,  -109,     1,    29,   104,    37,   -62,    15,  -131,   -39,  -126,  -114,   -30,   -16,    13,    -1,     2,   -49,   -51,     7,   -20,   -71,    17,   -10,   -88,  -104,   -37,  -234,  -143,     6,    37,    70,   107,    28,   -31,   -77,   -99,   -43,  -223,   -97,   -56,     3,   -15,    -7,   -31,  -127,   -60,     9,   -25,   -64,    27,   -36,   -61,   -95,   -86,  -227,  -110,     9,     0,    19,    75,   125,    75,   -97,   -83,   -57,  -221,   -64,   -52,    47,     2,   -18,   -11,   -80,   -26,    11,   -30,   -74,   -32,   -26,     8,   -54,   -43,  -116,    -4,    42,   -23,  -105,     1,   138,   107,   -84,  -154,     2,    15,   -86,    -9,    35,   -12,   -67,   -40,   -69,  -109,    -1,   -27,   -32,   -27,   -59,   -21,  -114,   -53,   -46,  -109,    95,   -10,   -41,    50,    73,   -13,   -44,  -121,   -94,    -5,   -33,  -154,    15,    58,   -89,   -43,    22,    94,     4,    17,   -10,   -29,   -27,   -61,  -139,   -76,  -129,   -86,   -24,    51,   -44,    11,   109,   -27,    -1,   -76,  -120,   -44,    60,   -17,    50,    61,   -79,   -51,   -41,   159,    19,     1,  -150,    59,     5,    -6,   -47,   -49,   -38,    92,    28,   -16,    25,    10,    64,   -47,   -14,  -134,  -147,   -75,   122,    12,    21,    77,   -87,    12,    10,   121,     9,   -12,  -146,     9,     9,   -21,   -14,    32,    98,    60,  -152,    29,    31,   -66,   -42,   -53,   -23,   -80,   -98,    38,   139,   -53,   -66,  -119,   -96,    85,    65,   -19,    -4,     1,   -11,    16,   -15,   -77,     5,    49,   -36,   -54,  -134,   -89,    34,    -9,   -20,   -62,    17,     6,     0,    13,    36,   -56,  -109,   -16,   -12,   -27,   100,    19,   -15,    -1,    15,    51,    -3,   -91,   -76,    -3,   -34,   -58,   -53,   121,    71,    98,    38,  -102,     5,   -13,    70,   -33,    86,   -39,   -95,   -30,   -95,   -57,    10,   -51,     4,   -11,    17,   -58,    -7,   -50,   -32,     5,   -34,   -76,   -46,    60,    32,    -3,    29,   -74,   -72,   -17,    26,   -78,    14,   -45,   -69,   -74,    -2,   -85,     1,   -26,    -9,    20,     5,   -29,   -24,   -94,   -69,   -97,   -30,   -57,   -61,   -40,    20,    16,    17,   -41,   -57,   -79,    19,   -84,  -103,   -65,    42,    44,   -50,   -83,   -24,    20,   -13,     3,   -22,   -18,   -51,    -3,   -69,   -36,   -95,   -60,  -200,   -42,   -66,   116,    57,    -9,    15,   -25,    56,  -130,    38,   -19,  -109,  -101,   -97,     7,    -3,    83,   -16,   -11,    14,   -17,   -20,    -8,   -24,   -60,    37,  -106,  -104,   -40,   -21,    51,   100,    52,    -2,   -72,   -43,  -170,   -52,   -56,  -144,   -90,   -39,    50,    62,    91,    20,    18,    -1,   -54,   -52,   -29,   -61,  -122,   -32,   -41,   -32,   -23,    88,    31,    43,    34,    13,   -29,   -43,   -73,     4,  -121,  -186,   -67,    -3,   -17,    89,   -14,    34,    26,    12,   -46,   -51,   -21,   -83,  -183,   -11,    -3,   -51,     2,     8,    14,   -21,     6,   -31,  -114,    82,   -29,    36,   -40,  -137,  -123,   -55,    31,   -34,    -7,    46,    20,    16,    16,   -35,   -23,   -34,  -149,    12,    -9,   -26,   -67,   -47,   -12,    14,   -27,   -31,   -44,    44,    18,    74,   -11,  -115,   -48,   -97,    79,    62,    -5,    13,     2,   -23,   -52,   -18,    18,    74,   -52,    21,   116,     8,    66,   -19,     6,    -4,     7,    25,   114,    95,    29,    65,   -42,   -22,   -64,   -71,   -21,   149,    14,   -15,   -14,   -14,   -26,   -21,   -19,    96,    17,   -14,    17,    83,   115,   -17,  -101,   -95,  -134,  -173,   -66,  -130,   -82,   -76,   -45,  -120,   -11,   -72,   100,    84,    15,    14,    -4,   -16,     2,   -11,   -13,    -6,   -18,   -28,   -57,  -255,  -207,  -144,  -124,   -34,  -160,  -152,  -169,  -141,  -147,  -240,   -93,   -72,   -68,    -4,    -9,   -18,     9,    15,   -18,    -8,    -6,   -57,  -118,   -87,   -76,   -75,   -64,   -52,   -72,  -120,  -126,  -133,  -128,   -94,   -94,   -24,   -54,   -10,   -62,    -6,    -7,   -13,     9,    -4,     5,   -16,    -5,    18,     0,   -18,    14,     1,     4,   -14,    19,   -11,   -13,    -5,   -15,   -27,   -21,    -3,     3,    12,   -12,     2,     6,     4,     2,   -14,   -18,   -12,   -20),
		    52 => (    5,    11,   -11,   -16,     9,     5,   -19,    15,   -10,     1,    13,    19,   -27,   -23,    16,    37,     7,    16,    15,    -7,     5,   -17,    12,   -14,     5,    20,     8,    -5,     6,    -6,    17,   -20,    19,    19,   -19,   -13,   -10,    12,    17,   -13,    12,    16,   -37,   -27,    21,    28,   -13,   -84,   -41,    -6,     5,    10,    12,    12,     8,    20,   -10,    -5,   -28,   -31,   -28,    19,   -23,   -35,    79,   119,   143,    71,    60,   -40,     0,   -54,  -145,  -107,    -5,    39,     4,    40,   -41,    31,    61,    36,   -17,     5,   -16,   -12,   -32,  -121,   -97,  -109,   -33,   -59,    40,    41,   -18,   -21,   -46,    26,    55,   -26,    -7,   -15,   -24,    95,   -29,   -22,   -33,  -146,   -75,    34,   -38,     1,     0,   -12,   -20,   -34,    89,   -22,   -15,    16,     3,    22,   -35,     2,    57,    22,    -8,    40,   -62,    33,   -74,   -25,    50,   -77,   -39,  -133,  -142,    62,  -105,   -49,   -12,   -15,     2,   -46,    15,  -115,  -127,  -170,   -82,   -13,    84,    11,   -58,    48,    29,    22,   -50,    25,   -18,    -4,    -2,    27,    -8,    67,  -115,   117,   -86,   -11,   -12,     3,     4,   119,    94,  -102,   -79,   -43,    38,    79,    78,     6,    12,    92,    21,    -1,   -36,    21,     7,   -15,   -32,   -84,   -30,   -19,     9,   -92,   -93,   -13,     4,     0,   -30,   154,   116,    82,   -30,    19,   -25,     5,   -20,    36,    26,    48,    12,    59,    73,    67,    22,    56,   -34,   -59,    99,    12,   -80,   -94,   -76,   -63,   -57,   111,   -18,   113,    74,    62,   -81,   -31,   -38,    59,     4,   -16,   -31,   -59,   -24,    14,    57,    84,   -14,    95,   -67,    -2,    90,    82,  -220,  -136,   -95,   -67,    20,   -37,    33,    23,   -33,    23,   -53,   -58,   -28,    77,   -78,     9,    43,  -108,   -32,    17,    46,    25,   -19,    94,     4,   -55,   -58,    83,  -181,  -117,   -55,   -26,     3,    -4,    10,    64,  -124,   137,    69,   -10,   -28,     5,   -73,   -91,    -3,    51,   -32,   -34,   -26,   -43,   -12,    23,    50,   -11,   -41,    85,   -38,   -42,    17,   -24,     4,   -57,   -17,    82,    15,    29,    66,     5,   -33,   -81,  -174,    -3,   -57,  -101,  -119,   -99,     5,   -37,   -93,   -19,   -47,    -8,   -44,    40,   -14,     6,   -90,   -17,   -14,     1,  -112,    -9,    25,  -122,   -49,   -90,  -112,   -83,   -99,   -93,   -37,  -153,  -187,   -49,     2,   -20,  -104,   -21,   -68,   -31,   -18,   -58,   -27,    47,    -7,   -48,    -4,    13,     8,   -13,   -19,   -47,  -172,  -151,  -256,  -151,  -115,  -147,  -191,  -110,   -86,   -43,   -35,   -83,   -72,   -90,   -75,   -85,    31,   -68,   -18,    49,    85,   -43,    14,   -60,   -76,   -28,  -100,  -181,  -198,  -204,  -318,  -202,  -103,  -108,   -34,   -60,     2,   -43,  -114,   -40,   -39,   -35,   -88,  -139,   -16,  -156,   -16,     7,   105,    56,    15,   -53,   -12,   -46,  -191,  -103,   -93,  -134,    24,   -12,   -49,    51,    -3,    64,    19,   -97,    14,   -16,  -118,  -136,  -135,   -80,  -149,   -78,    35,   -45,   120,   169,     1,    -4,   -75,  -122,  -217,   -76,   -88,   -63,   -32,    34,    39,    42,   -70,    28,    35,   -42,   -62,   -25,   -57,  -124,   -85,   -34,    56,   -47,    49,   116,   154,   103,   -15,   -11,     7,   -87,   -75,   -95,    -9,   -26,    -5,     9,    48,    19,   -67,   113,    72,     2,   -18,   -28,   -17,  -107,   -65,   -37,   -30,   -38,   -85,   198,   115,    94,   -11,   -14,   -29,  -168,   -59,   -45,    53,    77,   -33,   -50,    15,    -6,    36,   -11,   -16,   -24,   -17,    51,   -61,   -80,  -100,    63,    78,    76,   145,   240,   -14,   126,   -11,   -36,    35,   -83,  -100,   -34,    78,    50,   -52,   -77,    38,    23,     8,   151,   132,    38,    64,   -13,   -30,   -63,    11,    80,    35,    73,   -22,    68,    63,   129,     7,   -18,    76,    -9,    -9,   -53,   182,    60,    43,    56,   127,   106,    76,   206,    72,    57,   115,   -12,   -22,   -19,   124,   115,    45,    33,    24,    95,    43,     2,    14,    40,    39,    96,    31,    25,    92,    61,   -23,    53,    42,    48,     7,   154,   122,    95,    60,    81,    37,    59,    67,    55,    94,   202,    94,    94,    93,   -26,    10,    -7,    -4,     0,   -11,   100,   140,    75,    18,    81,    19,    32,    20,    11,    51,    40,   -38,   -88,    -5,   -84,    32,    88,   149,   176,   141,   -13,  -132,   -42,   -16,   -16,    14,   -94,   -50,    28,   104,    55,    40,    92,    39,   132,    98,    70,    25,   -27,   -83,   -55,   -61,    -3,    73,   103,   186,   130,   104,    15,   -68,     6,     8,    -1,  -101,   -70,   -24,   -57,     5,    55,   139,   -41,    12,    10,    91,   -43,    58,    27,   -98,   -31,    -4,     3,  -111,   -61,    -9,   105,   210,   117,    66,     5,    14,    -4,   -65,    -9,   -84,  -203,    93,   -31,  -105,  -206,  -267,   -79,   -41,   -17,    90,    66,   -67,    24,  -138,  -178,   -16,    27,  -147,   -66,    36,   110,    75,    -7,    13,   -15,   -12,    -4,   -68,  -125,  -140,   -91,   -88,  -133,  -229,  -185,  -107,  -118,  -120,   -73,  -178,  -166,  -133,   -13,   -58,   -76,   -47,     6,   -19,    -2,   -18,    13,   -20,    16,   -16,    10,   -10,     0,   -25,     2,    17,    -5,   -61,  -102,    -7,   -42,   -10,    -4,     4,   -22,   -12,     8,   -38,   -69,   -34,    -8,    -9,     4,     0,    -2),
		    53 => (   -6,    -9,     5,   -11,    -6,   -13,    20,   -20,    11,     5,     4,   -15,   -20,   -17,    -6,    -4,   -13,    -8,    -9,    -7,    18,   -14,   -15,    -6,    13,    -8,     0,     1,   -11,    -2,    13,     2,   -11,    -6,    13,    -9,    18,   -20,     4,    -6,   -16,   -14,   -37,   -10,   -46,   -20,     1,   -12,     0,     3,    17,     6,    16,    19,     5,   -19,    13,    19,     6,   -14,     5,    12,    12,     2,   -79,   -94,    67,    82,    55,   -36,   -78,   -80,  -117,  -119,   -83,   -41,   -16,   -55,   -64,   -88,   -27,   -18,    -5,     0,   -11,     2,    -5,   -46,   -19,    -4,   -29,    37,    17,   -22,    62,    67,    46,    51,    12,   -50,    29,    63,    75,   -33,   -31,   -46,   -18,  -146,   -66,   -15,    -5,     3,   -14,    36,    10,    -1,   -26,    17,    21,    53,    24,   -19,   -37,   -65,   -90,   -99,     0,   -41,   -47,  -121,   -56,     3,   -77,   -64,    79,  -161,  -135,   -71,   -22,    -5,    -1,    10,    18,   -31,   -16,    57,    79,   132,    13,   -90,  -130,   -62,   -45,   -55,    -1,   -22,   -15,   -17,   -23,    20,   -21,   -54,   -76,   -61,   -59,   -17,   -57,   -18,     2,    28,    -4,    37,    12,    -2,    15,   -17,  -106,   -75,    61,   -18,     9,   -36,   -58,   -38,   -17,    -2,     3,   -81,   -65,   -29,   -28,   -22,   -23,  -126,   -72,   -28,    18,    38,    55,   -79,  -180,   -74,     3,   -56,   -93,   -37,   -37,    14,   -32,    -3,    11,    11,   -19,    43,    -8,   -82,    19,   -52,   -13,   -69,   -45,  -101,   -74,   -32,     2,   -20,    48,  -110,  -149,     1,   -50,   -80,   -47,    29,    29,   -21,     6,   -59,    15,   -46,    10,     7,    68,    17,    35,   106,    62,  -141,  -235,   -77,  -102,     3,   -13,   -91,   -75,   -86,    15,     8,    53,   -10,   -28,   -34,    46,    74,   110,    57,    51,   -34,   -55,   -38,   -61,   -39,    69,    44,    44,  -110,  -281,  -113,  -114,   -18,    -2,   -97,   -44,    64,    29,    24,   120,    11,   164,    77,    87,    70,    -3,    -5,   -18,   -51,  -140,    -9,    59,    63,    43,   -20,    54,   -33,  -261,   -25,   -82,     9,    -9,  -100,   -43,   148,   134,   126,    29,    79,    48,   109,    41,   -77,  -166,  -161,  -135,    45,    32,    43,    68,    84,   130,    24,    30,    -8,  -156,  -145,   -32,   -20,    -9,  -100,   -88,   151,    85,    60,     1,    34,   -97,   -91,  -127,  -284,  -208,   -47,    70,   125,    44,    16,    61,    -7,   -29,   -67,   -44,   -97,     1,    14,     2,    14,     9,   -66,  -188,    63,   -96,   -64,   -48,   -60,  -131,  -265,  -274,  -174,   -36,    45,    93,    20,    23,   -11,   -56,   -73,   -49,   -29,  -143,  -109,    86,   -50,   -46,   -14,   -33,    28,   -29,   -50,  -127,  -152,  -219,  -202,  -199,  -102,   -44,   -78,    44,    71,    38,    29,   -23,    19,  -102,   -65,   -86,   -61,  -151,   -30,   126,   -34,   -72,   -46,    -9,    65,    29,    17,   -43,   -78,  -168,  -222,  -164,    -7,    41,   -35,    52,   107,   175,    -1,    58,   -21,   -26,    -8,   -34,     7,   -74,   -41,    98,   -39,    87,    16,    -1,    15,    49,    96,    21,   -62,   -90,   -62,  -132,   -88,   -95,  -182,   -22,    15,   -35,   -87,    58,    41,   -54,    10,    12,   113,   -26,   -83,    55,  -104,    37,     5,    -4,     9,    22,    22,     7,   -10,   -35,   -85,  -170,  -220,  -275,  -303,  -368,  -299,  -191,  -116,    72,   -20,   -92,    67,    56,   111,    36,   -77,   -32,  -137,   -18,    -7,   -37,    14,   114,    29,   142,    13,   -63,    -1,   -27,  -143,  -132,  -199,  -288,  -221,  -135,  -127,   -10,    89,    67,    72,    24,   -18,    47,   -32,  -177,   -51,     9,   -46,    -4,   -59,   -72,   -61,    37,    61,    -3,     3,   -49,    39,   -21,   -65,   -48,     1,     6,   -39,   -37,     5,   -44,    -1,    18,     6,    84,    -1,   -55,    33,   -26,   -42,    12,   -14,   -70,   -11,    36,    66,    77,    53,    16,    91,    78,   112,    48,     1,   -36,  -107,   -41,   -76,   -61,    16,    75,   -14,    26,   -65,   -83,   -58,   -16,   -21,   -11,    45,   -32,     4,   -31,    42,    20,    79,    89,    29,     6,     1,    14,   -37,     5,   -76,   -72,  -109,   -26,    34,    53,     0,   -41,   -59,   -94,   -40,   -35,    -1,   -20,    11,   -50,    10,    12,   -26,   -48,   -65,    -9,   -16,    19,    12,    25,    26,    35,   -20,   -11,     7,   -11,    70,    -8,    17,  -109,   -99,   -87,   -42,   -27,    14,     3,     9,    55,    80,    90,    61,   -23,   -37,   -25,   -19,   -99,   -41,   -74,   -28,   -34,    57,    13,    51,    57,     1,    26,    44,  -110,   -88,    77,    48,     4,     4,   -10,   -10,    -5,    66,    81,     0,   -71,   -38,    12,    51,     3,    16,    43,    10,     8,   -36,    72,    66,   -40,  -111,   -28,   -37,   -80,  -127,   -82,   -50,   -24,     1,    -4,    16,     4,   -86,   -67,    27,    49,    27,   -47,   -41,  -143,  -123,   -97,  -181,  -120,    -7,    -3,   -95,   -97,   -97,   -55,   -65,   -59,  -111,    -4,     2,    12,     3,   -13,    -1,     4,   -62,  -151,  -139,  -102,  -114,  -151,  -134,  -191,  -163,  -139,   -71,   -52,   -58,   -82,  -198,  -182,  -154,    -9,   -64,   -15,    -4,    12,     8,    -1,     6,    -6,   -13,   -12,   -18,   -13,   -29,   -26,   -36,   -30,   -96,   -72,   -89,     0,   -67,   -62,   -83,   -64,   -66,   -62,   -90,   -39,   -22,   -14,    -3,   -11,    -6,    19,     6),
		    54 => (   -9,    -9,   -10,    14,     5,   -10,    10,    -2,    -6,   -20,     7,     2,   -24,   -25,   -25,   -19,    15,   -19,   -19,    -3,   -19,   -19,     7,   -15,   -19,   -12,     8,    14,    -5,    18,    13,    17,    17,    -9,   -85,   -70,   -21,     4,   -38,    -4,   -33,    24,    75,   -17,   -19,   -11,   -19,   -11,   -42,   -28,   -26,   -17,   -18,    19,    -2,    -1,   -18,    -3,    -9,   -33,  -118,    -9,   -51,   -84,  -126,   -41,   -28,   -20,   -37,   -80,   -63,  -110,  -150,   -61,   -38,   -18,   -96,   -79,    -8,   -25,   -16,   -59,    -3,     2,     2,     2,   -35,   -54,   -93,   -32,   -68,   -89,   -40,   -17,   -45,   -25,    11,   -43,   -77,   -12,    14,    57,   -72,   -53,   -73,   -27,   -44,     2,   -11,   -38,     9,     2,    12,     4,   -32,   -22,   -38,   -57,   -94,    53,   119,    62,   -49,  -147,  -189,  -117,   -98,   -91,  -159,  -198,  -205,  -131,   -59,   -46,    16,   169,   124,    76,  -147,   -28,   -17,   -15,   -45,    16,   -54,    -5,   -51,    42,   174,    50,  -108,  -187,  -128,   -73,   188,   107,    78,   -34,  -192,  -236,   -84,   -77,   -14,    52,    32,   -52,   -24,   -21,     6,    10,   -17,   -70,    71,    98,   -35,    72,    77,   -76,  -218,  -253,   -43,    27,    31,    90,    80,    24,  -183,  -350,  -316,   -34,   106,   112,    69,  -161,    39,  -114,    -6,   -64,     4,   -71,    48,    75,    38,    55,   -15,   -39,  -121,   -78,  -115,    -9,    89,    89,    59,    52,  -264,  -366,  -168,    47,   154,   167,    17,  -197,    12,  -139,   -42,   -65,    -9,   -88,    -6,    90,    56,    66,   -24,   -28,   -86,  -120,  -152,    11,    64,   141,   -50,  -179,  -326,  -169,   -27,    82,    49,   -23,   -13,   -70,    40,  -101,   -12,   -25,   -32,   -98,    27,     6,    55,   130,     1,   -60,   -81,  -153,   -56,    -4,   110,    60,   -28,  -172,  -161,   -68,    58,    63,   -26,    30,   -25,   -46,    42,   -88,     8,   -37,   -90,  -104,   -37,     3,    24,    16,  -100,    32,   -31,  -124,    47,    -9,    97,    29,   -26,  -102,  -105,    -3,    40,    -6,    10,   -64,    15,    48,   -17,   -78,   -17,     8,   -88,   -52,   -76,    36,   -24,   -32,    14,    54,    -8,    27,    30,   -94,     8,     8,   -55,  -106,   -75,   -23,    -1,    11,    28,    -2,   -72,    -6,   -61,  -138,     5,    -5,   -61,  -211,   -63,    48,   -36,     8,    25,    20,    55,   -81,    27,    22,   -13,   -54,   -65,   -58,  -100,    15,    40,    19,    15,   -88,   -16,   -59,  -158,  -116,    -8,    19,   -66,  -143,   -95,   -15,    -1,    39,    -5,    45,   125,     4,   -91,    55,   -88,   -65,    40,     2,   -25,    50,     7,    10,     5,   -23,   -94,  -127,  -148,    -8,    14,    -7,   -61,  -130,   -38,     1,    71,     5,     5,    45,    64,    11,     5,    70,    37,   -41,    -4,    62,   -32,     5,    19,    47,    51,   -53,    -5,   -86,   -39,    10,   -15,    -9,    -1,  -125,   -12,    20,    38,   103,    79,    64,    57,    42,    46,    -4,    31,   -16,   -64,    15,    14,    16,   -38,   -47,    15,     0,   -51,   -60,   -26,    27,    16,    -9,   -17,   -99,   -57,    33,    93,   112,    54,     1,   -54,   -23,    -6,   -15,     6,    81,    39,    13,   -21,     5,    39,   -35,   -83,   -75,   -25,   -48,  -112,   -38,    -8,     7,   -32,   -58,   -34,     8,    31,     7,    62,   -46,    -4,   -45,     6,   -13,    75,    28,    21,   -28,   -44,   -51,   -47,   -26,   -11,   -51,  -107,   -99,   -59,   -46,   -56,   -14,    -6,    86,    71,   -26,   -64,   -75,   -52,    26,  -130,  -125,   -67,    12,    68,   -17,   -39,   -49,   -36,   -84,  -139,   -60,   -70,   -83,   -45,   -74,   -28,   -50,   -19,   -45,   -52,   124,    37,  -178,  -124,   -65,   -33,   -19,  -178,  -105,   -63,   -97,     6,   -21,   -43,   -33,    42,   -61,  -110,  -121,  -102,  -109,    -8,   -59,   -36,   -38,    -2,    -1,     0,   -53,    -3,   -55,   -54,   -68,  -109,    26,   -82,   -11,     4,   -91,    82,     8,   -50,    -4,    76,   -75,  -177,     7,   -42,   -31,    56,   -85,   -22,    15,     6,    -5,   -41,  -160,   -86,    10,   -90,  -118,    26,    36,   -10,    21,   -28,  -152,    -3,   -49,   -17,   -42,    19,   -24,  -127,   -14,   -45,    20,    13,  -102,   -50,     6,     3,    -9,    14,   -92,   -90,    18,   -21,    36,    66,   -63,   -24,    -8,   -46,   -85,   -32,   -50,    17,   -56,    15,    86,   -26,     9,    47,   -21,    58,    10,    13,    14,   -20,    -1,     2,   -53,   -69,  -137,   -40,    29,    32,     5,   113,    51,    29,   -89,   -65,   -98,   -93,   -70,     9,    30,    61,   -13,   -47,     2,    36,    55,     0,     9,    -6,   -16,     7,     0,  -116,  -103,    44,    33,    29,    17,    13,   101,    74,   -64,   -20,   -15,  -149,     3,    31,    37,    80,    11,    76,    38,    -9,   105,     9,    -8,    12,    -5,   -19,   -16,   -77,  -169,    30,     0,    -8,    -9,    54,    61,  -148,  -214,   -67,     9,  -128,    29,   -78,  -127,     5,    10,    65,     6,   -18,   -35,    -6,    11,    11,    -8,    16,   -89,   -26,   -91,  -109,   -45,   -67,   -82,  -120,   -87,  -104,  -137,   -32,     9,   -29,    26,  -104,  -134,  -139,  -157,  -115,    -8,   -15,    10,     4,    20,    -6,     5,     7,     9,    -8,   -16,   -39,   -52,   -55,   -36,   -96,   -78,   -61,   -72,  -127,   -16,   -59,  -103,   -89,   -77,  -104,   -68,   -81,   -14,    -1,    -3,     6,     2),
		    55 => (  -15,    -1,    10,    -6,    -2,    15,     3,    14,   -10,   -16,    13,    -7,     5,   -28,    12,    11,    16,   -15,     4,     0,    20,     9,    18,    -5,    -1,   -12,     6,     7,    -6,    -2,   -16,     2,    -2,     0,    -2,   -25,     6,     0,   -13,   -64,   -35,   -25,   -79,   -99,   -89,  -103,   -73,   -84,  -117,  -114,   -40,   -10,    -4,    11,    -8,     1,   -13,   -14,   -62,   -62,   -29,   -31,   -61,   -58,  -101,  -158,  -142,  -165,  -201,  -255,  -127,    40,    52,    76,    38,   -33,    -8,   -90,   -93,   -21,   -83,   -61,    16,    -9,    10,    12,   -31,    -1,   -26,   -97,  -183,  -118,  -241,    50,    92,   -13,    30,     1,   -62,  -112,   -95,    -4,    56,   116,   -15,    94,     3,   -85,   -46,    52,   157,     0,   -11,   -43,   -79,     1,  -105,   -18,    -6,    21,     2,   -21,    37,    -9,    37,   -52,   -25,   -64,  -103,   -63,    68,   -92,   -84,   -16,   -50,   -43,   156,   105,    24,   -51,    -9,    12,   -80,     0,   -81,   -26,   -65,    12,   -59,     5,    -2,   138,   110,   -36,    44,    88,   -12,   -75,  -182,   -34,   -14,    -2,    16,    77,    -3,    97,    35,   -10,    19,    -1,    -7,  -114,  -116,   -57,     3,    51,    48,   -12,    -2,    97,   136,    17,    16,   -50,   -70,   -89,   -93,   -15,   -37,   -30,    32,   128,   125,   155,   -15,    19,    13,   -65,    15,  -190,  -173,   -74,    55,   126,   110,    94,   100,    39,   -17,    15,    54,    -3,    73,    24,  -104,   -28,    28,     1,    10,    -3,    34,    34,   -40,    69,   -19,   -51,  -146,  -245,  -124,    79,    -4,   -89,   -20,    34,    37,    -9,    -9,    12,    72,    76,   -12,    51,   -85,  -163,   -44,   -44,    15,    -6,   176,    67,  -127,    36,     1,   -16,  -112,  -178,   -68,    71,    39,  -105,    23,   -52,    12,   133,    81,   120,   171,   106,    11,   -47,  -173,  -190,  -190,   -95,    32,    -3,    97,   107,   -67,   -48,    -2,    -8,  -141,  -296,   108,   116,    71,    35,   -52,   -38,    59,   107,   193,   136,   127,   143,     5,  -180,   -93,  -126,  -123,   -75,  -247,  -210,    79,   114,   104,   -63,    13,   -30,   -12,   -65,    30,    63,    47,   -22,   -33,   -43,    -4,    43,    87,    94,    35,   104,    46,   -18,   -59,  -154,   -89,   -70,  -251,  -284,   -13,   -14,    47,    20,   -11,   -15,   -24,   -42,    80,    32,    -3,    13,     1,    -9,     2,   -89,    17,    15,   -16,    20,   -57,   -69,     0,   -36,  -104,   -30,  -183,  -121,  -280,  -118,   109,  -118,     2,    -8,   -51,   -12,    -3,    63,   -47,     3,   -14,   -13,    -2,    42,    13,    15,   -19,    26,   -34,   -94,    -7,    47,    13,    15,   -42,  -148,  -228,  -173,     3,   -81,    20,   -18,   -20,    14,  -117,   -18,   -37,   -24,   -54,   -14,   -12,   -46,    -4,   -69,    17,   -53,    55,   -11,   -50,    17,    51,   -18,     1,   133,     9,  -113,   -69,   -44,     5,     9,   -60,   -41,    17,     0,   -11,   -17,  -143,   -95,    23,   -11,    11,   -48,   -11,     4,   -30,   -16,    10,   -49,   -72,  -146,    -7,   127,    57,  -113,  -108,  -122,     5,   -38,  -138,   121,    13,    43,  -166,  -243,  -116,  -127,   -61,   109,   -14,   -18,   -27,   -76,   -29,   -76,     1,    40,   -43,   -48,   -12,    57,   -40,  -243,  -142,  -136,    -6,   -29,  -213,   214,    46,     5,   -49,  -220,  -151,  -115,   -50,   -12,   -80,   -52,   -57,   -48,    27,    74,    25,    87,     2,    -4,    20,    46,  -135,  -243,  -197,  -200,   -26,    18,  -144,   210,   204,   115,   -13,  -125,  -173,  -243,   -35,  -104,   -63,  -101,    -5,   -12,    48,    59,   -17,   -46,    41,    62,    67,   112,   -13,   -36,  -214,   -67,    -1,   -55,   111,    11,   164,   154,    45,   -82,   -35,  -137,   -58,   -70,   -18,   -16,     1,    55,   -44,    36,   113,    -3,   129,     7,    81,   117,   127,    72,  -132,  -144,   -19,   -57,    87,   -21,    73,    85,    16,     2,     8,   -23,   -84,     2,   -14,    61,   -21,   -41,    61,    89,    12,   -74,    61,   -22,   156,    67,    66,   120,  -115,    -4,   -13,   -20,  -104,  -194,   -13,    72,   -42,   -68,    77,    71,    -3,   -32,   -42,    -8,    37,    97,    89,    45,    88,    83,    22,    91,   -15,   103,    40,   171,    60,   -24,   -24,    -9,  -158,   -65,  -121,  -111,   -65,    14,    21,    42,    49,   -20,    -1,    28,   -25,     3,    30,     1,    23,    80,   -54,    -1,    -3,   177,   184,   221,   142,     3,    10,    13,    29,    36,   -55,   -36,    15,   -25,   -96,     7,   -26,   -14,   -41,    33,    35,   -18,    32,    27,    70,    73,   -29,    34,   -49,   127,   124,   152,   102,    -6,    20,   -13,  -101,   -28,   -80,   -50,   -64,    40,    53,   138,    97,    84,   -23,   -59,  -106,    22,   -29,    98,    79,   103,    38,   -55,    30,    -2,   145,   -96,   -55,     5,    19,     3,     1,    74,  -151,  -189,   -66,   -30,    27,   -66,   -95,   -94,     5,   -53,  -118,     1,   108,   149,   135,    95,    22,   106,   168,   143,   142,   -53,   -19,   -11,    19,    14,   -19,   -42,   -67,  -144,  -187,  -173,   -65,   -14,    40,    31,     0,   -33,  -156,    51,   -29,    45,    41,   158,    43,    -5,   -39,   -79,   -45,    15,    16,    11,    -8,    19,    18,    -5,   -35,   -33,   -13,   -37,   -39,   -44,    18,    19,    25,    12,  -198,  -149,   -44,   -66,   -46,   -91,  -111,  -126,   -70,   -13,    12,    15,     8,     4),
		    56 => (   -1,    -7,    -1,    -9,    10,   -10,    16,    -6,   -12,     5,    -1,   -20,    31,    43,   -12,    19,   -16,    17,     8,     2,    19,     7,     9,     4,    -1,     4,    10,    -9,    15,     4,    -2,   -18,   -19,   -17,    43,    49,    93,    57,    43,    33,    14,    67,    -9,   -28,   -21,   -14,     2,    18,   115,    57,    38,     8,    -6,    -7,    -1,    -5,    -1,    -8,    -8,    -6,    61,     1,    33,   103,    88,    79,    50,   -31,   -45,   -51,   -45,   -20,     2,   -13,   -12,    52,    64,    85,    66,   107,    42,    40,   -14,   -13,   -13,   -16,   -90,   -91,   -19,    68,    61,    46,    33,    55,   -15,   -71,   -93,  -183,   -82,   -44,   -11,   -78,    36,   111,    64,    45,    23,   103,    73,    14,    -8,     6,    19,     2,  -107,  -115,    81,   110,    69,    14,   -39,    35,    11,   -99,  -127,  -188,  -122,   -10,   -28,   -54,  -122,     7,     9,   -37,   -80,     8,    80,    67,   125,   135,   -15,    19,   -58,  -104,   164,    92,    36,    21,    26,    10,    -3,   -49,   -73,  -138,   -53,    45,   -25,    21,   -51,   -56,   -60,   -24,   -45,    25,    50,    61,   137,    94,    -7,     0,    31,   -23,   122,    35,    66,    23,   135,    56,   -59,  -130,  -136,  -147,   -33,   -40,  -113,   -49,    -5,  -107,   -65,    -8,   -20,    -5,    18,   -77,    30,   160,     2,    -6,    10,   -37,   130,    52,   -23,    73,    59,    77,   -41,  -115,  -156,   -85,     0,  -107,  -134,    -6,    -7,   -18,   -20,   -63,   -70,   -86,   -84,   -33,    57,   138,    -1,     8,    10,   -43,    97,    30,   -24,    54,    13,    -9,   -89,  -154,  -171,     4,    13,  -121,   -21,    53,    27,    48,    54,    18,   -68,   -23,   -20,   -46,    61,   -84,   -10,   -11,   -22,   -85,    61,    22,   -32,    50,   -17,   -76,  -165,  -185,  -163,   -56,   -23,   -48,    36,    93,    12,    40,    68,     7,   -28,    11,   -17,   -82,   -27,   -27,    -8,   -13,   -31,   -80,    95,    63,    36,   114,    12,   -81,  -129,  -156,  -124,   -26,   -16,    18,    17,    79,   -69,   -38,   -43,    32,     5,    12,   -38,   -32,     0,   -15,     1,     9,    16,   -23,    76,    73,    51,    26,    -8,   -61,   -99,  -121,   -72,   -10,    16,   -11,   -35,  -139,   -93,   -25,   -60,     1,    35,    49,    13,     8,   -30,   -45,   -19,     6,   -21,   -41,    48,   118,    -6,    26,    -9,   -64,   -97,  -134,   -39,   140,    25,    18,    21,   -52,   -48,   -75,   -34,    40,    78,    65,    53,   -11,   -15,   -85,    16,    19,   -13,   -37,    22,    22,   -20,     5,    33,   -50,   -61,  -147,     5,    75,   -29,   -74,   -10,     7,   -55,   -53,   -34,    34,    32,    61,    51,    -4,   -12,   -19,   -11,    -4,     9,   -55,    12,    25,   -25,    30,     0,   -11,   -81,   -53,    68,    88,  -128,   -90,    -3,    13,   -19,   -18,   -73,   -24,     9,    45,    36,    -7,   -27,   -32,   -18,     1,     8,   -32,    50,    18,   -33,   -13,    -7,    -8,   -70,    -3,    -1,    45,   -52,   -20,     9,   -24,   -10,   -75,   -78,     0,    37,    78,    29,   -15,    15,  -125,    12,    10,   -34,   -14,    66,     9,   -57,   -45,   -49,   -35,   -39,   -24,    49,     2,    27,   100,     9,    11,    49,   -82,   -47,    -8,    48,    40,   -15,    22,    -1,   -58,     6,    11,    -4,    51,     0,    15,   -28,   -46,   -37,     6,    31,     7,   -34,    52,     3,    20,   109,     2,    40,   -16,   -72,    -7,   -10,    46,     1,    -1,   -21,   -52,    10,     2,   -11,    15,   -35,    20,   -77,   -65,   -67,   -13,    -2,    48,   -43,    18,   -43,    44,    26,    14,    78,    28,   -12,   -33,    32,    51,    -5,   -16,    -2,   -44,   -18,   -16,   -17,    62,     9,   -11,   -81,   -99,   -84,    -6,     7,    -6,   -24,     0,    22,    55,     7,    16,    77,    81,    54,    23,    -4,   -63,   -35,    22,   -86,    -9,     4,   -26,   -13,   -48,   -41,   -57,   -23,  -112,  -100,   -38,    16,   -36,   -35,    27,    22,    59,    35,    81,    71,   -52,     2,   -47,  -114,   -57,   -42,    40,   -30,    -1,   -17,    14,   -14,   -46,   -14,   -56,    -5,   -57,   -46,    15,     1,    -4,     3,    63,    27,    35,    25,   -46,   -64,   -35,     4,   -29,   -68,   -54,   -52,   -41,   -21,     8,    -7,   -17,    -4,   -54,     1,   -34,   -80,   -46,    13,    -2,   -37,   -54,    -6,    49,   -37,    23,   -22,   -39,  -108,     9,    -6,   -58,   -84,   -94,  -100,   -34,     1,    17,     4,    15,     5,   -30,   -39,     1,   -30,   -55,   -37,   -42,   -20,   -56,    -3,   -82,   -50,    29,   -55,  -114,   -54,   -46,   -37,   -10,   -56,   -61,   -74,    -4,   -25,   -13,    -6,   -17,   -20,   -19,   -14,   -25,     9,    -6,   -27,   -12,   -59,   -29,   -12,   -20,   -39,   -17,   -10,   -21,   -41,   -90,   -52,   -25,   -13,   -16,    -8,     7,     9,   -18,   -14,     4,   -20,    15,   -21,   -25,   -48,   -31,   -20,   -32,     3,   -22,   -32,   -24,     5,    -2,   -10,     6,     3,   -19,   -71,   -28,    -1,    25,   -16,    -8,    -7,    -4,   -19,    15,     7,    15,   -18,    -2,    -8,    -4,   -19,    10,   -21,     0,    -6,    -4,     9,    -4,    12,   -18,   -10,     5,   -39,   -21,   -12,     5,    -4,     2,     0,    -8,   -20,   -10,    17,   -20,     1,    -1,    -8,   -15,   -19,    -9,   -24,   -18,    -9,   -19,    -1,   -14,    -4,   -14,   -14,    11,    13,   -19,    -1,     8,    -6,    16,   -14,     5),
		    57 => (   -7,   -18,    14,   -10,   -15,    13,   -14,   -16,   -10,     6,    -7,    -4,     9,   -14,   -12,   -16,    18,    -2,     0,    -8,     2,    -5,    -7,    -1,    12,    12,     1,    19,     3,     4,     3,    -9,    12,   -14,    16,     8,   -13,    -9,    -9,   -77,   -87,   -76,   -50,  -168,  -199,  -211,   -45,     6,   -19,     1,   -14,     0,   -14,     4,   -16,     1,   -12,   -10,    -9,   -19,    12,    11,   -38,   -39,  -122,  -123,  -181,  -163,   -98,   -61,   -46,  -107,   -84,   -47,   -59,    -3,  -100,   -88,   -78,   -68,   -63,   -29,     6,     7,    -4,    -8,   -11,   -46,   -39,  -134,  -212,  -210,  -189,  -125,  -189,  -276,  -277,  -196,  -180,  -167,  -117,   -80,   -73,  -130,   -63,  -102,  -301,  -197,   -93,   -48,     3,   -18,     8,    10,   -14,   -81,   -90,  -151,  -205,  -284,  -311,  -373,  -399,   -63,   -17,   -31,   -53,   -92,  -213,  -293,  -241,  -161,  -118,  -108,  -183,  -247,  -249,  -141,   -31,    14,    19,    14,     7,  -107,  -154,   -62,  -121,   -82,   -21,    52,   -49,    47,    80,    71,     1,   -23,   -48,  -147,  -198,  -256,  -263,  -166,  -168,  -365,  -270,  -236,   -21,     7,     5,    -9,   -57,   -49,   -37,    50,    38,    34,     8,    36,   109,   103,     6,    19,   -90,   -39,    39,   -57,   -15,  -106,  -138,   -70,  -114,  -126,  -161,  -168,  -104,   -76,    12,    66,   -56,    16,   -18,   143,    88,    96,    74,    86,   110,    -4,    40,    66,    58,    11,    53,    71,    94,    50,   -34,   -20,   -25,   -48,  -121,  -258,  -161,  -101,   -71,    44,   -12,    72,     0,   122,     8,    35,    20,   -46,    62,    72,   -88,  -110,   -73,    44,    70,    45,    73,    58,    56,    49,   -30,    -5,  -117,  -147,  -153,   -70,   -15,    50,    57,    50,    72,     9,   -26,   -13,    -6,   -27,    14,    54,   -18,   -39,   -96,     7,    17,    95,    84,    22,    -2,    79,    26,    65,  -114,   -24,   145,   201,   -13,    92,   -14,   -48,    46,  -101,    14,   -55,    18,    26,     3,    42,   -70,   -94,   -14,    12,    74,    75,   100,    62,    56,   -22,    66,   -22,   -17,    77,   129,   173,    -8,    -2,     2,   -42,    61,    50,   -71,   -44,   -13,    61,    25,   -72,   -29,    78,   -22,    -5,    68,    36,    85,    53,   -55,    15,    89,    71,   -31,  -124,    -8,   111,   -11,    51,    76,     8,    82,   115,     9,   -74,    74,   -26,   -83,   -29,   -28,   -26,   -24,    89,    67,    81,    35,     7,   -11,    23,     6,    43,    14,    66,   115,   181,     2,    29,   110,     0,    82,    97,   -28,   -42,    30,     2,    -5,   -12,   -52,     4,   -54,    26,    12,    13,    -8,    14,   -38,   -19,    93,    32,    89,    98,   -19,   -51,    -3,    44,    39,    15,     3,    71,   -73,    46,    40,   -21,    -3,   -22,    12,   -48,   -35,     4,   -43,    53,    -4,    43,   -29,   -38,    24,   -39,   -26,  -194,  -177,   -28,    17,     0,   -19,    -9,   -41,   -62,     3,    23,    19,    44,    53,    25,   -24,     8,    47,    71,   -41,     7,    37,    42,   -15,    -5,   -57,  -118,  -166,  -198,   -22,  -131,     7,     1,   -26,   -93,    22,    51,   -53,   -64,   -37,    32,    40,     5,    39,   108,    66,   156,    35,    20,     8,   -46,   -71,   -46,   -16,   -38,   -73,  -179,  -134,  -131,   -16,   -21,   -70,  -136,    37,    20,   -12,   -73,   -64,  -136,   -37,   -52,    78,    93,    70,    64,   -13,   -45,   -61,   -54,   -36,   -28,    -1,    -9,    83,  -106,   -57,  -140,    30,    12,    39,  -228,     9,   -23,   -89,   -70,   -64,   -71,   -58,    -7,    16,    25,    39,   -42,  -125,     8,    -4,   -56,    94,    87,    26,    91,    27,  -164,    18,   -93,    18,    24,   -12,   -87,   -64,   -13,   -43,  -105,    -4,   -58,   -76,   -17,    43,    63,   -18,  -134,   -11,     4,   -16,   -14,    31,   109,   -37,   -86,    64,  -173,  -152,   -51,    -9,   -10,   -45,   -49,  -180,  -135,  -106,   -72,  -136,   -50,  -129,  -122,   -54,    34,    16,   -70,   -18,     9,  -146,   -14,    15,    27,   -66,  -169,   -69,  -149,  -129,    13,   -13,     4,   -69,  -122,  -167,   -19,   -42,   -42,   -52,  -120,   -33,   -46,   -37,    31,   -44,   -25,    20,     1,  -112,   -54,   -65,    84,   -64,  -148,  -213,   -56,   -39,     1,   -29,   -29,   -92,  -115,    -6,    19,    -2,   -46,    49,    -6,   -46,   -18,    21,   -53,    -5,    10,    90,   -11,   -24,    30,    83,    -8,   -93,  -381,  -204,   -19,   -63,     0,     7,   -19,   -73,  -136,    26,    34,    30,    23,    86,    45,     1,    36,   108,    64,   129,    20,    66,    60,     4,     0,    61,   -14,   -93,  -333,  -179,   -93,  -150,    -9,   -15,    11,    57,   -45,   130,   128,   127,   118,   112,     6,    60,    86,    98,   203,   178,    11,   115,    82,    18,    70,    64,    39,   -26,  -231,  -125,  -131,   -99,    14,    -2,   -12,   -15,    51,    56,    74,    62,    73,    65,    85,   149,   141,   108,    91,    38,   -53,   175,    69,    48,    51,    -3,    93,   106,   -33,   -31,  -102,   -72,    13,    -4,    11,    15,   -68,   -55,   -97,     7,    71,    74,   110,   116,   121,   112,   -96,  -173,   -18,    71,    12,    31,   109,    59,    90,   113,    38,   -50,   -12,   -15,    -4,   -10,    11,   -12,    -5,    39,    43,   -28,   -47,    -6,    52,    89,    18,    -9,  -132,   -30,    34,   -52,    61,    37,    44,    29,    93,    45,   121,     9,    -1,   -16,     6),
		    58 => (    9,    -7,    -4,     3,    11,   -16,   -12,    20,    -7,     8,   -14,   -19,    -8,   -17,     2,     9,     5,   -16,    15,    -6,    12,     1,    20,    -6,     2,     2,    -1,    19,     5,     4,   -12,   -17,   -14,    12,     3,     6,    -6,     6,    18,   -29,   -55,   -34,   -40,   -22,   -60,   -59,   -66,   -27,    11,    13,   -11,    20,     4,    16,    -6,    10,   -14,   -18,   -12,    -4,    -8,   -17,   -33,   -46,  -122,  -118,  -170,   -85,   -10,   -11,   -67,   -66,  -101,    23,    13,   -55,   -54,   -55,   -53,   -21,   -20,   -17,    -4,   -10,    -4,    -4,   -32,   -44,   -29,   -66,  -128,  -238,    23,    59,    57,   -10,   -63,   -79,   -55,    67,   -74,   -97,    17,   -61,   -48,   -56,    56,   109,     3,   -40,   -62,    17,    -7,   -59,   -53,  -147,  -124,  -140,   -78,    82,   180,   152,   119,    61,   -20,   -10,    53,    60,    50,   126,   -24,   -78,  -105,  -127,   -60,  -108,  -139,    14,    72,   -28,     6,    16,  -104,  -123,  -102,  -148,   -14,   202,    74,    86,    50,   103,   112,    50,    11,    31,    54,   114,    -6,   120,    -8,    18,    46,   -37,   -49,   -35,  -105,   -42,     8,   -19,  -160,  -133,  -141,   -72,   -49,    94,   -40,     9,    78,    14,   -11,    31,   -14,    37,    -8,   -28,    31,    34,    78,     5,   -13,    57,   -40,   -67,   -33,   -25,     8,  -108,  -131,  -156,  -130,   -98,    -2,    12,   -18,    -7,   -18,    82,    -2,    25,   -77,    56,    27,   -15,   -25,    22,   -48,   -21,   -38,   149,    89,  -149,  -100,    48,    36,   -74,  -115,    15,   -14,   -11,   -18,    80,    34,    16,    21,     5,   -16,    17,    -8,   -16,   -23,    -8,    55,   133,   -53,   111,    86,   141,   152,   -89,   129,   142,    11,   -37,  -149,    34,    79,   -44,     4,    70,    37,    -1,   -52,     2,   -13,     1,    44,   -23,   -29,    40,    17,   -15,    91,    84,    90,    63,    29,   -41,   128,  -163,   -12,   -13,  -179,  -121,   164,    49,   -58,    56,    58,    29,    78,    29,    30,   -21,    78,  -131,  -101,    10,   -20,     3,    26,    96,    43,    91,    67,  -134,    52,   -64,    12,   -20,   -83,    -2,   151,   130,    31,    90,    27,     9,    33,    -1,   -41,   -40,    28,  -115,  -104,   -77,     9,    -3,    41,    60,    69,    82,   101,    33,   152,   -32,   -10,    10,  -123,    32,   148,   261,     7,    12,    91,    40,    -4,   -53,   -83,   -80,   -11,   -59,     5,    -7,   -63,   -40,    54,    58,   136,    15,    60,   -58,    78,  -139,    18,   -13,   -75,    -8,    52,   145,    48,    26,    63,     9,    -9,   -21,   -20,   -32,   -19,    23,     3,  -105,   -51,   -40,    68,    29,   117,     7,   -78,   -84,    61,    21,     3,   -32,   -32,   -94,  -140,    19,    91,  -125,    70,  -163,  -112,   -32,   -64,   -73,     6,    14,   -43,  -112,     3,   -95,  -133,    40,    -6,   -40,  -109,   -16,   -69,   -46,    12,    12,   -56,    49,  -235,   -57,   -77,   -90,    39,   -95,   -32,   -32,  -113,    13,    41,   -62,   -48,    12,   -87,   -38,   -66,  -105,   -33,  -130,  -168,   -39,  -181,  -107,    13,   -22,   -34,    65,  -223,   -94,  -115,  -185,   -99,    -9,  -118,   -80,   -14,    61,    -6,   -34,   -86,  -155,   -77,    -9,   -83,  -121,   -65,   -41,   -63,   -63,  -205,  -106,     6,   -22,   -48,  -109,   -62,  -113,  -126,  -120,   -17,   -79,   -77,  -127,   -32,   -40,   -63,  -119,   -57,   -50,   -54,   -27,    11,   -30,   -32,   -18,   -22,  -197,   -95,  -152,   -24,   -27,   -73,  -202,     2,  -113,     3,    34,    16,   -16,   -39,   -53,    22,    -7,   -73,  -214,    -8,    19,     4,    38,   -18,   -37,     8,    -2,     7,  -183,   -79,   -99,    11,     8,  -151,  -187,   -42,  -113,   -70,    33,   120,    31,    22,   -45,   -79,   -71,  -129,   -87,   -25,    91,     9,    41,    45,   -65,    28,    93,   122,  -240,  -179,  -118,     7,     4,   -57,  -155,  -121,    25,    60,    16,   106,   -41,   109,    -5,    54,     3,   -81,   -29,    94,    65,    16,     3,    78,    83,    76,   196,    45,  -293,  -183,     8,   -49,   -79,   -71,   -85,   -98,    21,   132,    17,    83,   134,    59,    52,    31,    72,    62,   158,    -6,   107,  -113,    50,     9,    12,   148,   128,   -52,  -222,  -138,    -1,   -53,   -67,   -37,   -70,    58,   133,    79,   121,   106,   106,   147,   145,    66,   109,   183,   187,    30,    23,    44,   -42,     1,     4,   125,    72,   -70,   -12,  -139,   -10,   -17,    12,   -21,   -35,   128,   -12,    48,   -29,    57,    60,    15,    21,   121,   122,   119,   133,   118,   101,   119,   168,    40,   -47,   172,    87,   -42,   -16,  -142,     1,    16,     4,   -56,   -86,   -51,   -54,   -30,   -43,    47,    85,    38,    16,   111,    35,    50,    81,   173,   -19,   -10,   -22,    17,   -86,    22,    29,   -81,  -192,  -100,   -16,    18,    -4,   -60,     6,  -238,  -190,   -12,   -16,   -79,  -141,   -75,   -79,   -48,   -39,    53,    66,   -22,   -45,    37,   -19,  -135,  -123,  -129,   -66,   -77,   -48,   -29,     2,     5,     8,     2,   -54,  -108,  -188,  -175,   -42,    31,    11,   -92,   -49,    44,    29,  -153,  -324,  -149,   -88,   -74,  -239,  -205,   -97,  -112,   -41,   -10,     7,     0,   -13,     0,     3,    -9,    11,   -47,   -40,   -51,   -32,   -66,   -59,   -14,   -19,   -80,  -131,  -154,  -123,   -65,  -102,   -52,   -57,     1,     0,   -41,     0,    -5,   -17,     6,    -6),
		    59 => (   15,   -10,    18,    -5,   -16,    14,   -10,   -13,    18,    -2,    16,   -13,     7,    10,    -7,   -18,   -12,   -20,   -12,    -7,    19,    -8,   -19,    18,    18,    14,    11,   -13,     7,    14,     3,   -16,   -15,    14,     5,     0,   -20,    -6,     2,   -23,   -34,   -44,    17,   -26,   -11,   -33,    -3,    15,    10,    16,     7,   -15,   -12,   -17,   -18,    15,    -8,   -15,     7,    15,   -19,    12,   -17,   -13,   -32,   -21,    -9,   -33,   -15,   -18,   -60,   -18,    14,   -18,    10,   -14,   -16,    10,    -8,     4,   -11,   -14,    -4,    12,    -5,    -9,    12,   -15,   -28,   -39,   -32,    -4,   -50,   -79,   -24,   -62,   -21,   -84,   -58,   -65,   -16,    12,    33,     4,   -80,   -60,   -25,   -23,     5,   -24,     5,    20,    17,    -4,    12,    -4,    -6,   -21,   -80,   -27,   -24,    -3,   -40,     4,  -113,  -152,  -127,  -104,   -87,   -86,   -42,  -111,  -123,     0,   -16,     2,   -14,   -85,   -70,   -19,   -17,    -2,    -1,    -6,   -20,     8,   -17,   -51,  -159,   -62,   -75,     7,    23,    -1,    26,    -3,   -37,  -123,  -154,   -86,   -17,   -25,     2,    -7,     8,   -78,   -39,    11,    -8,    10,   -23,   -14,   -57,   -87,   -75,  -119,   -27,    53,    11,    92,    91,    74,    -9,   -43,    58,   -26,  -199,  -185,   -88,     3,     7,   -14,     0,     3,   -12,   -54,   -19,    -1,   -22,    13,   -40,   -95,  -148,  -113,    -9,   -70,    24,    82,     9,    41,   -45,  -123,   -95,  -102,  -214,  -276,   -96,    18,    -5,     3,   -35,    -1,   -18,   -45,   -39,   -22,   -40,    50,    15,  -102,    86,   -23,    73,     6,    -6,    17,   -26,    14,   -23,   -92,  -102,   -56,    27,   -67,  -148,   -26,   -26,   -36,   -45,   -13,    -9,    -2,   -13,   -71,   -65,    28,    -6,   -64,    65,    61,    27,    51,    83,   -43,   -49,    22,    14,   -80,  -124,    55,    52,   -51,   -95,   -77,   -94,   -38,   -72,   -95,   -44,   -45,    -6,   -23,   -32,    30,   -20,  -102,    86,    47,    36,    15,     9,  -170,  -147,    26,    98,   -19,    57,    -4,    -4,   -50,   -87,   -97,  -109,   -71,   -62,   -78,   -13,   -73,   -12,  -108,   -46,    52,   -47,  -114,    39,    92,    69,    18,   -33,   -16,    60,   206,    -6,   -18,   -18,    72,   -29,   -12,  -146,  -162,  -104,   -98,   -34,   -69,     3,   -66,    16,   -41,   -45,    68,   -36,    36,    35,   -16,    -6,    80,    38,    15,    66,   137,   -53,  -110,   -24,    58,     0,    -6,   -56,   -89,  -143,  -108,   -64,   -54,   -61,   -73,    13,   -44,   -34,   -54,   -70,     6,   174,    24,   -82,    13,    29,   -37,    -1,   -26,   -37,   -24,    -8,   -14,   -62,    38,   -64,   -85,   -81,   -78,   -37,   -43,   -53,    -2,   -17,   -10,   -32,   -38,   -50,   -45,   112,    12,   -44,   -34,    88,    -3,   -63,   -39,    29,    33,   -24,     3,     4,    -2,   -59,  -108,  -115,  -116,   -52,   -83,    -6,    -6,   -21,    -5,   -33,   -42,    56,   -77,   -74,    14,   -22,   -57,    43,    16,   -41,  -117,   -51,    29,    33,    -4,   -29,   -28,  -179,  -161,  -111,  -103,   -30,   -20,     0,   -50,   -14,    -1,   -56,    -9,    -4,   -46,  -172,   -17,    31,   -65,    22,   190,    67,    26,    11,   -81,   -67,   -68,   -24,   -70,  -234,   -88,   -49,   -37,   -32,   -23,     5,   -82,    -8,   -10,   -71,     7,    -5,   -63,  -135,  -161,   -16,  -121,   -42,    51,    91,    59,    12,    10,   -93,   -99,   -64,   -53,  -153,   -98,   -35,   -58,   -88,    67,   -61,   -40,   -20,     1,   -65,    -5,     6,    -1,   -42,  -100,  -130,  -123,  -129,   -53,    69,   -35,   -30,   -42,   -25,    -3,   -91,   -32,   -64,  -110,     2,   -38,  -102,   -14,   -51,   -41,   -19,    -6,   -51,   -13,     0,   -31,   -17,    -3,   -27,   -22,  -106,  -166,  -155,  -147,  -111,    61,    32,    10,   -60,   -61,   -99,  -112,   -56,     0,   -71,    74,   -51,   -43,    -9,   -25,    -2,   -31,    -7,    -3,    -6,   -79,    -5,   -78,   -87,  -145,  -189,  -114,    -7,    15,   -15,   -25,   -51,   -58,   -45,   -36,   -43,   -50,    15,    48,   -66,     3,    13,   -19,     9,   -29,   -16,    57,   -24,   -27,   -11,    12,    18,   -21,   -49,   -18,    18,   -62,   -12,     2,    -2,  -106,   -39,   -68,   -36,   -18,    38,    78,   -87,   -20,    -4,   -12,   -26,    52,     0,    19,    34,    32,    38,    60,   -28,    21,    59,    27,    23,    39,   -12,    41,   -25,   -96,   -65,  -109,   -22,     1,    27,   -21,    -5,   -12,    16,    13,   -43,    25,   -18,   -16,    42,    -8,    32,   -27,    19,   -23,     1,    -7,   -12,    59,     4,    37,    55,   -39,   -44,   -52,   -12,    38,    22,    20,   -43,     1,    -4,    -4,    -6,    -8,   -21,    14,    -1,   -55,     6,   -41,    48,   -49,  -135,  -103,   -32,    27,    50,    35,    38,    48,    38,     8,   -12,    29,    20,    30,   -11,     3,    -4,    -6,    34,    -9,   -12,     7,    10,   -31,   -24,    29,   -64,   -83,   -53,    21,  -101,   -80,    16,    76,    22,   -82,  -100,   -87,   -76,   -37,   -28,    29,     6,    14,     9,   -11,    14,    34,     4,    -1,     4,     9,    21,    53,   -40,   -89,    79,     7,    82,    45,    26,   181,    68,   -83,    16,     7,   -17,    27,    26,    14,    -1,   -19,   -19,   -12,     1,   -13,   -14,   -18,    35,    46,    23,   -58,   -27,    19,    -7,   -60,   -76,   146,   136,   -13,   -31,    67,    28,   -55,   -43,   -12,    -6,    -4,    17,     5),
		    60 => (    6,     1,    11,    14,    15,    -2,    16,    14,    -4,     3,     7,    19,     2,    -3,   -18,    11,    -6,   -17,   -16,   -17,    13,    12,     1,   -17,     0,     3,    -5,    19,    -1,    -8,    18,     5,    -1,     9,    -7,   -43,   -37,   -49,   -88,   -39,    13,    24,  -115,   111,   136,   139,     6,   -19,   -28,   -24,    12,    -3,    13,    11,    -1,    -1,    -3,   -14,    17,   117,   142,   -40,   -65,    21,   -28,   -78,  -127,  -109,  -137,  -263,  -136,   -64,    -9,  -100,   -67,   -70,   -75,   -65,  -185,   -71,   -89,   -17,     8,    18,    13,   -11,    15,   125,    42,  -119,  -140,  -121,  -117,   -94,   -65,  -148,  -207,   -98,  -114,  -124,    48,    51,     2,   -96,   -97,  -142,  -202,  -101,   -74,   -83,  -148,    16,    -1,    -1,   -12,   -35,   -48,  -245,   -89,  -104,    10,   106,   -12,    19,  -118,     0,   -45,    43,   108,    52,    -8,     3,   -89,   -89,   -35,   -53,  -165,  -279,  -114,     9,    -6,   -20,   -62,   -40,   -57,  -124,    54,   -22,    25,   154,    97,    83,    19,    12,    67,    61,    62,    67,    62,     3,    -6,   -16,   -69,   -49,  -155,  -242,   -56,   -30,     9,     5,   -87,    -8,  -161,    44,    98,    94,    85,    61,   105,    50,    12,     7,    54,   -56,    22,   -20,   -78,    27,   -17,   -95,    -4,  -185,  -105,  -280,   -80,   -27,    -3,   -41,   -76,   -87,   -93,    -5,    86,    86,   -43,    44,   -27,    17,    26,    33,   -89,  -100,   -43,   -23,   -33,   -87,   -27,   -81,   -19,    -5,   -98,   -53,  -145,    25,   182,  -114,    -7,  -123,  -114,     8,    11,   -91,    18,    31,   -45,   -88,     7,   -26,  -148,   -12,   -32,    72,   -13,   -43,   -50,    20,    -1,    69,  -115,  -267,  -139,   -32,   -22,   -33,    67,    -4,   -28,    30,   -92,   -48,   -19,    41,   -36,    33,    74,    28,    31,    69,    49,    64,    32,    42,    33,   -28,    -2,    68,   -28,  -162,   -43,   -30,   -28,   -24,    85,    33,    13,   -58,   -24,   -57,    15,    57,   -17,   -26,    -4,    60,   182,   135,   124,   150,   -24,    55,    36,   -51,    28,    70,    -4,   -96,  -120,     1,   -13,   195,  -118,   -16,   -35,  -114,   -41,   -60,   -77,   -34,   -55,   -12,    49,   218,    82,    99,   241,   186,   161,    97,    77,    38,    38,    46,   117,  -115,  -122,   -11,   -14,     6,  -121,   -41,    63,  -117,  -105,  -123,   -99,   -22,   -44,    11,   116,   166,   114,   137,    96,    89,    93,    62,   -46,     5,    -8,    31,    60,   -57,   -97,   -64,     4,    17,     1,   -51,    84,   -17,    10,   -69,   -22,   -79,   -60,    35,    46,    14,    -6,    21,     3,   -38,   -20,   -32,   -42,    30,    19,    95,    34,    52,  -169,   -60,   -16,     0,   -21,  -157,   -58,   -29,   -72,   -22,    -6,   -47,   -50,     5,   -46,   -30,  -153,  -176,  -177,   -76,    44,   -30,    67,   142,   145,    81,   135,   115,  -145,   -17,   -13,    13,   -99,  -143,   -30,   -69,   -90,    39,    -5,  -106,   -95,   -72,  -111,  -108,  -238,  -136,   -94,   -27,   -55,    -8,    85,    60,    16,    61,   101,   125,  -154,  -135,   -19,     2,   -58,   -69,    54,   -36,  -102,    24,   -21,   -55,     3,   -51,   -90,  -130,  -135,   -18,  -111,   -98,   -35,    59,    52,   -32,   -51,   -89,   -15,   -44,  -219,   -49,     6,   -12,   -77,     5,    24,    16,   -62,    40,   -19,    24,    47,    73,    30,    81,   -52,   -52,   -83,   -19,   -18,    52,   -15,  -129,   -31,   -45,   -25,  -140,  -138,    38,   -10,    -4,   -65,   -46,    74,    67,    50,   -31,    20,    79,    90,    37,    12,   -51,  -104,   -35,   -36,    27,    22,    20,   -96,   -75,   -45,    49,  -121,  -132,  -108,   -76,    14,    30,   -22,   -41,     2,   107,    69,   119,    90,    24,     1,    19,    94,   -41,   -60,    -2,    -7,    12,    13,    98,   -47,   -71,   -21,    48,    -6,  -218,   -29,   -21,     4,    33,   -94,   -72,   117,    75,    57,    94,    50,   142,     0,    44,   136,    39,     9,    50,     1,    36,    -9,    19,   -87,  -108,   -51,   -31,   -75,  -254,    20,     7,    13,   -18,   -97,   -56,    10,   -15,   101,   141,   114,    84,    57,    17,    79,     8,   -24,    53,    33,     1,    33,    27,   -39,   -78,   -13,    15,  -128,  -123,   248,    -2,   -13,    -9,   -52,   -56,  -168,   -93,   -20,   134,   106,    16,   144,    67,   -17,   -46,    35,    91,    55,    42,   -36,   -31,   -98,   -99,   -41,    -7,   -87,   -52,   151,    30,     6,    15,   -49,  -113,   -38,  -106,   -87,   -12,    96,    78,    56,   -70,    74,   -22,    19,    43,    37,   101,   -22,  -108,  -171,  -115,  -143,   -46,   -97,  -132,  -128,   -20,    20,   -14,   -36,   -59,    34,    63,  -110,   -65,   -60,   -30,   -56,  -182,  -117,  -109,  -103,    59,   -21,    -6,   -66,  -155,   -89,  -161,  -135,  -100,   -85,   -44,   -11,     2,    11,    11,   -17,   -37,  -157,   -98,  -173,  -259,  -144,  -151,  -165,   -97,  -150,   -89,  -104,  -131,  -288,  -248,  -250,  -281,  -196,  -224,  -159,   -71,   -14,    -5,    18,    18,    -5,    -1,    -9,     3,   -51,  -158,  -219,  -106,   -84,  -151,  -108,  -122,   -80,   -94,  -122,  -195,  -162,  -146,  -145,  -177,  -156,  -183,  -114,   -74,   -43,    -8,   -10,     2,    -2,     2,     0,     3,     0,     2,   -10,   -27,   -48,   -88,     5,    -6,     1,  -116,   -40,   -20,    -2,    13,   -66,   -60,   -46,   -88,   -43,   -67,     5,    11,   -16,    20),
		    61 => (  -10,   -13,    11,    -4,   -18,    12,   -16,    11,     1,    -6,   -18,     3,     5,    10,   -15,    -2,   -18,   -17,    -7,    13,   -13,    -1,    -5,   -15,     3,    19,    -9,    -8,    19,     0,     2,     1,     1,     9,    -2,     3,     3,     9,    -5,   -10,   -32,   -33,    27,     7,   -30,   -22,     1,    17,    16,   -14,    -1,     7,    17,     6,    10,    17,     1,    14,    10,     6,   -11,   -12,   -10,    15,   -11,   -16,    -4,    -2,   -74,   -77,   -74,  -157,  -158,   -67,   -46,    -8,    43,   -50,   -37,   -13,   -43,   -40,    11,    -8,     6,     4,   162,   108,    18,   -29,     6,    62,    26,    17,   -25,   -15,  -125,  -315,  -242,  -188,  -127,  -115,   -74,     1,    -9,   -20,   182,    33,   -10,   -49,    -6,    20,    20,   -17,   136,   113,    49,   -42,   -74,   -46,  -121,   -57,  -102,  -118,  -198,  -217,    99,    49,    76,    54,    46,    41,    10,    47,    49,   -60,  -102,  -123,  -106,   -88,    15,   -18,   104,   158,    95,    27,   -34,   -57,  -238,  -144,  -223,  -212,  -209,  -123,     5,    48,   -30,   -57,  -137,   -71,   -30,    38,    87,    -5,   -80,  -133,  -117,  -112,   -10,    -5,   -83,    69,   136,   -68,    96,   146,   -91,  -220,  -247,  -236,  -120,   -45,    -9,   -46,   -28,    13,   -53,   -31,    49,     1,     9,   -25,  -105,  -104,   -66,   -59,   -19,  -115,  -142,   -25,   -92,   104,   110,   136,  -165,  -162,  -360,  -205,  -110,   -49,    -7,     7,    56,    46,    -2,    73,    86,    15,   -72,   -45,  -121,   -86,   -72,   -51,    -1,  -110,  -117,    42,   -90,    74,    96,    31,  -102,  -121,  -152,  -176,  -201,   -98,    -9,    57,    51,    47,    22,    45,    38,    13,   -50,   -91,  -166,   -67,  -140,   -20,    12,   -11,  -106,    22,   -51,   -70,    85,   125,    71,    29,   -33,  -201,   -58,  -151,   -12,    94,   152,    40,    55,    10,   -17,   -59,   -57,   -45,  -105,   -33,    -9,   -38,   -16,    48,  -117,   -40,   -55,  -106,    -5,    97,   -36,   -23,    63,   -19,   -66,  -128,    -8,    33,    58,    42,   -29,   -55,  -144,  -191,     6,   -18,   -90,    -4,     0,   120,     9,    10,   -22,    56,    -7,    93,    64,  -134,  -180,   -67,    43,   -46,  -184,     5,    20,    45,    39,     2,   -64,  -166,   -60,   -36,     3,   -38,   -23,    -1,     6,    96,    -1,    11,   -50,    92,   -25,   120,   111,   -42,   -69,    13,   -18,   -68,   -54,    42,    78,    19,    40,    53,   -97,  -133,   -41,    97,   -28,   -53,   -82,    67,    -8,    84,   -13,    -3,   -29,    62,    34,    47,    95,    27,    61,    69,   -37,   -87,   -76,     0,    83,    -8,    20,    86,  -162,  -269,  -142,    81,   -62,   -67,   -93,     3,    16,    17,   -11,    -4,    62,    39,   132,   -64,   -71,  -198,    60,    -7,    16,   -52,   -55,    32,    34,   -46,    50,   -36,    11,  -123,   -85,   134,    80,   -13,   -46,   109,   127,    -2,     8,     1,    11,   138,    62,  -156,    -6,   -23,    68,     9,   -32,    36,    -8,    30,   -56,   -54,    92,    62,  -180,  -193,   -62,    17,    -8,   -71,   -94,    59,    59,   -29,     1,    19,    60,   -28,    -7,    12,     1,  -112,    10,    -3,  -140,    23,   -48,    49,   -19,   -17,    90,    16,  -104,  -197,  -110,    50,     3,    53,    66,    29,    -2,   -27,   -20,    12,     6,  -117,    34,   -12,    21,   -35,   -51,   -65,   -95,    68,    13,    44,   -17,   -78,   -19,  -157,  -136,  -105,   -76,    24,   -46,     5,    35,    58,   -18,   -18,   -20,   -10,   -19,   -26,   -46,  -152,  -114,  -117,   -24,     1,   -22,    31,    15,    36,   -25,   -61,  -140,  -136,   -88,  -127,  -114,    17,     3,    60,    21,    67,     8,    80,   -17,   -12,    65,    34,    -2,  -125,   -40,   -76,   -16,    56,    10,    39,   -20,    50,    -5,    11,  -100,   -69,   -39,  -124,   -90,   -11,   -72,    68,    94,   110,    25,    72,    -1,     1,    63,    -9,    61,   -30,   -20,   -64,     2,   -60,    13,     6,   -41,    31,    65,   -29,   -10,  -121,    -9,   -42,    71,   -41,   -19,    44,   140,   121,    14,   -10,    74,    95,    78,    59,    31,    84,   -52,   -12,     5,   -42,    32,   -70,    -4,     4,    14,    14,   -74,  -157,    -4,    56,   131,    43,   -10,    71,   119,    63,     5,    -8,    60,    91,    60,    55,   -18,    36,    15,   -99,   -85,   -28,   -68,   -68,    -8,    -5,    78,   128,    56,    13,   140,    65,     4,   -21,    25,    89,    16,   -16,    41,     5,    18,    16,    -4,   -15,   -27,   -19,    77,   107,   137,   148,   -16,   -33,   -17,    31,    37,   156,    63,    99,    74,   -11,  -120,  -123,   -31,   -35,    47,   107,   159,   -17,     8,     4,     8,   -40,  -148,  -140,  -128,   -17,   -11,   140,   -53,   -38,   -44,    11,     9,    96,   -21,   -12,   -23,    28,    -9,    57,     9,   -59,   -47,    67,    46,     0,    13,     7,    16,   -32,   -77,   -60,   -49,  -208,    -7,    94,  -259,  -214,     1,   -25,    72,   -33,  -113,  -214,  -115,   -65,  -108,   -76,   -57,   -42,   -15,    11,     0,   -14,   -16,    -2,    -7,     9,   -29,   -70,  -157,  -196,  -174,  -177,   -68,   -95,  -170,  -174,   -91,   -47,    49,  -105,    -9,   -30,   -17,   -31,    -5,    -3,    18,   -19,   -15,   -10,    -5,    14,    15,    -2,    13,    12,    -3,   -14,    -8,   -26,   -85,   -72,    -3,   -13,   -64,   -23,   -39,    11,    19,   -14,     5,    -5,    -7,     4,     3,     7,     6,    17),
		    62 => (  -11,     7,     3,     8,    18,    -9,     5,     4,    -6,     0,   -19,    -7,   -12,    11,    31,    19,    15,   -12,    14,    18,    -1,    11,    -7,     2,   -14,    -4,   -18,    -2,    17,     8,    -6,   -18,    -2,    -4,   -17,    11,    10,    33,    16,    -9,    -2,     3,    -9,   -54,    51,    23,     5,   -83,   -22,   -20,    -1,     1,     2,    14,    -1,    14,    10,     9,   -13,     3,   -27,   -17,    19,    -9,    19,   -18,    41,   145,   112,   177,    71,   -26,   -47,   -55,  -101,  -249,  -183,   -44,   -39,   -15,     1,    29,    -4,    -1,    -2,   -10,   -18,   -69,   -66,    43,   102,   -12,   -24,    78,   -37,    18,   -31,    10,    -1,    28,    83,     4,  -131,  -111,  -124,   -75,    69,     9,    -4,   -10,    15,    -4,    16,    14,   -46,    40,    47,    66,   172,   165,   -44,    13,    93,    97,    67,   149,   102,    92,     3,    18,    15,   -72,    25,    39,    23,  -109,  -118,   -41,   -70,   -20,    10,    15,    26,     7,   -19,   -72,   -55,   102,   -17,   -57,    35,    14,    55,    44,     3,    52,    56,    -6,    10,   -17,   -87,    57,   130,    18,   -61,   -66,   -78,   -39,     8,     5,    48,    33,   -30,  -116,    35,    42,   -25,     3,   -20,   -42,     0,   -24,    53,    -7,    -3,   -64,    28,   -86,    11,    54,   167,    36,   -61,   -87,   -45,   -24,   -11,     3,   -15,    84,    -3,   -38,  -115,    -7,    52,   -20,    46,    -5,    16,    37,    98,    71,    -9,   -46,   -50,  -105,    29,     0,    75,  -120,   -96,  -131,   -27,   -33,   -58,    45,    40,    11,    86,   -56,   -88,   -43,    27,    -1,    79,    77,   -17,   -48,   -69,    17,    16,     9,   -20,    -5,     3,    -6,    18,     2,   -63,   -78,   -92,   -24,    -5,   -45,   154,   -39,    67,    87,  -106,    13,    -9,     6,    -7,   -69,    15,  -180,  -292,   -29,    43,    32,    -6,   -19,    -2,    -4,    -6,    56,  -137,   -73,    40,   -45,   -14,   -26,    86,    35,   -26,    -9,   -42,    99,    35,   -71,   -62,   -77,  -156,  -228,  -109,   -89,    13,     0,   -52,   -10,   -78,    28,  -135,    62,   -55,   -35,    54,   -23,     3,     2,   -37,    67,    75,   -27,    -2,   -21,   -28,  -170,  -131,  -217,  -247,  -254,   -57,   -28,     5,   -77,   -97,   -77,   -29,   -43,   -64,   101,     4,     4,   -49,    -7,    13,   -10,   -52,   -30,    -7,   -19,   -72,  -212,  -166,  -194,  -191,  -149,  -186,   -68,   -10,   -72,    54,   -13,   -86,   -78,   -12,     5,   -62,    67,   -10,    33,    90,   -42,     4,    14,    64,     1,   -46,  -114,  -190,  -279,  -314,  -302,  -156,  -129,   -58,    88,   -47,   -56,    38,    -5,   -43,  -115,   -92,   -33,   -82,    16,   -37,    -8,    92,    13,     0,   -28,   -35,   -10,   -11,  -130,  -157,  -218,  -234,  -156,   -30,   -19,     8,    25,   -74,   -71,    -8,   -24,  -103,   -71,   -91,   -18,     3,   -29,   -32,     7,    61,    62,   -15,   -47,    -5,   -16,  -136,  -102,   -39,   -85,   -27,    66,    90,    56,   -43,    35,   -27,   -61,   -15,   -71,  -107,   -74,  -138,    15,    -9,   -43,   -19,    56,    63,   133,   -17,    -2,    -9,   -56,  -115,   -76,     3,   -82,   -50,    34,    24,    41,     9,    11,    21,  -136,   -25,   -83,  -160,   -85,  -138,   -38,     2,    -8,   -42,   149,    66,    54,     9,     4,    12,   -15,   -94,   -28,  -110,   -52,   -17,     7,    16,    46,    74,    41,   -18,   -46,   -73,  -126,  -185,  -112,    16,    -3,  -102,  -103,   -77,    73,   -26,    56,    18,    13,   -41,    35,    90,   -24,   -20,   -28,    95,    60,    24,    26,   115,   -27,   -23,  -159,  -118,   -90,   -27,   -41,    11,    18,    -5,   -70,   -52,   197,   -71,   130,    12,   -15,    30,    87,    80,    11,    -8,    66,   128,   -28,    59,    56,   116,    66,   -80,   -56,   -89,  -130,   -36,   -10,     4,     1,   -92,  -118,    69,    74,   112,   143,    -2,    -9,    91,   109,   110,    98,   -94,    44,   -13,   -13,    30,    57,    84,    45,    -4,    63,    11,    82,  -108,    17,    28,    39,    -2,   -17,    63,    77,   101,    19,   -10,    46,   112,    95,    70,    57,   -60,   -42,   -44,    28,    30,    -2,    54,   -18,    -6,    28,    63,   -52,     9,    97,    21,    61,    69,    65,   186,   212,    70,    -9,     4,   -10,   101,    96,    27,     0,   -18,    12,    35,   -45,    48,    18,    29,    -8,    61,    67,    14,  -153,   -35,    53,    68,   -24,    41,   -58,    -6,    29,   -83,   -43,   -14,    -8,   -17,    21,   -58,    43,    -4,    31,    98,    -9,   -18,    50,    -2,   -47,    38,   105,    27,   -98,    71,    33,    -1,    78,    54,    81,    67,    46,   -60,    -6,   -10,     0,   -66,   -35,   -73,  -117,  -195,  -284,  -181,   -78,     9,    23,    35,    37,   145,    11,   -68,    27,    92,    88,   -79,    53,   217,   128,   127,    47,    53,   -16,     4,   -12,   -30,   -21,   -30,   -62,   -47,   -96,  -181,  -185,   -36,   -11,   -34,    -3,   100,   118,    59,   167,   -17,  -165,    13,    36,    28,     4,    65,    61,    49,    14,   -10,     4,   -20,     3,    -7,   -18,   -51,   -43,   -50,   -26,   -15,   -80,    -4,  -107,  -107,   -70,  -177,  -121,   -86,   -37,   -15,   -10,   -59,     8,   -19,   -16,     4,    15,    20,    18,     9,    17,    16,    15,   -20,    12,    13,    11,   -15,   -13,    -9,   -15,     3,    14,   -16,   -17,    13,   -17,   -49,   -38,    -6,   -15,     4,   -12,     2,    17),
		    63 => (   13,    16,    17,     1,     3,    12,   -14,    -1,    -8,   -15,    -4,   -12,   -13,    -6,    -3,   -22,    20,    -7,   -18,    -7,     5,    -7,     2,   -16,     7,   -14,    20,   -12,    19,     3,    -5,    -9,    11,   -19,     5,   -13,    -6,    11,   -17,   -39,   -31,   -48,   -56,   -50,   -29,   -90,   -46,    -4,    11,   -12,    17,     5,     0,    -5,     6,    -5,    10,     3,    13,   -11,     1,    -3,    -1,   -41,  -145,  -132,    70,    65,   -52,  -104,  -142,    -2,   -49,   -36,   -20,   -27,  -103,   -80,   -66,   -76,   -34,     0,     2,    20,    19,    17,    -4,   -34,    -7,    41,    42,   109,    82,    -6,   -46,    79,    70,    59,   134,    45,   -71,   -31,   -60,   -48,    26,     2,  -173,  -257,  -129,   -94,    13,    10,   -14,   -17,   -62,    72,  -133,    15,   129,    48,    23,   -49,   -41,   -37,    18,    62,   101,    -2,    -4,  -124,   -84,   -31,   -51,    35,    18,  -317,  -286,  -148,  -128,    18,   -13,     7,   -18,    -6,   -49,   -32,    64,     8,   -59,  -103,   -20,    80,    95,    15,    37,   -18,    35,    23,   -14,    35,    38,   149,    69,   100,    79,  -269,   -49,    12,    14,   -10,    50,    17,    59,   -27,    34,    91,  -117,   -10,    37,   108,    42,    38,   -59,   -59,   -41,    25,    43,    -1,   118,   136,     3,   -20,    69,  -189,  -138,   -37,    14,    29,     8,    57,   180,    55,   124,    43,    12,    -8,    33,    91,    54,     9,    67,    59,  -101,   -31,    10,    90,     1,    24,  -108,   -20,    32,  -175,  -223,   -67,   -44,    -1,     4,    24,    62,    22,   -33,   -59,    17,    12,    12,    38,    -8,   -58,    78,    46,    33,   -63,    53,   126,    59,    93,   -67,   -43,   -39,  -229,  -221,   -35,    10,   -77,   -19,   -42,    48,    46,    -8,   -36,     6,   -35,   -57,    -6,    -9,    32,    70,    36,    88,    67,    41,    37,   -39,   -53,   -41,   -57,  -263,  -280,  -261,   -92,    -4,  -100,   -68,   -66,   -19,   -78,   -88,   -12,   -37,    11,   -37,     9,    65,    55,   -55,    -1,    33,   127,    33,  -114,   -19,  -182,   -99,   -23,  -177,  -131,  -199,   -84,   -15,   -92,  -103,    16,   -38,   -36,   -30,    37,    -6,   -61,    -3,    31,     7,   -48,   -56,   -51,    -4,   188,    79,     1,   -27,   -97,   -96,   -87,  -240,  -306,  -176,   -17,    -1,   -59,  -128,     0,   -44,    13,   -21,   -63,   -42,   -11,    -5,    38,    87,    -3,   -44,   -22,    49,   106,    87,   100,    65,   -29,   -22,   -38,  -318,  -161,   -82,     0,   -12,   -37,   -95,     2,  -102,   -72,   -54,    -2,    -5,   -88,   -39,   -10,    79,   -17,   -28,   -62,   120,   102,    21,    81,    50,    19,   -69,   -39,   -23,  -198,  -152,   -52,   -30,    42,    -6,   -44,   -97,   -13,     4,   -13,   -30,   -58,    12,    40,    19,   -22,   -61,   -34,    30,   114,    84,   146,    58,    95,   -18,   -16,    53,  -211,  -142,   -23,    -3,    33,    -4,    -1,   -37,   129,   118,     3,    -4,   -36,   -73,   -12,   -59,   -12,   -78,   -47,    37,    57,    44,    94,    52,    23,    42,    29,    99,  -142,   -79,   -42,    -1,    21,     6,    43,    -8,    39,   134,    68,   -32,    -2,   -11,    10,    24,   -50,   -68,   -74,    75,   116,    71,    30,    98,    82,   -18,   -57,    -2,  -197,  -213,   -75,    -6,    -6,   -10,    99,   -22,   -22,   114,   127,   -61,   -46,   -14,     8,    47,   -27,  -112,    13,    80,    78,   -22,   -53,   -14,   -14,   -31,   -43,  -216,  -199,   -96,   -22,   -52,    18,    29,   105,     9,   -21,    97,    44,    12,    32,    67,    31,    -4,  -125,   -36,    62,    67,    -2,   -51,     2,    29,    20,   -47,   -80,  -192,  -202,   -47,   -52,     7,   -82,   -19,     5,    93,    94,    62,   108,    47,    44,    64,   -10,  -142,  -156,   -75,    -5,  -121,  -130,   -41,   -21,   -13,   -52,    76,    16,  -121,  -184,  -182,   -91,    -7,   -45,   -52,   -30,    32,   118,    72,    89,   -20,    29,    40,    55,  -143,  -121,   -76,   -78,  -139,  -149,   -81,   -47,   -56,  -118,   103,   -14,   -32,  -136,   -39,   -19,    -7,   -14,    46,    11,   -28,    38,    77,    13,   -19,    -2,    51,   132,    23,  -103,   -15,    10,    -3,   -56,   -12,    25,   -26,     1,    36,    -7,   -96,  -148,   -66,    16,   -39,   -33,    62,     2,   -24,    36,    59,   -40,    29,   -25,   130,   147,    92,   -80,   -33,    81,    13,    19,    51,   -29,    -2,    -7,    92,   -41,  -193,  -124,  -102,   -15,    -2,    19,    23,    21,     0,    -2,   -25,    18,    19,    78,   128,   155,    33,   101,    74,   104,    56,    37,    79,     8,   -19,    32,   -26,   -80,   -88,  -113,  -157,    -3,    -2,    -1,   -41,   101,     6,   -26,    -2,    94,   133,   134,   143,    15,    27,    34,    68,    76,   128,    42,   -45,   -74,     5,    21,   -22,    -2,  -174,  -133,   -70,   -16,   -10,     3,    13,   -56,   -53,    94,    84,    87,    96,   119,    67,   -19,    36,    -3,    58,    80,    96,    87,    58,    75,    86,    -2,   -89,  -241,  -151,   -51,   -32,     4,   -20,    19,     1,   -57,  -132,    93,    61,    74,  -102,  -103,    25,    20,   -39,  -111,   -94,   -48,    42,    21,   -19,   -35,   -34,   -89,   -85,   -57,   -20,     7,     7,    -1,   -19,    -1,     9,    -5,    -3,   -39,   -14,     7,   -32,   -66,   -82,   -88,   -45,   -82,   -89,   -60,    -2,   -21,   -56,   -74,   -56,   -41,   -22,    -4,     5,    -9,   -15,   -12),
		    64 => (   -7,    -7,   -20,    -4,    10,   -13,    13,    12,    -6,    -3,   -18,   -16,   -30,   -38,   -13,   -16,     5,   -19,   -17,    -8,    -3,   -10,   -19,    -5,    -2,    -3,     4,    16,    -4,    19,   -11,    15,     6,   -11,   -72,   -57,   -41,   -29,   -79,   -63,   -20,   -73,   -29,   -51,   -35,     5,    12,    -4,   -15,   -10,    -8,   -26,     3,   -10,    -6,    -4,    11,    -5,    -2,    15,   -12,    -5,   -93,   -76,   -95,  -148,  -135,  -158,   -97,   -70,   -30,   -33,   -25,   -23,   -34,   -21,   -67,   -16,   -30,   -36,   -16,     3,    -9,    13,    -1,   -13,    13,     8,   -44,   -56,   -19,   -44,  -140,  -204,  -111,    -8,   -47,  -120,   -88,     1,    -2,   -23,    93,    32,   -49,   -17,   -62,     3,    47,    -9,    19,    -1,   -15,     0,   -22,   -39,   -58,     0,    14,   -21,   -46,   -77,    -2,   -27,   -54,   -74,   -57,   -73,   -47,   -66,    -4,    46,   -49,   -37,    29,   123,    48,    43,   -66,   -35,    -4,    16,    -6,   -26,   -25,   -79,   -19,   -76,    40,     0,    62,  -123,  -216,  -279,  -235,   -67,    94,    68,  -117,  -122,   -71,   -85,   -19,    89,     8,    56,   -66,   -19,    17,    14,   -17,   -91,   -72,   -23,    65,    27,    40,    85,   -88,  -215,  -249,  -374,  -266,   -45,    27,    81,   -33,  -171,   -56,    13,    80,   105,   -45,  -108,    26,   -49,   -18,   -91,    -1,   -76,   -71,     2,   -11,     2,    86,   127,    45,  -130,  -314,  -431,  -140,    74,    52,    65,  -150,   -19,    47,    98,   210,    58,  -139,  -128,   -32,  -122,   -49,   -74,   -28,   -96,   -83,   -36,    44,    -2,    32,   129,    54,   -81,  -376,  -279,   -77,    28,   100,   -11,  -129,   -89,    23,    79,    22,    61,  -158,   -21,   -98,  -102,     7,   -33,   -11,  -110,   -72,   -20,   -71,    60,    93,    89,    66,   -46,  -139,  -110,   -43,    -2,    38,   -38,   -37,     1,    -6,    14,     3,    86,   -63,   -41,   -68,   -39,   -11,    18,     3,  -112,   -12,     2,   -21,    44,    63,   137,    91,    11,  -133,  -170,   -29,    71,    22,     6,     9,   -19,   -64,   -59,   -50,   -14,    51,    33,   -37,   -60,    13,   -32,   -20,   -72,    22,    39,    28,    13,    95,   132,    53,   -61,  -120,  -116,   -82,   -30,   -18,     5,   -61,   -30,    13,   -23,    13,   -47,   -21,    49,   -47,  -113,    17,   -31,    20,  -148,   -56,   -14,    53,   -29,    18,    86,    44,   -11,   -16,    20,   -23,    31,    -6,     9,   -11,    27,    74,   -14,     8,  -117,   -99,   -21,   -54,  -108,   -14,    -3,   -39,   -96,  -110,   -75,    56,    40,   -24,    94,    39,     1,    -1,    49,    16,    52,    -5,    18,    63,   115,   -23,    19,    19,  -151,  -152,    -6,   -62,    16,   -18,    29,  -115,   -27,     8,   -43,   -50,    32,   -75,   -50,    -6,   -19,     7,   -25,    31,    93,    24,    73,    62,    15,    25,    66,   -56,  -167,  -125,    22,   130,    14,    14,    -9,    78,    13,    96,   -10,    80,    -8,    85,   -57,   -42,   -69,   -82,     2,   -43,    63,    20,     3,   -27,    14,  -116,   -20,    28,    69,   -97,    47,   165,    19,     8,     4,   -59,    57,   -20,   -88,   -73,    49,   -15,    25,   -17,   -43,   -27,   -26,   -77,    27,   -22,    -9,    -7,   -63,  -175,     1,    22,   -13,   115,   144,    48,   -18,    17,    -6,   -30,    10,     7,   -65,   -58,    30,    26,    10,   -37,   -49,   -68,   -47,   -93,    29,     4,   -36,     0,   -91,   -77,    60,   -18,    29,    54,   156,   123,   -41,    -8,    -2,   -27,   -15,   -14,   -87,   -66,    15,    -9,     1,   -74,  -124,  -126,   -39,   -59,    40,   -62,   -44,    26,   -30,   -48,   -14,   -26,    12,   -59,   -29,     7,   -35,    18,   -22,   -54,    24,   -39,   -74,   -23,    36,   -48,   -44,   -66,  -115,  -104,    -3,   -17,    60,   -12,   -52,    87,   -31,  -110,   -40,    -7,   -47,   -61,   -80,     4,   -38,    16,    -2,    -1,   -54,   -71,   -73,   -69,    50,   -32,   -35,   -87,   -45,  -125,   -50,   -26,    10,    25,   -16,    13,    33,   -16,    22,    42,     8,   -19,  -128,    -2,     1,    14,    15,   -66,   -78,     0,    -2,   -26,    50,    21,   -41,   -75,  -186,  -110,   -18,    82,    19,   -20,   -25,    -6,    26,     7,    -1,   -37,    72,    -4,  -138,   -66,    -9,    10,     6,     7,   -48,   -74,     9,    22,   -13,    35,   -66,  -111,  -128,   -84,   -21,    20,    21,   -45,   -94,   -22,    90,     8,    28,    44,   113,   -55,   -58,    38,    -2,   -11,    11,   -16,   -18,   -44,   -56,     6,    -9,   -39,   -13,   -44,  -147,   -26,    36,    29,   -14,   -47,   -99,    43,    68,   -50,    99,     6,   -50,  -115,    41,    14,    -4,    -3,    -9,    -9,     5,   -56,   -46,   -44,   -71,    18,   -17,   -49,   -58,   -43,   -20,    41,    54,     1,    -1,    30,    22,    25,    38,    82,   -56,  -137,    11,   -36,    19,    -7,    16,    -7,    -2,   -24,   -11,   -46,   -34,    37,   -25,   -71,   -69,    -5,    51,  -110,   -60,   -54,    39,    38,    20,    82,    46,   -42,   -47,   -59,   -33,   -27,    12,    16,   -20,   -10,   -40,   -20,   -39,   -18,    -6,    19,     9,   -58,   -35,   -34,  -224,  -247,  -233,  -121,   -17,   -54,  -134,  -176,  -162,  -200,    -9,   -56,     1,   -17,    -3,    13,    11,    -4,    -7,    13,     3,   -32,   -73,   -80,   -46,   -35,   -81,   -78,   -71,   -79,   -28,   -84,  -134,   -99,   -78,   -91,  -103,  -110,    -3,     9,    -5,    -2,    19),
		    65 => (  -15,    15,     6,    -5,   -15,     1,    -3,    13,   -20,   -19,     7,    -7,   -12,    -2,     6,     8,     8,    -8,   -20,   -17,    13,   -20,   -15,    10,   -16,   -12,   -18,   -11,    -3,    -2,   -17,    -8,     3,    -5,   -12,    15,    18,    -5,   -27,    -6,   -20,   -24,   -30,   -37,   -39,   -32,   -38,    -4,   -15,    -9,    11,    12,     5,   -14,    -5,   -18,    -1,    10,   -20,    15,   -20,     0,     2,   -10,   -32,   -10,   -19,   -92,   -88,  -101,  -125,   -61,   -75,    75,     5,    39,    98,   -28,    -6,   -27,   -38,   -24,   -17,    -2,     6,   -17,    -5,    -6,    17,   -17,   -40,   -31,   -52,   -77,    18,   -30,   -72,   -27,   -23,    30,   -67,    69,    53,    52,   123,   133,    83,   -93,   -73,    36,   129,    11,    -6,    15,   -45,   -26,   -30,   -42,  -112,   -54,   -99,    78,    75,    -2,    12,  -113,   -65,   -33,  -125,   -32,    68,   -54,   -54,    33,    -5,   -46,   -16,    95,    76,   -72,   -11,    15,   -67,   -49,   -39,   -63,  -208,  -221,   -50,    83,    18,    -9,    44,   102,   -20,  -213,   -80,   -58,   -84,   -46,    90,    51,    50,   -51,   -52,    61,    96,   -32,   -14,   -19,    84,   -43,   -72,  -158,  -204,  -215,  -112,   -22,    59,   -30,   109,   105,   -11,   -65,   -72,     0,   -16,    33,   101,    41,    86,    -7,     6,   175,   182,    59,    18,   -18,    81,   -95,   -53,   -54,  -181,  -177,  -102,    61,     9,    -8,    86,    70,   -59,    55,    92,    94,   105,   114,   127,    30,    80,    -9,   -48,    75,   182,     4,    -6,   -41,   -79,   -77,   -45,  -190,  -161,   -81,   -15,   -23,   -57,   -45,    -8,   -50,     7,    56,    83,   105,   181,   138,   106,   -18,    30,    67,    -7,   -22,    97,    55,     9,    -6,  -127,  -137,  -128,  -121,   -75,   -67,  -100,     0,   -28,   -35,   -65,   -43,  -102,  -101,   -52,   105,    45,   -15,   -81,   -63,    -9,   -30,   -46,    76,    15,    92,    17,   -23,   -11,   -22,    21,   -71,   -26,  -141,   -57,    43,   -60,     2,     9,   -59,  -130,  -298,  -312,  -244,  -194,  -267,  -231,   -85,  -107,  -239,  -106,     9,   105,   117,   -13,    -6,     3,   -25,   137,     2,  -141,   -88,   -50,     4,     5,   -42,     3,   -44,   -73,  -192,  -247,  -345,  -316,  -292,  -323,  -199,  -160,  -198,  -128,   -69,    18,   103,     7,   -11,     4,    36,    67,   -60,  -120,   -47,   -38,   -23,    42,    14,    -4,   100,    17,   -14,   -54,  -133,   -86,  -133,  -157,  -214,  -214,  -163,  -130,   -55,   -13,   -51,    -3,   -19,     5,    59,    31,   -44,   -22,    10,   -46,   -71,   -29,   -39,   -18,    48,    59,    46,   -48,   -53,   -64,   -75,   -22,  -170,  -278,  -166,  -134,   -45,    -8,   -55,     3,   -33,   -25,    87,    27,   -74,   -33,    41,    17,    28,    -1,    23,    31,   -10,   -37,    22,   -50,   -28,   -52,    -7,    80,   -23,   -62,   -50,   -51,   -30,   -14,   -14,    28,   -30,   -97,   -59,    38,     5,    64,   -66,   -35,    63,   -11,     3,    22,   -50,   -16,   -31,    30,   -40,    -5,   -46,    38,   102,   -45,   -26,    39,     8,   -26,   -62,     9,   -21,   -59,   -55,   -26,   -14,   -69,  -106,    -5,    11,    40,    53,    16,    52,     5,   -64,    -6,    19,  -101,    14,   -18,   -45,  -103,  -128,    -5,   -59,  -101,   -68,     0,   -19,   -79,     0,    14,   -82,   -94,   -34,   -78,   -25,    72,    65,    32,    75,   -43,   -31,   -28,   -26,   -37,    11,    44,   -55,   -81,  -156,   -22,   -71,   -19,   -89,     3,   -21,   -68,    30,    29,    -9,  -127,  -183,  -124,  -159,   -81,    55,   -24,   -22,  -106,   -89,    65,    28,    21,    -1,    84,   -71,   -55,    -4,    22,   -17,   -85,   -50,    17,     1,   -52,   -86,   132,    -4,    -2,   -87,   -97,  -219,  -201,  -228,   -80,    15,   -59,  -125,     1,    58,    21,   -25,    76,   -72,   -63,    55,    59,   -44,   -13,   -26,     5,   -24,   -38,   -45,    24,    64,    22,    14,   -30,  -119,   -17,   -89,  -155,   -21,   -24,    26,   -54,    17,    18,    62,    53,   -29,   -11,    37,   -13,   -21,   -38,    15,     3,   -15,   -95,    -7,    98,    57,    11,    12,    -3,    31,    43,   -10,   -13,    49,    19,    14,   -43,   -46,    20,    84,    17,   -52,    58,    41,   -36,   -19,   -65,     4,    17,    12,  -109,   102,    43,   -61,   -29,   -49,    31,   126,    98,    79,    19,   -61,    36,   -42,   -24,    33,   -14,    -5,    22,    -5,    -9,   118,   -10,   -32,   -16,   -18,    -4,    10,    45,   126,   114,    57,    80,    12,    18,   -74,    28,    62,    27,     6,   -17,    12,   -64,   -31,   -18,    15,    20,    -2,    33,   126,   -25,   -80,    14,   -15,    19,    15,   -67,    26,   -34,   -34,    -7,     6,   -30,     9,    18,   -38,   -24,   -13,     7,     5,   -61,   -39,    48,   -28,   -70,    28,   164,    39,    62,   -92,   -51,    -9,   -17,   -20,   -18,   145,  -111,  -113,   -44,   -70,  -106,    11,   -61,   -50,    14,    82,   -27,   -24,  -177,    31,    36,    19,    51,   134,   205,    99,    61,     1,     4,     1,     1,    10,     0,   -10,   -17,   -35,   -31,   -37,   -55,  -101,   -25,    74,    87,    46,  -169,  -198,  -166,  -172,   -82,    42,   -62,    55,    48,   -20,   -16,    -1,   -10,   -13,    19,     0,    -9,     2,     2,   -18,     5,   -13,   -19,   -32,    -3,     7,    19,    32,   -43,    -6,    -6,    -4,   -26,   -12,     9,   -23,   -49,   -21,   -12,    -6,    19,     5),
		    66 => (   -2,     8,     4,   -13,    15,    17,    -6,    -7,    10,   -19,    -5,     6,    67,    81,    11,   -14,    -6,     0,   -16,   -12,    -5,    15,     8,    14,    15,   -11,     2,     1,    -5,    15,   -10,   -18,     3,     4,    38,    36,    17,     6,    88,    11,    38,    96,   -43,   -39,   -20,    18,    54,    84,    92,    75,    69,    61,    -3,    20,    -4,     0,    -4,   -16,     5,   -23,    27,    61,    40,    -9,    22,    75,    67,    69,    46,    69,    58,   -29,    59,    62,    82,   132,   111,    62,   188,   126,    95,    77,     2,     6,    16,    11,  -111,    61,   -13,   111,   124,   117,   160,   163,   188,   190,   244,   157,   213,   149,    38,    16,    20,    16,   -62,   -78,   -54,    -4,    76,  -154,  -132,     5,    12,   -14,   -86,     8,    62,   101,   110,   154,    77,   165,   144,    78,   142,    24,   164,   136,    36,    61,    27,    85,   102,    55,   -28,   -42,   -49,  -105,   -41,   120,   -19,   -10,   -43,   -90,   141,    63,    85,    99,    63,    71,   128,    30,   -73,    65,   136,    70,    19,    99,    12,   -40,    24,   -86,   -15,    10,   112,    53,   106,    39,     8,     1,     2,     8,   106,    39,   115,    64,   -16,    48,   -27,   -64,    39,    32,    34,    14,     9,     3,  -127,    30,   -11,   -75,   -75,   -66,   -17,    42,    98,   139,     8,   -17,    -7,   -39,   109,    75,    41,    39,    10,   -38,   -61,   -28,   -91,  -121,    44,   -43,   -18,   -40,   -39,    12,   -39,   -23,   -27,   -24,    41,    12,    86,    94,   -12,   -45,   -57,  -210,   123,    42,    23,   -47,     3,    64,   -56,   -62,   -37,   -73,     3,   -96,  -170,   -74,   -42,   -15,    41,    43,   -40,   -75,   -75,  -170,   -13,  -132,     0,   -17,   -73,  -115,    97,   -23,   -68,   -47,    15,   -39,   -59,   -73,  -107,  -129,     0,     6,   -69,  -165,   -28,   -31,   -15,    81,   -15,   -19,  -115,  -207,  -128,  -114,   -12,   -17,   -81,   -63,    29,    10,   -71,   -76,   -18,   -46,   -28,  -106,  -130,   -60,    16,   -52,  -143,   -87,  -120,   -89,    16,     9,   -97,   -82,  -141,  -152,  -127,  -125,    -5,   -20,   -15,  -128,    28,    17,    -7,   -19,   -62,   -23,   -53,  -101,    11,   -11,   -20,   -86,   -74,   -65,   -77,   -41,   -39,     9,   -86,   -20,   -65,  -130,  -138,   -95,    20,   -16,   -60,  -120,   -19,    33,    90,    26,   -32,    31,    -7,    15,   -30,    50,   -67,   -44,  -107,   -69,   -97,   -71,    52,    38,   -59,    57,    83,    -9,  -186,   -95,    -7,    12,   -42,  -106,   -48,    41,   -12,   -49,   -46,    83,   104,    70,    68,    35,    46,    16,   -24,  -122,   -34,    51,    58,    62,   -40,    64,    45,   -59,  -194,    -3,    -1,    -8,   -19,  -102,  -144,    47,   -60,  -100,    30,    35,   103,   102,   109,    56,    23,   -73,   -15,   -70,    30,    36,    18,    46,    47,   -54,   -27,   103,  -155,   -33,     1,    -7,   -61,   -70,  -161,   -58,   -54,   -18,   -48,   -16,    27,    54,     1,   123,    81,   -51,   -55,  -131,     8,    68,   -10,    21,   -95,    12,     2,    89,   -66,  -187,    13,    -2,   -93,   -73,   -37,    30,    28,    42,   -46,    55,    53,    22,   -36,   -67,   -43,   -40,   -46,   -61,    87,    98,   -40,   -32,    30,    -5,   -30,    68,  -101,  -154,   -18,     6,  -108,  -108,   -72,    92,     5,    35,   -21,   -72,   -40,   -18,   -37,   -64,    11,    39,    39,    67,    54,    64,    53,   -24,   -21,   -45,   -23,    61,   -95,  -218,    16,   -14,  -103,  -168,   -31,   -12,   -70,    16,    -9,    20,    68,  -114,    -7,   -14,    -1,   -79,     7,    65,   167,   134,    13,   -51,     5,    27,    21,   102,     8,   -94,    13,     1,  -123,  -136,    16,    50,    44,   -17,     9,     6,   125,   126,    72,    31,    19,    36,     5,    92,    -4,   136,   -13,    -8,   -22,   -52,  -108,    33,   -64,    -4,     2,    -7,  -112,  -169,    -7,    -7,     4,    53,    19,    30,   107,   116,    98,   -62,    27,    28,    23,    65,    71,    61,    64,    -7,   -12,  -123,  -148,   -42,   -40,    -3,   -10,   -18,  -143,  -153,  -116,  -136,   -38,    90,   113,     0,    57,     6,   166,    77,    32,    18,   135,    84,    73,    44,    28,   -44,   -30,  -131,   -67,    -7,   -12,   -22,     3,    10,  -104,  -119,  -215,  -269,  -357,     1,     4,    66,    34,    21,     7,     2,    11,    91,   107,   154,    96,    12,    31,    29,  -109,   -95,  -237,   -63,   -26,   -17,    -4,    18,    17,  -130,  -162,  -185,  -170,   -24,   -45,     7,   -71,    20,    80,   -22,    40,    87,     6,   -72,    21,     3,    11,    55,  -132,  -163,  -157,  -108,  -128,    20,   -18,     7,   -11,   -20,   -52,   -61,   -90,  -172,  -234,  -306,  -211,  -270,  -133,  -132,   -84,    22,    43,    62,   138,  -210,   -32,  -112,   -95,   -88,   -68,   -43,   -18,    -1,    11,    13,    -6,    -9,   -18,   -39,   -69,   -67,   -49,   -64,   -75,    27,    61,   -38,   -33,   -57,   -98,   -96,   -53,  -156,  -144,   -27,   -77,   -76,   -61,    16,    -9,    17,     6,    16,     1,    -4,   -17,   -29,    13,   -22,    -7,   -22,   -17,   -35,   -13,     6,    -9,   -31,    -5,   -20,    -2,   -22,   -19,    18,   -18,   -19,    11,    14,     9,    16,     1,     9,   -14,    18,     7,     7,    -1,    -2,    20,    -7,   -11,   -14,     9,     9,   -12,     0,    -8,   -17,     3,     6,   -19,   -23,   -11,    10,   -17,    -4,     7,     3),
		    67 => (  -14,   -15,    13,   -14,     2,     7,     7,    14,   -19,   -15,    14,     9,    15,     3,    -5,     2,    19,    11,    13,    17,    -8,   -15,    14,    18,     7,    17,   -16,   -19,    11,   -12,    -4,     0,     8,    -6,    17,    -9,    13,     7,    -7,   -21,   -20,   -29,   -32,   -74,   -75,   -47,    -6,     4,     3,   -13,    -8,   -12,    11,    13,     4,    12,   -13,   -11,    19,   -12,     1,    -6,   -19,    -9,   -31,    23,   -16,   -70,  -114,   -49,   -51,   -48,    16,    -6,   -17,   -18,   -22,   -24,    -7,    18,     4,    -4,     3,   -12,   -15,    14,   -14,     0,   -30,   -60,   -69,  -112,   -49,   -20,   -49,   -75,  -136,  -139,  -100,   -97,   -63,   -49,   -22,     2,   -18,    16,   -41,   -12,   -31,   -27,    15,     1,    17,     0,    -1,   -14,   -51,   -12,   -84,   -85,  -120,  -147,  -212,     8,    18,     8,   -32,  -100,  -234,  -175,  -130,  -137,  -103,    11,   -66,   -83,   -90,   -56,   -24,   -16,   -11,   -15,    -3,   -53,   -77,   -30,  -157,     6,   155,    30,   -31,     2,    50,   -19,    56,    15,    23,    -2,   119,    -6,   -81,   -40,   -34,   -71,  -122,   -18,   -27,   -10,    -8,     6,    56,   -40,   -39,   -32,  -101,    42,    67,   107,    51,   -18,   -26,   -29,   -34,    47,    22,     4,    75,    29,  -148,   -67,     8,   -80,   -81,   -57,   -59,   -30,    15,    44,    62,    -2,    35,     1,    43,    39,    57,    43,   -14,   -41,   -79,   -83,   -92,    -8,    76,    79,    60,    97,   144,    26,   -60,   -64,  -109,   -62,   -55,   -31,   -81,    24,   154,    10,    62,    43,    25,   100,    90,     8,   -18,   -36,   -25,   -70,     9,    91,    23,    22,    39,    47,    95,    52,   -11,  -140,   -90,   -19,   -41,   -30,    28,    32,    36,    76,    72,  -109,   -27,     6,    33,    -7,    28,   -60,   -37,    28,     4,   -23,    29,    83,   -26,   -21,    43,   -71,   -42,   -86,   -54,   -12,   -78,    30,    23,    10,   -23,    19,   105,   -27,   -26,    17,   -43,    38,    24,   -69,  -133,    25,   -10,    16,    15,   -19,     3,    21,   -26,   -98,   -26,   -73,   -74,   -12,   -54,     4,    26,    28,   -16,   -78,     0,    14,   -38,    60,    26,   -42,    15,    -2,  -133,   -87,    -2,   118,   -11,    -4,     1,   -10,   -81,   -55,   -76,  -157,   -85,   -92,   -72,    27,    14,    14,   -62,   -19,   -61,   -17,   -65,    57,   -12,   -87,   -50,  -147,  -152,  -104,   -62,    76,   -36,  -103,   -33,  -137,   -81,   -80,  -147,  -145,  -161,   -41,   -48,    10,   -10,    52,    58,   -25,   -18,   -17,   -53,    -4,     9,   -59,   -83,  -139,  -276,  -180,   -97,   -20,   -51,    -6,   -41,  -128,  -111,  -111,  -134,  -176,  -155,   -21,   -94,   -45,    -4,    64,    21,    66,    -8,    48,  -108,   -55,  -105,  -164,  -290,  -228,  -148,  -109,   -82,     3,   -80,    27,    65,    16,   -46,    31,   -94,  -116,   -44,   -24,   -75,   -29,    15,    -8,    -2,    52,    41,   -24,   -75,  -200,  -122,  -110,  -158,    15,   -28,   -21,   -95,    -4,    -8,    73,    85,    21,    51,    46,   -23,    10,    15,    39,   -25,   -36,     8,     8,     3,   -53,   -34,    -1,  -126,   -63,   111,   -38,   -34,   101,    33,    -5,   -20,    85,    35,    15,    76,   -47,   -14,   -81,   -51,   -23,   -19,  -123,   -59,   -17,    17,    -1,   -58,   -48,   -74,  -141,   -70,   -50,   -29,     5,   -87,     8,   -23,     7,   -27,    33,    25,    73,    45,     5,  -140,  -148,  -121,  -101,   -39,  -192,  -107,  -133,    25,     7,    27,   -70,   -62,   -20,   -53,     7,   -44,    24,    -7,    11,   -83,    60,    24,   104,    -9,   114,   -58,    40,    65,    12,   -97,  -125,   -74,  -147,    13,   -93,    -7,     9,     5,    -8,   -19,  -134,   -50,   -50,    45,   -37,   -36,   -95,   -44,   -42,    98,   139,   -62,   -55,   -46,    41,    68,    74,   -46,   -15,    26,   -61,   -80,   -69,    -2,    54,   -28,    -5,   -23,  -108,   -84,    -3,    28,    41,   -21,  -201,   -60,   -27,    41,    32,   -58,  -106,   -43,   -18,    61,    -7,   -49,  -166,   -87,   -47,   -83,    14,   -23,    13,   -25,   -40,   -33,  -113,  -155,  -142,    31,   -41,   -67,  -109,   -22,     6,    57,    22,    86,  -114,   -48,   -72,   -44,    16,   -57,  -197,  -107,  -106,    -6,    -6,   -29,     9,   -16,   -11,   -25,   -94,  -127,  -123,   -72,   -94,   -51,  -106,   -62,    72,    17,    61,    18,    32,   -78,   -40,   -55,  -166,  -249,  -179,  -106,   -61,  -100,     6,    -2,    19,   -27,   -66,  -139,  -144,  -126,  -193,  -163,  -225,  -154,  -133,   -76,   -35,   -37,     3,   -26,  -119,  -177,  -123,  -113,  -119,  -112,   -88,    28,   -59,   -91,   -16,   -19,   -16,    11,     0,   -54,  -141,  -167,  -166,  -242,  -230,  -169,  -113,   -29,    -2,    26,    87,   -17,   -30,  -159,   -99,   -14,   -43,   -13,   -77,   -49,   -52,   -14,    -6,   -10,     0,   -92,     0,    13,   -60,   -92,  -130,  -132,  -208,  -126,    34,   -56,   -48,   -17,   109,    11,    29,    -7,    55,    75,    52,   -33,   -61,     2,    -9,   -15,    -7,     3,   -10,    -1,    -5,   -46,   -50,   -14,    60,    35,    37,   -50,   -37,    53,    79,    42,    16,    -2,    27,   226,   185,   114,    32,   -21,   -31,   -10,     1,    -1,    -1,   -12,    -7,    -2,    10,    38,     7,    -9,   -35,     2,    81,   112,    67,    51,    49,    20,    88,    78,   134,   200,   127,    59,   -10,   -39,    18,     3,   -16,   -11,   -18),
		    68 => (   13,    19,    15,     4,    -9,   -16,     7,   -19,     6,   -11,   -19,    -2,    -7,     8,     3,    12,    11,     6,    -6,     4,     5,     5,    -8,    -4,    -1,   -19,    20,     6,    16,   -10,   -10,   -13,    17,    13,    17,   -16,     7,     1,    14,    -7,     5,     0,    -4,   -17,   -84,   -72,     4,     0,   -10,   -19,   -17,     9,     4,    -6,    12,    -8,    -5,   -18,   -15,   -13,   -20,     3,     7,   -18,    21,   -23,   -45,   -12,     1,   -15,    10,    -9,   -42,    -5,     2,    -2,   -16,   -45,   -20,   -40,    -6,   -16,    17,    14,   -16,    -8,     2,    -7,   -17,   -35,   -21,   -43,   -32,   -29,    -2,     1,   -16,     5,   -66,   -46,   -15,    -7,    25,   -17,   -41,     7,    18,    17,   -16,     5,   -32,    12,    17,   -11,     7,   -30,   -20,   -20,   -59,   -60,    15,     3,   -13,    59,    58,   -41,    -3,  -103,   -84,   -18,    33,     7,    25,   -36,   -40,    -4,   -26,     9,     3,     2,   -17,   -19,     0,   -34,   -92,  -110,    -5,   -16,     3,     4,   -47,   -24,   -49,   -45,    13,   -24,   -66,   -27,   -34,   -42,   -14,   -31,   -50,   -28,   -16,    42,     2,   -32,   -18,     3,   -40,   -81,   -14,    15,   -15,    44,   -12,   -40,   -63,   -97,   -38,   -91,   -51,    -2,    -7,     6,   -23,   -34,   -26,   -57,   -23,   -15,   -16,   -29,   -18,    -1,     9,    -9,   -31,     1,    21,    94,    18,    24,    10,   -19,   -23,   -58,    13,     7,    23,    34,    29,    18,     7,    21,   -58,   -19,    17,     3,    27,    -4,     7,   -19,    -6,   -43,   -14,    76,   117,   127,    47,   -16,   -73,   -52,   -16,    27,    12,    18,    -7,   -49,   -65,   -37,   -36,   -35,     7,    14,    21,   -24,   -18,    11,   -35,    -6,     5,   -52,   -68,    62,    99,   115,    44,   -41,  -104,   -63,    38,   -65,   -65,   -37,   -50,   -96,   -85,   -21,   -39,    42,    50,    54,    14,    -4,     5,    55,   -30,   -23,   -13,   -35,   -68,    38,    28,    90,    76,    47,   -50,    14,    43,   -11,    -1,   -34,   -37,   -52,   -43,     2,   -32,     3,    20,    -6,   -40,   -42,    -6,   -56,   -28,   -31,    -1,    -9,   -87,   -46,   -39,    -7,    75,    95,    64,    94,    68,    20,   -20,   -37,   -52,   -27,   -28,   -38,   -75,    -7,   -23,   -21,    14,   -21,   -42,   -29,    -2,   -73,     5,     7,   -53,  -113,   -88,   -21,    10,   -39,    37,    18,    63,     7,    -1,   -82,   -83,     0,     0,   -18,   -15,   -55,   -53,    40,    15,   -21,   -32,   -53,   -56,   -89,     4,   -24,   -81,  -124,   -48,   -75,   -77,   -78,   -77,   -66,   -37,    11,     8,   -48,    22,    25,     7,   -53,   -48,   -89,   -70,   -14,   -10,   -19,   -52,   -88,   -54,    27,   -33,   -22,    17,  -122,   -53,   -47,   -67,   -99,   -92,  -138,   -67,   -94,   -55,    -4,   -22,   -72,   -77,    -9,     2,   -33,   -76,   -29,   -12,   -16,   -63,   -28,  -140,   -15,     4,    18,   -26,    25,     3,   -27,   -49,   -89,   -56,   -79,   -59,   -32,   -45,    -4,    -7,   -25,    -7,   -26,    -7,   -46,    -6,   -54,   -43,   -46,   -54,    27,   -49,   -58,    11,   -29,    -7,    33,    -3,   -27,   -64,   -38,   -16,   -72,    -2,    18,     2,   -39,   -82,   -88,    31,    37,   -41,   -29,   -11,     0,     2,   -39,   -38,    14,   -64,   -46,    18,    -2,    -2,    50,   -17,   -48,   -42,   -32,   -52,   -50,    52,    59,    -8,   -58,   -61,   -96,   -51,    27,     4,   -44,   -33,    18,    38,   -54,   -25,   -31,   -18,   -27,    -4,   -17,   -11,     7,   -39,   -30,   -43,   -32,   -58,   -49,    20,     3,    25,     4,   -82,   -66,   -65,    50,    17,   -20,   -74,   -34,    64,   -18,   -33,    12,    -6,   -57,    10,     9,   -23,    -9,   -46,   -19,   -15,   -30,  -112,    -6,    45,    48,    -9,     7,   -56,   -68,   -68,   -13,    57,    19,   -21,     9,    34,    41,    -2,     9,   -41,   -45,   -14,    -6,   -40,   -33,   -38,   -25,   -12,   -36,   -73,   -12,    23,    62,    27,   -72,   -89,   -59,   -84,   -17,    30,     7,    -2,    -6,    61,    18,   -18,    -5,   -53,     3,   -28,   -32,   -13,   -55,   -17,   -19,   -71,   -52,   -42,   -31,   -25,    21,    29,   -15,   -45,   -41,   -79,    10,    27,    13,     9,    15,    64,    -1,   -23,   -27,   -25,    -5,   -63,   -26,   -25,   -39,   -26,   -48,   -38,   -28,   -43,   -56,   -13,   -12,   -25,   -18,   -38,   -28,   -49,    26,   -13,   -10,     1,    46,    19,   -19,   -68,   -26,    -8,     5,    15,    17,    -2,   -32,   -32,   -60,   -59,   -43,   -21,   -45,    -8,   -67,   -30,    37,   -30,     1,    26,     6,   -18,     4,    33,    59,    23,   -36,    -3,    -1,   -87,     0,   -13,    18,   -23,     4,   -16,   -40,   -35,    17,   -31,    -9,     1,   -60,   -55,   -60,    19,    46,    51,   -47,   -81,   -51,    -3,   -51,   -60,   -19,   -22,   -28,   -11,    16,     9,   -14,   -33,   -29,   -31,   -34,   -45,   -52,   -36,     3,    49,   -35,   -46,   -32,     1,    19,     3,   -12,   -39,   -32,   -61,   -47,     1,    -6,   -23,   -13,   -37,   -17,     0,    -9,    -5,   -10,     1,   -32,   -25,   -53,   -26,   -60,   -54,   -50,   -55,   -41,   -75,   -64,   -20,    -2,     2,   -81,   -98,    -7,   -63,     1,     9,    11,     1,     3,    -5,    19,    16,     5,    -6,     9,    -4,   -12,   -10,   -31,   -27,   -12,     2,   -27,   -22,   -14,   -32,   -26,   -54,   -12,    -7,    -9,   -18,   -15,    -3,    15,   -17,     4),
		    69 => (  -13,   -17,    13,    14,    15,    15,     1,    19,   -18,    13,    18,    16,    -5,     7,     3,     9,   -17,   -13,    19,   -12,     3,    -8,     6,    -5,     3,   -14,    -2,     5,     4,    13,    19,   -16,     4,    -1,   -13,   -35,   -43,   -38,   -31,   -51,   -61,   -92,   -48,  -106,   -92,   -97,   -49,     3,    12,   -16,   -50,     4,    16,   -15,   -14,   -13,   -14,    -6,   -15,   -73,   -82,   -15,   -14,   -86,  -109,   -47,   -53,   -78,     7,     0,  -226,  -126,  -117,   -73,  -129,   -93,  -171,  -192,  -139,  -116,   -70,   -36,    16,     4,     3,    -5,    -9,   -95,  -122,  -107,   -67,  -116,  -255,  -319,  -429,  -383,  -256,  -332,  -306,  -332,  -434,  -377,  -120,  -162,  -267,  -233,  -193,  -110,   -96,   -61,    19,    11,    18,   -14,   -53,   -85,  -139,  -176,  -251,  -175,  -195,  -215,  -133,   -37,    15,   -20,   -69,   -69,   -59,  -125,  -230,  -451,  -287,  -237,  -236,  -124,  -106,  -172,  -123,     9,    -8,     3,   -53,   -79,   -63,  -103,  -108,   -70,  -157,    26,    29,     9,    58,   124,    41,    48,   105,   104,   -15,   -64,  -132,   -55,  -262,  -111,  -164,  -169,  -118,   -30,    -9,    18,   -53,  -172,  -127,  -157,   -82,   -51,    -5,    81,    82,   -40,   -33,   120,    52,   123,   194,   121,    27,    42,   -28,   -14,   -33,    30,     5,   -56,  -128,  -150,     2,   -60,  -110,  -145,   -92,  -168,   -23,   -16,   -29,    33,    30,   -22,    70,   146,   134,   114,   235,   141,     0,    43,    71,    -8,    38,    37,     0,    13,  -140,  -115,  -102,  -131,  -101,  -114,  -125,   -12,    47,   -22,     1,    38,    13,    10,    95,    84,   129,   195,   156,   108,    97,   118,     9,    48,    32,    75,    79,     5,  -134,   -74,   -18,   -91,  -133,  -140,    85,    32,    80,    39,    46,    86,    17,   -24,    39,   112,   104,    66,    48,    38,    32,    26,    93,     1,    -6,   -35,   -42,  -142,  -174,  -116,    -8,   -63,  -189,   -89,    84,    86,     4,    15,   -11,   -14,     5,    -6,    63,    44,    25,   -81,     2,   -49,    -2,    -5,    24,   -87,   -52,   -42,  -111,    74,  -182,   -73,    -9,  -293,    -2,   -62,    25,    99,    42,   -35,   -87,   -24,   -24,   -68,    -2,  -111,   -94,  -100,    -4,    26,   -74,   -37,    64,   -42,  -126,   -81,  -106,   -11,  -152,   -61,     3,   -31,   -21,   -58,    68,    41,    31,   -41,   -98,   -99,   -36,     2,   -85,  -107,   -52,   -82,   -44,    23,   -61,   -92,    22,   -69,   -60,   -11,  -126,  -213,  -128,   -89,   -20,   -62,   -94,   -66,    32,   -30,    26,    18,     4,   -60,   -15,   -61,     5,   -33,   -51,   -94,    22,     2,   -29,   -48,   -64,     4,   -76,   -73,   -55,  -154,   -94,   -26,   -34,   -55,   -58,   -14,    44,   -22,   -11,    27,     3,   -10,     7,   -36,    50,   -92,   -61,    37,     8,     0,    42,    34,   -10,   -61,   -87,  -178,   -79,  -185,  -111,     1,    -1,    -9,  -131,   -56,    23,    16,    47,    11,    66,    42,   -67,   -93,   -79,   -26,    47,    38,    73,    39,    62,   101,   121,    45,    21,  -131,   -74,  -177,   -40,  -117,    11,   -30,   -91,   -59,     1,    73,    71,   -19,    32,     8,   -23,  -106,  -109,   -30,    86,    59,    11,    82,   -26,    60,    94,    21,    -4,   -91,   -33,  -224,  -120,  -130,    -4,    -5,  -130,    11,   -82,    23,   -69,   -34,    -3,    28,   -37,   -69,   -19,   -46,    61,    19,    14,    31,   -51,     5,    27,   -44,  -181,  -212,   -66,  -271,  -160,   -91,    46,     5,  -154,   114,   -72,   -66,   -14,    -1,  -115,   -55,   -68,   -92,  -142,   -19,   -60,   -36,    50,    29,  -118,    22,     9,   -91,   -61,   -69,   -91,  -213,  -137,   -61,    13,   -32,  -132,    55,   -14,   -70,   -97,   -37,  -123,   -48,     1,   -34,   -22,   -69,    -4,   -71,    39,   -39,   -25,    15,   -14,   -81,    -1,    73,   -43,  -141,  -103,   -40,     9,   -41,  -252,    20,   -93,    27,    -8,  -163,   -45,   -78,   -46,   -52,  -103,   -73,   -51,   -75,    16,    15,   -50,    17,   -67,  -102,     3,   140,   126,    60,   -75,     3,    16,   -12,  -213,    29,   -35,    42,    36,   -38,   -55,  -109,    27,   -20,   -76,   -52,   -10,   -41,    83,    70,   -18,   -73,  -114,   -16,    31,   102,    91,   -15,  -206,     8,     7,    -1,  -163,    60,   -59,    -7,   -45,   -67,    -4,   -52,     0,   -89,    32,   -44,    77,    15,    96,    88,    10,   -73,   -37,    18,   124,   126,    99,  -148,  -148,    -8,    -1,    10,   -23,    33,   -56,    10,    19,   119,    51,     3,   -45,   -14,    10,    44,   102,    83,    65,    46,    37,    -3,   -33,   -14,    47,    99,   152,   -69,  -102,    10,   -19,    -3,   -75,  -107,   -38,    50,   140,   176,   109,    77,    29,    60,    24,    45,   -92,   -57,   -69,    43,   174,    83,    91,    16,   -71,    20,    31,   -70,    -7,    -8,    -8,     2,    77,   -92,   -16,    69,   120,   158,   108,   101,     3,    41,   -26,   -69,    53,   -28,   -15,   114,    92,    45,    80,   -37,   -15,   -59,     2,     5,   -29,     9,    -5,   -16,     3,    70,     5,    42,    82,   145,   -33,    39,    -4,   -55,    46,   -39,   107,    99,    43,     5,    49,   -18,   146,    34,   -46,    90,    37,    -3,    17,    -2,    11,     9,    -9,    13,    -3,   -71,    29,    20,    28,    -3,    37,    56,    70,    41,    54,    19,    54,   -85,     1,    30,   -48,  -116,   -85,   -76,     9,    -9,    20,   -16),
		    70 => (    4,   -13,    -8,     7,    18,    -9,   -13,     4,    -5,    17,    -1,   -10,    -1,     0,   -14,   -13,    12,   -19,     5,     6,   -14,    17,     1,    -9,    20,    -3,    -7,    -3,    13,    19,    19,     1,     1,     2,     1,    -5,    12,   -19,   -12,    -1,    15,    39,   -23,     8,   -15,    10,    11,     2,     2,    -5,    15,    18,    -1,     3,     6,     5,    -5,    -1,     8,   -12,   -12,   -16,   -22,     9,   -30,   -33,    -2,   -35,   -46,   -79,   -32,    17,   -38,   -57,   -26,   -17,     0,   -20,    -5,   -21,   -11,    10,   -20,    -6,   -18,    19,   -18,   -18,   -10,    26,   -37,   -42,   -42,  -155,   -85,   -53,    10,    56,    29,   -84,   -18,   -14,     2,    10,   -36,   -86,   -84,   -39,    15,     8,    -7,   -16,    12,    16,    20,     9,   -31,  -138,   -43,    -9,   -50,   -18,   -30,    83,   112,   127,    60,    35,  -106,  -127,   -33,    19,  -100,  -114,   -57,   -36,   -35,   -67,   -37,     0,   -12,    -9,   -40,   -14,   -27,   -90,   -30,     7,    11,    -3,    15,    39,   135,    36,    36,    63,   -25,  -118,   -90,    59,   -61,  -119,     8,    25,    -7,   -95,   -78,   -50,    18,   -22,   -12,   -28,    25,    36,    49,    46,    53,    15,     1,   115,    16,   -17,    14,     3,    78,    51,   -60,     1,   -44,   -27,   -15,   -27,   -20,  -141,   -71,   -29,     0,   -13,   -32,   -76,    14,    50,    73,    59,    21,    50,    11,    59,   -10,    17,    92,    53,   106,    33,    28,    42,    57,    37,   -73,   -28,   -29,   -30,   -79,   -61,    18,   -16,    73,   -62,    55,     5,    42,   -47,    -8,    76,    60,   -20,   -47,    76,    59,   -20,   -56,   -60,    73,     5,    27,    72,   -15,     4,   -62,   -46,  -118,   -49,    17,    -4,   101,   -14,   -21,   -45,   -81,   -73,    56,    66,    82,   -13,   -28,    74,   -10,     9,   -40,   -11,   -35,    90,   -17,   -43,   -30,   -45,   -82,   -79,   -96,    16,    -4,    16,    95,    23,   -56,   -13,   -63,   -76,    48,    45,   -10,    -2,     3,   -84,   -24,    53,     7,   -45,   -78,   -67,   -89,   -50,   -46,    49,   -20,   -36,   -74,     7,     9,   102,     4,   -51,   -69,   -15,   -33,   -49,   -11,   -19,    43,   -49,  -151,  -227,  -171,   -27,   -54,   -78,   -79,   -84,   -34,   -46,   -33,   -32,    40,   -47,   -34,   -45,     8,     1,   -14,   -30,   -71,   -90,   -40,   -86,   -43,   -16,   -63,    -7,  -184,  -222,  -261,  -119,    62,   -41,   -58,   -24,    15,    12,   -14,   -41,   -96,   -70,   -68,   -47,    -4,    17,    27,    63,   -29,    -1,    13,   -53,   -39,    23,    27,     3,  -136,  -224,  -100,   -49,     2,    38,   -26,   -46,    30,    63,   -23,   -27,   -81,   -62,   -96,   -24,     2,     9,   -19,    57,    36,    -8,   -46,   -41,   -73,    51,   114,    -3,  -130,   -98,   -76,   -92,  -111,   -15,    25,    -6,    14,    57,    18,   -31,   -54,    -8,   -87,   -19,    -1,     3,   -26,    34,    59,    18,  -123,   -45,    18,    89,   147,     5,   -64,  -116,   -36,   -89,  -190,   -13,   -12,   -23,    71,    40,    71,   -52,   -68,    65,   -70,   -77,   -10,     4,   -13,    38,    39,   -63,   -92,   -51,   -13,    33,    71,    69,   -88,   -52,   -71,   -50,  -237,   -11,   -36,   -31,    58,   -32,    46,   -45,  -103,   -41,  -163,   -41,    -2,   -20,   -47,    25,    21,   -47,   -82,   -24,    -8,    38,    71,    21,   -24,  -122,  -168,  -304,  -127,    -7,   -73,   -26,    31,   -43,     4,     7,   -38,   -61,  -122,     5,     6,    -7,   -40,    -8,   -15,   -74,   -89,   -65,   -56,    38,    82,    23,   -41,  -107,  -226,  -241,  -162,   -88,    88,    -1,    60,   -33,   -10,    -2,   -55,   -61,   -83,   -28,   -16,    21,   -38,   -20,   -19,   -32,   -97,   -62,   -31,   105,    39,   -30,    18,   -51,  -104,   -75,   -39,   -27,     4,   -10,    40,    -9,   -58,    15,    13,  -153,   -34,     1,    15,    15,    -9,   -45,    36,    73,  -111,   -64,   -58,     6,    44,    89,   -71,   -25,    87,     3,   -36,   -22,    15,   -50,     8,    29,   -65,    44,    15,  -118,    47,    17,    -9,    15,    -4,   -18,   -24,    -5,  -146,   -31,   -72,   -45,    12,    56,    77,    76,    53,    68,   -68,   -49,   -25,    14,    57,    11,     8,    27,    27,   -16,    39,    55,     2,     0,    -5,   -26,   -47,   -22,   -63,   -31,   -34,    -2,   -45,    60,   -10,    44,    59,   -13,    30,   -33,     5,    46,    65,    32,    18,    38,   -17,     8,    40,    34,    -3,     8,   -14,   -55,     6,   -21,   -94,  -131,   -44,    50,   -16,   -38,   -20,    72,    48,    96,   133,   134,    34,   -72,   -62,   -29,   -17,   -51,    18,   -77,   -32,     4,    -4,   -14,   -30,     8,    50,   -27,   -65,   -56,   -92,   -40,   -35,   -47,   -36,   -30,   -48,    -1,    -9,    20,   -11,   -64,   -29,     6,     4,   -34,   -26,   -10,     9,     0,    11,    18,    16,   -10,   -22,    -3,   -40,    -8,   -19,   -12,   -14,   -29,   -23,   -35,    -7,  -145,  -106,  -117,   -61,   -81,   -97,   -65,   -58,   -13,   -19,    16,     5,    -6,     4,   -16,    13,    -5,     1,   -54,   -81,    -8,   -19,    -4,   -36,   -29,   -21,   -73,   -94,   -77,   -70,  -116,  -122,   -24,  -105,   -76,   -17,   -13,   -20,   -18,    -1,    15,     2,    19,   -18,    -6,    18,    11,   -10,     9,   -17,   -17,   -19,   -22,     6,   -40,   -22,   -13,   -15,   -14,   -17,    -2,   -12,   -38,   -29,   -20,   -11,     5,    -5,    -8),
		    71 => (  -10,   -19,   -17,   -13,    -9,    -6,     6,     1,     5,   -19,    -8,    10,     7,   -12,    14,    10,    10,     8,    18,     3,   -18,     3,   -10,   -19,   -12,    16,   -19,    17,   -11,   -11,     7,    12,     8,     8,    12,    13,   -20,     7,   -11,     9,   -11,    -9,    53,    18,    39,    -1,   -25,   -15,   -17,    12,   -12,   -18,    -5,    10,   -16,     7,   -12,    17,   -10,    -9,   -15,    12,    10,    13,   -62,   -70,   -39,   -35,   -90,   -49,   -69,    -1,    90,    -8,   -26,   -22,   -59,  -147,  -101,   -70,   -26,   -33,     1,   -11,    12,   -13,   106,     9,     4,   -32,   -34,   -12,   -66,   -96,  -107,  -134,   -10,    14,  -132,   -37,    64,    71,    74,    66,    74,    83,   -33,    -7,   -23,    -7,    -7,    18,     9,   -12,    85,    88,    24,    37,     9,    -9,    34,    -2,    31,   -12,    -6,    40,   -72,  -101,   -12,    27,    49,    81,   -46,    66,   -35,    14,   -19,   -64,   -87,   -35,    18,    10,    48,    16,    24,    41,    -5,   -18,   -64,   -43,   -43,     7,    72,     4,    58,    64,    25,   -90,    -9,    50,    38,    37,    27,    18,   -21,   -70,   -17,   -40,    -7,    -3,   -60,   -57,   -20,    29,    14,   -13,  -171,  -251,  -109,     9,   -25,   -48,   -34,   -20,     9,  -100,    65,   -16,    15,    62,    39,    16,    -8,     4,   -43,   -23,    10,   -14,   -74,   -68,   -84,    33,    36,   -82,  -160,   -75,     1,   -61,   -19,   -71,   -15,   -83,   -54,   -42,    39,    21,    45,    98,    32,   -22,   -39,     7,   -82,   -17,    -8,   -29,  -103,   -74,  -107,   -32,   112,    21,  -128,   -58,    13,   -24,    78,    73,     7,   -27,   -50,   -65,   -92,  -118,     7,    51,    68,   -40,   -64,   -10,   -86,    -4,    -5,    -1,   -55,   -86,   -65,    -9,    15,    67,    44,    11,   -83,   -43,   -37,    45,    13,    -8,   -71,   -64,  -113,  -160,   -64,   -23,    28,    72,   -30,   100,    78,   -34,   -11,   -30,   -63,   -39,   -47,   -52,   -82,   -47,    57,   -38,   -97,   -31,    15,    82,    21,   -77,   -25,     9,   -81,   -42,  -109,  -132,    57,    65,   -46,    81,    67,    70,    -4,    -3,   -24,   -22,   -45,   -52,   -81,   -78,  -108,  -128,  -107,    -7,    22,     1,   -34,   -82,   -67,     5,   -94,   -77,   -44,   -59,    50,    66,   -39,    73,    44,   118,    17,    16,   -29,   -40,     4,   -14,    -3,    -2,   -81,   -42,   -17,    14,    69,    66,   -17,   -30,    12,    91,  -112,  -105,   -39,   -37,   -49,   -22,    -2,   102,   125,   149,   -12,     9,    -7,     2,    -8,    44,    31,    16,    71,    75,   -34,   -27,   -24,  -109,    -6,   -20,    17,    21,  -149,  -141,   -92,   -81,   -90,  -138,   -87,   131,   104,    -9,    18,   -13,     6,    26,   -27,    46,    49,   -25,   150,   133,    47,   -84,  -124,  -100,    17,   -18,    72,    -8,   -67,  -118,   -47,   -72,   -60,   -26,   -11,    -9,    11,     1,    -4,   -12,     6,   -32,   -49,   -37,   -79,    41,    60,   137,     4,   -45,   -35,   -12,   -16,   -11,    44,   -13,   -29,   -89,   -87,  -105,   -77,   -75,   -97,    -9,    -5,   -35,     6,     8,     7,   -48,    -6,    34,   -73,    -5,    58,    32,    24,   -81,   -10,   -21,    18,   -98,     0,   -40,   -79,  -158,  -105,  -156,   -97,   -79,    -6,  -101,   -56,   -18,    18,    -5,    -7,   -51,    -2,    34,   -40,  -102,   -30,   -75,   -98,  -178,    25,    71,    19,   -12,     4,   -76,  -151,  -124,   -56,  -100,   -76,   -40,   -26,   -56,   -69,  -106,    38,    -7,   -30,   -12,   -86,   -72,  -113,  -135,  -141,  -229,  -177,  -196,   -85,   -20,    83,    15,    11,   -44,  -133,   -71,   -63,   -54,   -54,   -57,   -84,   -41,   -70,   -29,     3,   -13,    13,   -57,   -65,  -167,   -65,  -116,   -46,  -124,  -142,  -194,  -128,   -93,    90,    70,     7,   -16,   -73,   -30,   -78,   -55,    -6,    14,   -33,   -30,   -46,    -3,   -10,     7,   -27,    30,    54,   -27,    28,   -39,   -55,    47,    45,     3,    21,  -105,    99,    72,    70,    46,   132,    18,    69,   -67,   -83,   -13,    30,   -49,   -35,    -7,    31,     0,   -45,    69,    96,    54,    85,    75,    -9,   -42,    14,   -32,   -84,   -69,    40,    46,    97,     6,   103,    34,    92,    26,  -130,   -73,   -39,   -15,   -69,     1,    34,    30,  -135,   -67,   124,   167,   102,    54,    16,   -58,   -93,   -53,     2,   -44,   -25,   160,    63,   -46,    25,    11,    41,    15,   -68,   -76,   -53,   -11,     4,    -4,    16,    19,   -27,   -58,    21,     7,    64,   -81,  -117,   -48,  -131,  -100,    19,   -10,     2,    35,    15,     4,    16,   -24,    12,   -53,    -2,   -30,   -38,   -85,   108,    -9,    11,     8,     0,   -31,     7,    -7,   -27,   -28,   -75,    77,    67,    14,   -34,  -135,  -121,    29,   -25,    46,   -80,  -207,   -95,   -71,  -107,   -75,  -101,   128,   139,    18,   -12,     5,   -17,   -23,    -5,   -17,   -41,   -21,   -24,   -47,   -60,  -111,   -87,  -178,   -82,  -133,  -100,  -197,  -136,   -97,  -145,   -43,   -29,   -33,     0,   -19,   -31,     1,     0,    -1,    -3,   -11,   -17,   -28,    -9,   -38,   -10,   -43,    -4,    -1,  -136,  -100,    46,    28,    83,  -133,   -43,   -35,    -2,   -30,    -3,     6,    19,    -1,    18,    19,   -11,    -5,    -2,    -2,    19,    18,   -13,    -1,   -18,    19,   -42,   -34,   -20,   -26,   -50,   -45,   -34,    -4,    16,    13,   -17,    14,    -5,     4,     6,     1,   -14,    12),
		    72 => (  -15,    -6,    -3,   -20,    -6,    19,   -10,     9,    10,    -3,    12,    11,   -44,   -43,    28,    16,    14,    20,   -18,    13,    -5,    16,    -2,    13,   -11,     7,    -7,    -3,    -9,    -1,     3,     3,     3,    10,   -23,     1,   -87,   -54,   -86,  -110,   -77,  -108,   -52,   -74,   -26,   -53,   -74,  -159,  -113,   -36,   -28,   -34,    18,     3,     5,    11,   -13,    -1,   -26,   -22,   -67,    -8,   -10,  -104,   -37,    93,    82,   -11,   -25,  -163,  -132,  -214,  -147,   -37,     3,   -33,  -181,   -51,   -63,   -26,    42,    17,   -11,    17,     1,     9,   -28,   -78,   -37,    19,     7,    -2,    36,    35,    60,    -3,   -88,  -198,  -150,  -169,  -166,  -136,  -150,  -132,  -149,  -111,   -71,   -30,     6,     6,    19,     8,    11,   -18,   -56,    -9,    11,   -40,    50,    45,    14,   -29,    67,    12,   -60,  -174,  -152,  -126,  -145,   -88,  -141,  -138,   -90,  -104,   -69,   -60,     5,   -14,   -65,   -26,   -17,    14,   -38,    -1,    43,   -59,    89,    82,    91,     7,    52,   -49,    40,    -2,   -67,   -12,  -175,  -176,  -126,   -77,   -45,   -89,  -115,   -38,   -67,   -21,   -12,   -35,   -17,     5,   -12,    14,    37,   100,    66,    18,    57,    70,     0,   -20,   -16,    49,   -15,   -77,   -88,   -92,   -92,   -45,   -38,   -89,   -86,   -69,  -109,   -38,   -32,   -30,    -2,    -8,    -6,   -39,   -17,   -15,   -71,   -38,     7,    23,   -85,    -9,   -24,   -21,   -57,   -64,   -85,   -23,   -93,  -109,   -99,  -132,  -144,  -158,  -113,   -69,   -64,   -40,   -64,   119,   -25,     2,  -111,   -31,    27,   -29,     8,   -41,    41,   -37,   -49,    56,    57,    11,   -34,   -32,   -71,   -84,  -166,  -173,  -141,  -137,  -155,   -65,   -88,   -41,   -17,   -56,   -35,    37,  -129,   -20,     6,   -44,    -3,    -9,    29,    10,    25,    11,   165,    47,   -24,   -73,   -97,   -80,  -107,  -101,  -208,   -52,   134,  -116,   -39,   -51,     0,   -43,   -33,   -17,  -153,    53,    -8,    -4,    -2,   -61,   -69,   -34,    20,   -26,    38,   103,    80,   -59,   -92,   -57,   -60,  -105,  -105,    21,    80,   -59,   -86,   -76,    -2,   -11,  -112,   -45,   -58,   -45,   -46,   -30,   -49,     2,    27,   112,   -63,  -100,   -21,    32,     9,   -26,   -17,   -83,  -100,  -145,   -81,    10,   -18,   -84,  -154,   -17,   -14,   -20,  -133,   -18,   -12,    35,   -85,  -152,   -19,   -51,   -79,   -50,   -11,    -6,   -42,   -18,    43,   -22,   -12,  -104,   -82,   -28,    21,  -133,   -36,   -46,   -70,    13,   -14,   -20,  -103,    -5,   -22,   -32,  -120,  -161,   -37,   -63,  -114,   -66,   -40,     6,   -50,    40,    10,    19,   -51,   -60,    32,    95,   124,    21,   -35,   -23,    81,    78,    10,    -9,   -23,   -32,   -89,    -9,  -139,   -98,   -40,   -90,   -31,   -42,    -2,    29,    20,    32,    46,    -5,   -56,     1,    39,   100,    58,   -15,   -32,     4,   161,    79,    -4,   -28,    87,   -69,   -20,   -12,   -22,   -79,   -48,   -15,    21,     3,    72,   110,    39,    51,    -2,   -24,   -22,     6,    54,    12,   -53,   -82,    -2,    28,    44,    98,    11,     4,    94,   -21,    54,   -70,    10,   -22,  -129,   -31,    25,    73,    10,    55,    47,    43,    88,    49,    10,    42,    -7,    41,    36,    43,    30,    55,   -22,    94,   -19,    -6,   139,    21,    74,   -39,    71,     8,   -33,    15,    50,    61,    -9,    13,    70,    63,    74,    52,    72,   105,    65,    80,   -30,    20,    -5,   -41,  -105,    87,   -10,     9,    60,    49,    41,    32,   107,   -11,   -58,    17,    57,    63,   -44,    24,   -32,    50,    29,    12,    63,    37,    18,    64,    51,    75,   124,    65,   -76,    61,     2,   -71,    10,   110,   -15,    68,    47,    28,    -8,    81,    21,   -18,   -62,   -47,   -23,    58,    -6,    -5,   -36,   -52,   -54,     1,    72,   123,    73,    38,    69,   142,    -8,   -34,    22,    81,    10,   -23,    16,   -36,    40,   -14,     2,   -11,   -17,     8,    20,    -4,   -99,  -143,  -123,  -118,  -106,   -29,   -55,   -29,   -32,  -101,    56,    -9,    17,    -6,   -15,    46,    34,    25,   122,     3,    -5,   -14,    72,   -63,    24,   -45,   -57,   -60,  -187,  -281,   -37,   -55,   -94,  -113,  -122,  -165,  -165,   -83,   -75,    -3,    20,    12,    -7,    -8,    -6,    41,    24,   -53,   -57,   -63,   -85,   -34,   -39,   -78,   -66,  -174,  -270,  -250,   -75,   -44,   -99,  -150,  -184,  -136,  -134,  -113,  -180,    -2,    13,   -20,    17,   -18,   -25,   -38,   -48,   -82,    -4,    -5,  -118,  -127,  -231,  -198,  -262,  -211,  -247,  -237,  -164,  -175,  -163,  -175,  -153,  -212,  -165,   -94,  -169,    17,    -2,    15,   -53,   -17,  -189,   -52,  -119,   -33,    15,   -87,    13,   -55,  -359,  -256,  -225,  -187,  -212,  -234,  -199,  -192,  -182,  -193,  -149,  -150,    26,    64,    58,     1,    -8,     2,    -7,    10,   -49,   -34,    -9,   -27,  -142,  -190,  -206,  -128,  -202,  -188,  -132,  -161,  -165,  -125,   -96,  -163,  -168,  -141,   -38,   -41,    -1,    34,    41,     7,    -3,   -14,   -18,     9,     0,   -61,  -102,   -98,  -145,  -181,  -133,   -46,   -55,   -63,   -95,   -36,   -77,   -65,   -35,  -115,   -59,   -40,   -73,   -16,   -15,     2,     4,   -11,   -12,     4,     8,   -15,    -2,   -12,   -19,    -5,    15,   -26,   -46,    -9,   -26,   -69,   -40,    -8,   -35,   -31,   -57,   -33,   -43,   -45,   -41,   -15,    20,    19,    -4,     0),
		    73 => (   17,     2,   -17,    10,   -18,    13,    -7,   -14,   -14,     3,     9,    18,   -24,   -13,   -31,     1,    -6,    15,   -14,   -20,    11,     9,     2,     6,    10,   -19,    -5,     1,   -10,    12,    12,    -5,     2,    -2,   -12,     4,     2,     3,   -21,   -21,   -15,   -28,   -52,   -42,   -28,   -22,    -6,     9,     1,     5,    10,     1,   -12,    -8,    18,    -2,   -11,    -4,   -12,    -4,    -6,    10,     6,   -22,   -32,   -56,  -159,  -156,  -155,   -30,   -32,    -5,   -23,   -23,    12,    -1,   -48,   -11,     1,   -34,   -18,    -4,    -6,    -1,   -13,    -1,    -4,    -3,    -1,   -32,   -20,    -5,    23,     4,   -24,   -90,   -54,   -82,  -113,  -125,  -116,   -48,   -37,   -20,   -32,   -42,   -62,   -82,     2,    -1,   -18,     3,   -11,    -4,    16,    10,     1,   -13,   -33,  -114,   -86,  -207,    26,    72,   -16,   -16,    66,    17,     0,   -14,    -9,    -2,   -20,    63,   127,   -84,   -89,   -75,   -10,     2,    -7,     0,    13,   -13,     5,   -67,   -48,   -67,  -154,  -162,   -60,    71,    57,   -73,   -34,   -40,     1,   -52,   -41,   -62,     7,   -76,   -28,   -58,   -52,  -186,   -58,   -15,     0,     7,    40,    29,    -2,   -57,    21,   -34,   -22,    44,   104,    26,   -15,    37,   -23,    26,    36,   -77,   -33,   -93,     9,     0,   -58,   -10,   -44,   -89,  -130,   -41,    19,    17,    13,    -7,    16,  -183,  -146,   -66,    18,    11,    -5,   -82,    24,   129,     8,   -54,   -66,   -22,     3,   -26,   -30,   -57,   -35,   -92,  -135,   -82,  -101,   -13,    -2,   -10,   -13,   -31,     0,  -129,   -90,    10,    19,    18,   -39,   -29,    64,    54,   -14,   -36,    13,   -38,   -29,   -13,   -18,   -22,    -2,   -51,  -239,   -72,  -160,    19,   -19,   -27,    13,   -34,   -76,   -72,   -31,    44,   -15,    21,    47,    95,    62,   -23,   -22,   -54,    30,    54,   -38,    11,    21,   -18,    30,    19,  -192,   -70,   -92,   -79,     5,   -46,   -10,   -22,   -41,   -75,   -28,   -75,    36,     9,    32,   100,    57,   -91,  -109,   -41,   -53,   -37,   -63,    25,    84,   -66,    21,    -8,  -182,  -154,  -139,   -63,   -16,   -61,     0,    40,    92,    60,    26,     1,    89,    14,   -91,  -105,  -353,  -136,   -55,   -71,   -53,   -17,   -51,    18,    55,   103,   -11,    49,  -149,  -102,   -66,    14,    -6,   -38,   159,    29,   112,    72,     6,  -127,  -105,  -173,  -174,  -240,  -181,   -21,     7,   -36,   -34,   -71,   -44,   -14,    30,    74,    63,    54,   -99,    24,   -51,     0,   -10,   -62,   -76,   -97,  -108,   -90,   -74,  -272,  -241,  -183,   -99,   -59,    14,    98,    94,   -59,     9,   -14,   -30,     6,   -16,   -30,   -34,   -16,  -109,   -71,   -90,   -29,    -1,    21,    50,   -42,   -76,  -209,  -203,  -237,   -28,    68,    35,   -37,    -2,    53,    -6,    23,   -18,    48,     3,   -74,   -94,   -51,   -52,    10,   -62,  -146,   -89,   -29,   -19,     6,     2,   -21,  -106,  -223,  -290,   101,    97,    15,    24,    42,    84,    81,    72,    20,   -14,   -13,    13,   -20,  -115,   -71,  -135,   -58,   -63,   -84,    88,   -23,   -11,    16,    43,   -34,   -44,   -78,   -31,   -35,    51,    74,    75,    84,    70,    55,    66,   -18,    -6,   -47,   -14,   -56,  -133,   -90,   -84,    13,   -40,   -53,   -26,   -29,    15,    16,    38,    30,   -98,  -101,   -49,   -71,   -26,    33,   114,    42,   115,   103,    24,  -106,   -74,     4,   -27,    -7,  -133,   -94,   -67,   -47,  -149,   -55,   -17,   -11,   -37,   -24,    10,    39,   -92,  -173,  -190,   -59,   -93,    -6,    43,    78,   105,    16,     5,   -44,   -48,   -85,    35,   -13,    17,   -49,   -51,  -128,  -152,   -26,   -16,   -14,   -18,   -50,     7,   -10,  -146,  -135,  -161,  -144,  -192,  -138,  -172,   -67,  -125,   -46,   -88,   -45,    63,    39,    80,    12,   -68,    28,   -67,  -135,  -150,    -7,   -73,   -22,    11,   -48,    28,   102,   -38,   -13,  -151,  -245,  -258,  -387,  -512,  -379,  -300,  -107,   -14,   -49,   -14,    68,    95,    57,    22,   -36,   -67,  -178,  -141,   -93,   -24,    17,   -25,   -16,    75,   163,   100,    -1,   -14,   -98,   -20,   -77,   -80,  -121,   -82,   -61,     4,    36,    -6,    -3,    50,     0,    48,   -18,   -49,  -121,   -90,   -35,   -45,    18,   -13,     7,    20,    90,   168,   158,   114,    71,    64,    38,    87,    37,   -34,    21,    21,    22,    42,   -15,   -25,    -8,   -48,   -34,   -87,   -57,   -95,   -55,    -7,     0,    12,    16,    17,   -39,   114,   113,   100,    86,    18,   -28,    43,    -3,    64,   113,    -4,    57,  -116,    20,   -11,   -78,    54,    16,   -30,   -27,  -102,   -63,   -11,    19,   -13,   -10,    23,    72,   146,   -25,    76,    62,     8,    11,    56,    65,    42,    50,   -10,   -22,   -43,    29,  -206,   -57,    42,    52,    74,    77,  -126,   -36,   -51,     3,    14,    -9,    21,   -79,     2,   216,   140,   118,    50,    68,    10,   -31,    13,   -30,   -78,   -34,   -29,   -78,  -211,   -44,   -61,  -132,   -51,  -160,   -97,   -53,   -70,    17,     8,    17,     0,   -64,  -125,    -3,    12,   -27,   -26,  -103,    -1,    12,   -38,    17,     0,  -107,   -14,    47,    37,   -52,   -27,   -43,    16,   -13,   -16,    -6,    10,    -2,    19,   -13,   -18,    -2,   -13,   -46,   -16,   -12,   -14,  -118,  -105,   -83,   -57,   -71,   -74,   -76,     6,   -12,   -37,   -85,   -76,   -15,   -65,     3,   -17,    -8,    -1,    -5),
		    74 => (   -6,    -3,   -19,     2,     3,    16,    -6,    10,    19,    13,    12,    18,   -15,   -63,   -13,    -4,   -17,    -4,   -20,    19,   -12,   -15,    -6,     8,    -5,    20,   -11,    -5,     1,    -3,    20,   -15,    17,    16,   -76,   -74,   -27,   -67,  -121,   -69,  -145,   -87,    37,  -220,  -196,  -139,   -40,    -7,   -92,   -16,     0,   -32,   -18,     8,    10,   -13,    -5,   -12,   -32,   -84,  -123,   -84,   -41,  -113,   -70,   -71,  -191,  -248,  -190,   -44,    27,   -61,  -111,   -91,  -127,  -167,  -170,  -108,  -112,  -135,   -35,   -82,    14,   -19,   -16,    -4,   -52,  -155,  -254,   -86,   -98,   -10,  -174,  -199,  -120,  -168,  -287,   -96,    29,   -19,   -75,  -112,  -153,   -50,   -38,   -80,   -49,  -142,  -166,   -68,    -7,     8,    -1,     0,   -28,  -221,   -24,     8,    12,    34,   -10,  -115,   -85,   -80,   -22,    58,    71,    32,    18,    50,    81,     2,   -43,    17,   165,     7,   -18,   -33,  -150,   -44,   -12,     9,   -55,  -102,    19,    47,    32,   134,    73,    56,    53,   -23,    49,    83,   127,    31,    -8,    93,    33,   113,   -22,    73,    73,   124,   126,    70,  -143,     1,   -14,     8,   -47,   -29,    85,    57,    21,   139,   115,   125,    75,    44,    24,   127,   159,   208,   125,    27,   -57,    -1,    52,     6,   -13,   122,   160,    46,    33,   -85,    -2,   -82,   -70,    41,    90,    42,    86,   144,    64,   297,   190,   263,   144,   160,   146,   135,    79,    93,    31,   104,    44,   -44,   -31,    14,    64,   -64,   169,  -117,   -85,   -97,   103,    47,    48,     8,   112,    60,    -8,   249,   143,   162,    25,   -32,   -13,    40,   -48,   -49,   -47,   -18,    23,    16,  -112,   -39,    -1,    43,    78,  -128,     9,   -38,    82,   -67,    12,   -61,   -86,   -40,   -39,    -5,    44,  -107,   -40,    17,   -33,    18,   -78,    39,   -18,   -27,   -25,   -30,  -135,     0,   -28,   -79,   -77,   -68,    14,   -51,    45,   -44,   -42,   -94,  -164,   -72,   -77,    22,   -44,  -127,     0,  -102,   -87,   -45,   -42,    -6,  -104,    -1,  -130,   -69,   -32,   -81,  -176,   -50,   -12,  -102,    20,   -86,    45,   -67,   -85,   -69,    59,  -122,    16,   -53,  -110,   -34,   -14,   -36,   -61,   -21,    13,    69,   -89,   -79,  -214,   -87,   -59,  -130,  -212,   -52,   -86,  -165,   -14,    20,    16,   -69,  -116,   -34,   -14,   -81,   -15,    13,   -62,    35,   125,    62,  -118,     3,    24,    50,   -29,   -53,    -2,    64,   -29,   -84,    17,   101,   -80,  -136,    -5,   -39,  -114,  -105,  -117,   -13,     9,   117,    67,   -52,    37,   114,   144,   -15,    39,    20,    -1,    58,    69,   -19,     6,   -63,   -76,   -35,    12,    57,   -40,   -17,   -19,    65,  -201,  -137,    -3,    -4,    -4,   185,   105,    60,   105,    75,    48,   -32,   -42,   -16,    26,    24,   -35,   -17,   -85,  -105,   -25,   -18,    -5,    80,  -110,   -15,   -20,    17,    87,    20,   101,    -7,    68,    89,   106,    53,    18,    19,    93,    63,    20,   -10,    47,    96,   -26,   -46,     6,     9,    92,    55,   -39,   -11,   -72,  -111,    12,     4,  -125,    28,   -52,   -52,   -46,   -39,     4,    -6,    56,    55,     7,    -3,    22,   -14,    32,    41,    21,    44,    97,    67,    69,   -16,    43,    19,   -66,   -46,     5,    -9,   -80,  -104,     2,     7,   -57,    94,    16,   -20,  -107,   -43,    10,   -73,   -20,   -73,    80,   -18,   -33,    25,     4,    72,    29,   133,    40,  -158,   -28,   -53,   -85,   -17,   -29,     4,    14,    75,    41,    12,   -88,   -36,  -105,   -75,    40,   -48,    10,   -48,   -61,  -125,   -38,   100,   167,   103,    63,   114,    75,   -42,   -71,  -101,     6,   -76,  -112,   223,   -57,   -38,   -62,  -111,   -44,   -97,  -119,  -121,   -11,     8,    37,    54,    23,  -129,    -3,    50,    56,    41,    72,    11,    24,   -10,   -29,   -81,    14,   -24,   -58,    54,   -71,  -108,  -120,  -130,   -69,    52,     9,    12,     1,   -19,     6,    45,    71,   -18,    82,    76,   119,    76,    31,   -24,  -118,  -136,   -59,   -16,   -33,   -11,   -84,    70,    52,   -48,   -79,   -65,    20,    31,    -1,    37,   -86,   -42,   -26,    51,    59,    49,   -16,   101,   222,   170,   176,    53,   -41,  -190,  -127,     6,   -32,   -30,   -35,  -107,  -232,  -123,    -1,    41,    97,   -40,   119,    14,   -23,    -4,   -87,   -51,    89,    83,    -4,   168,   194,   213,   135,   111,     9,    -4,   -36,   -25,    19,    13,    -6,  -153,  -199,  -369,    65,   101,   156,   100,   177,   133,    55,     4,   -30,   -53,    32,   -13,    79,   183,   179,    77,   -75,    79,    -2,   115,   -36,    -3,     4,    11,     8,   -57,  -193,   -33,   153,   167,    46,   120,    19,   139,   -44,    -7,    -7,  -126,   -59,   -70,    95,   164,    -2,   -55,   -28,   -11,  -101,    96,   -95,    -9,     2,    -3,   -60,    -5,   162,   224,    74,   -60,   -43,    20,    84,    73,   -80,    45,  -104,    34,    14,   -23,   -26,   -19,   -26,   -39,   -36,    20,   -40,  -107,   -79,    18,     6,   -19,     1,  -144,   248,   210,   122,   -42,   -88,  -142,  -246,   -49,   -72,   -80,   -47,  -181,  -191,  -127,   -32,   -11,  -146,  -293,  -259,   -67,    14,   -17,    20,    12,     0,   -20,    10,    -8,   -30,    -5,   -85,   -95,   -63,   -75,  -101,  -123,  -100,   -34,   -74,   -31,  -157,  -232,  -185,  -110,  -119,   -54,   -84,     9,    20,     3,     0,     1),
		    75 => (  -14,    15,   -16,    -5,     0,    -6,   -13,    10,    -8,   -17,     3,    -3,    14,     7,     5,   -16,    20,     2,    13,    -3,    13,     9,    -4,    -5,    17,     7,   -13,   -13,   -11,    -1,   -16,    -4,   -17,    16,    -3,    -3,    16,    12,   -18,   -21,   -34,   -61,   -44,   -30,   -25,   -60,   -42,    -4,    -9,   -26,     7,    10,   -20,    20,   -10,     7,     5,    -6,   -16,   -16,     3,     5,   -46,   -29,   -98,  -101,  -117,  -120,   -62,   -77,  -186,   -30,    23,    22,   -16,    60,   102,     5,    -1,    28,   -50,   -10,    17,     0,     6,     4,   -21,    28,    54,   -81,   -95,   -99,   -60,   -31,   -33,   -52,    13,    30,    58,    69,    55,    -9,   -67,   -51,    20,    61,    17,    52,    25,    17,    25,    20,    12,   -12,     1,    44,     0,    -8,    52,    78,    23,    79,     4,   -98,   -59,    -7,    34,    80,    91,    10,    -6,   -62,   -18,     5,    43,    57,    42,    61,   -38,   -56,   -19,    -8,    10,    10,   -53,     2,    77,    42,    51,    10,   -19,   -76,   -89,   -18,     4,   -22,    -5,    -4,   -12,    99,    72,    -3,    63,    63,    58,    46,   -45,   -49,     7,   -19,   -84,   -56,    36,    51,   108,    33,     9,   -11,    -1,   -48,   -60,   -27,    -8,    -4,   -19,   -46,    22,   103,   110,    75,    57,    33,    57,    57,    40,    21,   -16,     9,     8,   -69,    17,   126,    17,    25,   -47,   -22,   -33,   -17,   -31,   -46,   -10,   -49,    -4,   -18,   -28,     7,    48,   -21,    60,    53,   118,    66,    49,    56,   -16,   -60,   -67,  -111,    23,     4,     5,    12,   -39,    11,     2,    52,    35,    37,    -6,   -67,   -63,   -94,    19,    26,   -32,     7,    93,   119,    57,    86,    53,    29,    -5,   -29,  -141,   -99,    10,    21,     8,     8,   -43,   -29,    45,    63,    95,    72,   -34,   -40,   -82,   -76,   -31,     3,    38,    95,   117,   112,    92,    18,    77,    23,    10,    -8,   -22,  -148,    -4,    -3,   -11,    39,   -41,    14,    -5,    93,   124,    13,    57,     3,   -91,   -32,     7,    56,   108,   162,   153,   117,   110,    56,     6,   -54,    14,   -21,   -14,   -94,    32,    -2,    21,    38,    51,   -17,   -37,    89,    72,     8,    60,   -55,   -78,  -124,    98,    85,   148,    58,    70,    73,    99,    87,    16,   -66,     7,    10,     0,  -112,    32,    51,    56,    56,    98,    67,   -58,     1,    25,     9,    15,   -29,   -83,    -9,    50,    98,    58,     2,   -21,    60,    39,    41,    94,   -69,   -19,    -1,   -13,  -122,     2,    38,    44,    83,    58,    85,   113,    50,    41,   -34,     3,   -81,   -48,   -40,     1,    84,    74,    80,    -2,   -52,   -53,    -5,    74,   -64,    16,     0,   -28,  -162,   -14,    22,    60,    72,    67,    50,   119,    14,    23,     7,    -1,   -65,   -30,    31,   112,    89,    78,    61,    47,   -44,   -76,   -74,   -52,     6,    19,   -23,   -40,   -15,    34,    57,    -5,    26,    63,    97,   113,   -11,    -9,     6,    58,    14,    -4,    44,    66,    94,    52,    48,    28,     2,    15,   -79,   -49,  -105,    -5,   -30,   -73,    -9,    39,   143,    37,    23,    59,    64,    58,   -68,    11,    22,    12,    45,   -50,    13,     4,    15,    80,   144,    66,     4,   -36,   -82,   -60,  -127,   -13,    -7,   -60,    32,    52,   136,    92,    80,   101,    90,   -31,   -39,   -65,     3,    67,   -49,    11,   -17,   -14,    -7,    59,    38,    70,    16,   -18,   -86,  -139,  -147,    -4,     5,   -88,    14,    24,   119,    90,    70,   109,    87,    -9,   -83,  -133,    36,    45,     4,    -9,   -36,   -46,   -64,   -19,     3,   -10,    35,    38,   -60,  -167,   -93,    20,   -21,    66,     7,    28,    59,    63,   123,    84,    -7,   -46,   -47,   -71,    42,     3,    17,   -44,    14,   -21,    11,    13,   -10,    -8,    57,    22,   -64,  -180,   -77,    18,   -12,    44,    37,    32,    24,    66,    83,   105,     2,   -41,   -64,    14,     7,   -42,   -28,   -21,    11,    56,    57,   -27,    28,    34,    68,   -72,   -17,  -125,    -7,     1,     3,    14,    12,    20,    58,    72,    98,    92,    72,     2,    42,    24,    19,    -2,   -22,    -4,    -7,    26,    62,    73,     8,    25,    17,   -80,    -5,   -76,   -18,   -12,    -8,   -88,   -10,    33,    18,    68,    45,   101,    58,    27,    98,    46,    13,     9,    11,   -35,   -46,   -37,    14,    24,   -48,   -32,   -44,  -108,    10,    70,   -14,     1,    -4,    22,     0,   -48,    -8,    43,    77,    50,    29,    -4,    47,    41,    43,    30,   -31,  -117,   -84,   -46,   -43,   -22,   -81,   -49,   -80,   -26,    34,    55,    10,   -20,   -14,   -23,     3,   -63,   -31,    56,    25,    22,    52,    58,    42,    20,   -29,    20,    -2,   -72,   -57,   -24,   -62,   -70,   -55,   -42,   -35,    22,  -131,   -45,     4,    13,    -5,    12,    66,  -119,   -97,   -11,    31,   -44,   -71,    70,    37,    40,    20,     0,    32,    45,    81,    60,   -16,    47,    24,    89,    26,     6,    -3,   -11,    -1,    -9,   -16,     0,   -61,   -92,  -124,  -142,   -24,    -6,   -34,   -26,    71,   -17,    22,    66,    38,    41,    13,   -32,   -17,   -64,   -48,    17,   -74,     1,    -1,    17,    -9,    -9,   -18,   -16,   -13,   -33,   -25,   -10,    -3,   -13,    -3,    16,     3,   -31,   -18,   -29,   -16,    -6,    11,   -12,   -47,   -27,  -100,   -75,   -29,   -11,    15,    12,   -10),
		    76 => (    9,    -6,    13,    -6,     1,   -10,   -20,     6,    11,    16,    -7,     6,     5,    10,    -9,   -14,     8,     5,     8,    -5,    15,   -10,     6,    -3,   -19,     7,   -13,    -3,   -10,   -17,    -9,    -4,    -7,    17,    25,    35,    60,    32,    22,    39,    35,    21,   -20,   -28,   -48,    11,    -6,    -7,   107,    44,    19,    32,    12,     7,     2,     5,     8,    -8,    23,    19,    91,    33,    -1,    65,    82,     9,   -28,     2,    -4,    20,   -46,   -25,   -28,    31,    -3,    25,    37,   135,   163,   131,   121,    57,   -15,    -8,     8,     2,   -42,   -41,    -7,     2,     6,   -14,   -12,   -10,   -28,   -19,  -123,  -117,  -119,   -63,   -78,  -100,    28,   124,   125,    80,    34,   117,   120,    10,   -95,   -14,    17,    14,   -32,     6,    43,    21,   -39,   -55,   -66,   -11,   -34,   -57,  -108,  -143,  -160,  -124,   -53,   -67,   -50,    13,    15,    98,     9,   111,    36,   -31,    60,    73,   -20,    -9,   -47,   -59,    41,    18,   -23,   -35,   -25,   -12,   -69,   -92,  -101,   -94,   -72,   -33,   -50,   -20,     0,     7,   -29,    33,    64,    99,   116,   103,   130,    75,   -17,   -11,     4,   -14,    17,    24,   -29,   -17,   -59,   -16,   -64,   -62,   -44,   -67,  -124,  -135,  -110,   -25,   -24,    29,     3,   -30,    16,    85,   115,    65,    51,   113,    13,   -11,     6,    -8,    54,    26,   -62,   -12,    -6,    41,   -91,   -94,   -84,  -149,  -101,  -152,   -50,     6,    26,   -41,   -44,    16,   -50,   -47,    32,    64,    44,   122,    -3,    -2,    -6,   -28,    67,     5,  -106,   -47,   -30,   -15,  -122,  -128,  -151,  -143,  -121,   -86,    22,    13,    38,     8,    -1,   -30,   -38,   -21,  -110,   -57,    97,   -62,    11,   -18,     2,   -52,    90,   -10,   -95,   -14,    26,   -19,  -109,  -130,  -141,  -142,   -78,    35,    43,    22,   -12,    18,   -24,   -43,   -37,   -79,  -100,   -66,   -50,   -33,   -10,   -17,    -4,   -32,    65,   -23,   -62,   -17,   -17,  -100,  -209,  -158,  -113,   -23,    -8,    44,   -37,   -52,  -104,  -133,   -26,   -35,   -73,   -82,   -68,   -57,   -48,   -62,     5,   -13,    21,   -48,    27,    16,  -107,   -96,   -87,  -203,  -121,  -114,   -52,     4,    45,    -1,   -51,  -161,  -204,  -129,  -127,   -75,   -55,   -71,  -104,   -13,   -22,   -35,   -20,   -10,   -21,   -77,    19,   -28,   -80,  -103,  -123,  -122,  -134,     8,   -43,    39,   -12,   -32,   -52,  -109,  -178,  -129,  -102,   -62,   -31,   -42,    -6,   -27,   -63,   -27,    18,    14,   -11,   -46,   -17,   -20,   -66,   -75,    -4,   -37,   -41,   -25,    34,    46,   -34,    13,     8,    -2,   -30,   -37,   -21,  -126,   -71,   -13,   -11,    -3,   -68,   -22,     4,    -1,     8,   -40,   -49,   -53,   -42,    11,    62,   -50,    17,   -30,    46,    10,    16,   -57,    30,    -2,   -19,     7,    11,   -80,  -146,  -122,   -13,     6,   -28,   -36,     3,     1,   -40,   -21,   -54,   -72,    42,    32,   -31,    19,   -39,    35,    71,    -7,   -23,   -35,   -11,    36,    11,   -52,   -91,   -97,  -128,   -55,   -35,   -22,   -21,   -57,    11,     9,   -36,   -46,    16,   -65,   -27,   -14,    19,    10,    -1,    12,    42,    27,     4,    22,   -19,   -48,    23,    12,   -77,  -118,   -69,   -30,   -48,    12,   -38,   -28,   -14,   -12,   -45,   -81,   -22,   -85,   -63,     9,    24,   -12,    92,   -45,   -34,   -87,   -59,   -44,   -57,   -80,    76,    50,    10,   -68,   -20,   -39,   -53,   -36,   -47,   -96,    14,   -14,   -15,   -12,    60,   -32,   -73,   -37,    -3,    13,    -4,   -34,   -78,   -58,    -1,    33,    -3,    -1,    89,   129,    88,    -2,   -34,   -55,   -29,    -6,   -94,   -14,    -4,   -14,    11,   -48,    43,   -43,   -54,     9,   -70,    34,   -21,   -77,   -26,  -104,     0,    60,    21,    40,   107,    79,    70,    11,   -79,   -56,   -12,     4,   -11,   -37,   -12,   -11,   -27,   -52,    55,     4,    77,    39,   -28,   -14,     4,   -35,   -36,    -1,   105,    20,   -35,   -46,    -3,    17,     0,   -41,   -65,   -61,     5,    -8,   -14,     1,    12,   -14,   -56,   -46,    24,    -6,     4,     5,    62,   -60,    37,    83,    73,    49,    35,     5,   -14,   -54,   -52,   -72,   -99,   -87,   -64,   -24,    -6,   -14,     5,   -14,    -2,    -1,   -25,     9,   -22,   -38,  -139,   -41,    65,   -27,     6,    69,   108,    44,   -74,   -81,   -39,   -92,   -69,   -78,   -78,   -19,   -20,   -58,   -40,   -58,     8,    14,   -17,   -18,     6,   -46,   -62,   -28,   -78,    46,    38,    15,    42,    67,    60,    15,   -16,   -44,   -19,  -117,   -93,   -72,    -5,   -21,    -5,     9,   -42,   -47,   -14,    10,    10,    14,    -9,    -7,   -28,   -37,   -19,   -22,   -55,   -47,   -23,   -43,   -22,   -50,   -19,   -18,    25,     1,    -5,   -56,   -19,   -28,   -22,    12,     4,   -24,     4,    -7,   -17,    18,   -15,   -15,     1,   -68,   -84,   -88,   -48,   -28,   -13,     3,     3,   -16,   -18,     8,   -24,    -6,   -18,   -21,   -61,   -22,   -17,   -35,     2,   -10,     5,   -14,    15,   -19,     1,    -8,   -13,   -34,   -31,   -24,   -19,     2,   -41,   -32,   -17,    -3,    -5,    -3,   -14,     7,     1,    10,   -42,   -17,   -30,    -1,     4,    14,   -13,    14,   -16,     8,    18,    12,    11,    17,   -16,    19,    17,    14,    12,     7,    -7,    -6,   -22,    -3,   -10,   -24,     9,    -5,   -19,   -30,     9,    -6,     2,   -16,     3,   -19),
		    77 => (    3,    -6,   -11,     9,    11,     3,   -19,    17,    -3,     4,   -12,    19,    -9,    18,    10,     6,     6,    -4,     2,   -14,   -14,   -19,    17,    11,     4,    -2,    16,     0,    11,     7,    -7,    -3,    -4,    -8,     2,    16,    11,    -4,   -27,    -4,    -8,   -14,   -22,   -69,   -88,   -56,    17,    16,    19,     1,    -2,    -1,    11,     1,    -2,    20,    10,    16,     2,   -12,     2,    14,    -5,   -21,    -5,     0,   -51,   -32,    -7,   -11,   -14,   -17,    -2,     5,   -20,    -1,    -1,    -8,     0,   -15,   -11,    -3,    -8,    14,    -7,     3,   -18,   -15,   -18,   -11,    -9,    12,   -49,   -49,   -44,   -59,   -30,   -45,    11,   -59,   -71,  -140,   -41,   -71,   -43,   -36,   -74,   -16,   -29,   -16,   -14,    17,     7,    -1,    10,   -12,   -54,   -27,   -46,  -134,  -109,   -93,  -128,  -196,  -225,  -168,  -117,  -220,  -163,  -186,  -172,  -102,  -110,   -42,  -148,   -86,   -53,   -40,   -16,   -16,   -19,    20,   -21,   -81,   -15,   105,    88,    62,   141,   136,     3,    55,    21,    45,   -32,    -4,   -20,   -76,    -4,   -44,   -81,  -165,  -168,  -123,  -160,  -135,   -40,   -16,    13,    -1,   -12,   -47,   -30,    58,    76,   107,   113,    -3,    20,    65,    98,   100,   125,    30,   107,    79,    55,    63,    75,    18,    50,    -9,   -21,   -49,     2,   -39,    -1,    15,   -27,   -14,   -45,   -36,   -52,    80,   -23,    19,   -13,    74,   121,   117,    46,    71,    46,   111,    12,    39,    60,    -7,     6,   -15,    17,   -21,   -29,   -20,   -53,    32,    -3,   -29,   -32,   -88,   -79,   -67,  -110,   -98,  -111,    -7,    13,   -32,    13,    24,   -13,    45,   -27,     4,   -72,   -41,   -88,   -83,   -81,   -31,   -56,   -64,     0,    -9,   -25,    21,     5,   -66,  -115,   -88,  -185,   -59,  -111,   -73,   -60,   -88,   -47,   -78,     8,   -89,     3,   -19,   -68,   -49,   -52,   -72,   -61,   -21,   -65,    38,    -9,   -32,   -74,   -66,    -3,   -78,     0,   -51,   -86,   -51,  -103,   -58,  -164,  -195,  -200,   -52,   -38,    16,   -30,   -45,   -11,  -138,   -35,  -112,   -75,   -37,   -77,    34,    -9,   -17,   -67,    -9,   -59,   -62,   -67,  -121,  -158,  -134,  -207,  -138,  -226,  -136,  -102,   -37,    -2,   -30,   -52,   -53,   -42,   -40,    57,    70,   -54,  -124,   -67,    56,    -3,     4,   -35,    18,    -3,   -55,   -86,  -164,  -136,  -189,  -129,  -163,  -127,   -81,   -68,   -25,    -7,   -95,  -116,   -44,   -60,    14,    21,   -25,    -5,    -7,   -39,    55,    15,    -7,    28,     0,   -26,   -62,   -40,     9,   -70,   -13,   -54,   -29,   -33,     1,   -11,    14,    42,   -49,     6,   -24,    66,    69,   -25,   -76,   -62,    -5,   -74,   -64,   -16,    -6,    -1,   -28,    50,    -1,    33,    71,     0,     8,    21,    43,    61,    41,    43,    38,    42,     6,    39,   135,     2,    14,    36,  -139,   -83,   -51,   -51,    17,     4,     0,   -32,    12,    68,    53,    48,    78,    76,   -20,    34,    -6,   -34,    11,     1,    35,    88,    53,   -12,   -26,   -65,    15,   -50,  -159,  -164,  -104,   -17,   -38,    19,   -13,   -39,   -46,    15,     5,   -15,  -100,    -2,    -7,   -12,   -66,    -6,    19,    15,    74,    32,     1,    -7,   -25,    14,   -31,   -93,  -124,  -147,   -92,   -64,   -52,   -12,   -12,   -48,   -44,   -69,   -35,    56,   -72,   -29,   -13,   -31,    46,     3,   -40,    29,   -26,   -63,   -60,    -6,    -7,    49,   -18,    18,   -26,    27,    40,    76,  -104,     6,     5,   -18,   -48,     2,   -49,   -55,   -28,    -1,   -91,   -56,    55,    27,   -36,   -21,   -22,  -159,  -107,   -19,     9,   -55,   -70,   -90,   -74,   -25,    55,   106,   -97,   -12,     9,    15,   -26,    43,   -66,   -12,  -118,  -127,   -28,   -57,     6,   -59,   -46,   -21,   -80,  -214,   -90,    -8,   -27,  -171,  -213,  -105,  -121,   -54,    69,   -52,   -32,    15,    24,    21,   -15,   -57,   -22,   -42,   -83,   -66,   -37,    -3,    47,   -56,   -51,   -41,   -92,  -124,   -61,  -171,  -162,   -63,   -87,  -101,   -50,  -118,  -135,   -30,   -16,    -8,     4,   -11,    -2,   -44,    43,     2,    15,   -35,     9,    10,    -6,    66,    28,   -45,   -24,   -64,   -28,   -96,   -70,  -136,   -91,   -42,   -28,   -63,   -67,   -22,     7,     8,    -8,   -28,   -26,    76,    -3,   -30,    25,    43,    -7,    -4,     9,    -5,    39,   -99,    -6,    45,    -6,   -45,  -123,  -157,  -100,   -24,    -4,   -99,   -31,   -47,     8,    10,   -12,   -29,  -133,   -11,   -90,    14,   -11,    -1,   -51,   -29,   -17,     4,    64,   -41,   -40,  -110,  -120,   -75,   -70,  -143,   -67,   -71,    -3,   -10,    -6,   -54,    -9,     1,    -5,   -31,   -87,   -38,   -67,    -6,    65,    38,    14,   -87,    10,    37,    53,   -16,    71,  -117,  -124,   -26,   -24,  -122,  -127,   -95,    20,   -18,   -67,   -32,    15,    13,   -18,    21,    34,    40,    19,   -93,    25,    50,  -105,   -15,    47,    61,   -44,   -27,   -85,  -144,   -74,   -42,   -52,   -82,   -59,   -31,    -4,     5,   -23,    -6,     5,    -3,    12,     5,   -69,   -23,   -57,    -9,    86,    87,    57,     4,     7,    68,    65,    79,     1,    -5,     7,    11,    18,    10,    -1,     5,    -3,     6,   -15,    17,   -13,     3,     1,   -12,    17,    25,     4,     7,   -11,    30,    -9,   -38,    -7,    22,    26,    20,     1,    -3,    -2,    25,    19,    -9,     1,    12,    29,    16,    13,    -1,    -7),
		    78 => (  -18,   -14,     3,    16,    10,    18,    -7,    -4,     4,    -1,   -10,    18,     6,   -11,    16,     6,    -8,    13,     6,     6,   -14,     0,    16,   -14,   -18,     9,    12,    17,    10,    17,   -14,   -12,   -18,   -17,     0,    -1,    19,    10,    -4,   -15,    11,     6,   -11,   -55,   -98,   -71,    -6,     5,    -4,    -1,     5,    16,   -10,   -19,   -13,    -1,    14,   -16,    -2,    12,    18,     2,    -7,     7,   -29,   -51,  -114,   -83,   -28,   -15,   -22,    -2,     4,   -29,   -40,   -21,   -24,   -50,   -75,   -34,   -37,   -29,    -6,     9,     0,     1,   -32,    -6,    -8,   -66,   -42,  -100,    57,    31,   -21,   -34,    -6,   -35,   -64,   -36,   -19,   -51,   -10,   -25,   -32,   -28,     6,    20,    -2,   -26,   -53,    14,    -2,     9,     6,    -3,   -60,   -99,    -9,     2,   -26,   -96,   -92,  -116,   -34,   -35,    -9,   -82,   -33,    70,    73,   -39,   -29,   -45,   -65,   -52,   -10,   -37,    20,   -27,    16,   -18,   -11,   -10,   -58,   -78,    21,    17,   -56,  -106,   -81,   -60,   -70,   -19,   -29,    -3,     6,    14,    47,    26,     8,     1,   -33,   -17,   -10,   -21,   -16,   -56,     3,    17,   -49,   -94,   -18,   -78,     1,    16,    -7,    -9,   -60,   -53,    12,    16,    -6,    37,   -17,   -11,     8,     3,    12,     0,    13,    -7,    -3,    -6,   -13,     9,     4,   -83,   -37,    -6,   -51,   -35,    26,    -3,    15,    19,    40,    -3,     8,   -55,    -9,    70,    17,   -16,    58,   -51,   -12,    -8,   -21,   -39,   -29,   -33,   -20,   -19,   -34,   -42,   -38,     2,   -47,   -32,    41,     2,   -11,    -5,    18,    -8,   -29,   -33,    -6,    68,    36,   -77,    16,   -20,   -74,   -29,   -20,     8,   -11,    28,    -7,     7,    -1,   -29,   -78,     2,   -19,  -100,    20,   -23,    22,    -9,    -8,   -69,   -48,   -26,   -14,    58,    24,   -75,    25,     3,   -17,    -3,    -5,   -31,   -61,   -12,   -44,   -98,     5,   -24,   -72,    19,   -20,   -90,   -84,    10,   -11,   -61,    14,     4,   -20,   -65,   -84,    28,   -50,    23,     7,     1,   -16,   -45,   -47,   -78,   -60,   -21,    57,   -70,     4,    10,   -37,    -4,   -45,   -87,   -79,    25,   -24,   -75,   -26,   -47,   -73,   -97,   -31,    47,    -5,     1,    44,    22,   -26,   -92,   -56,    37,    -3,    -2,    80,   -80,   -16,    11,   -50,   -44,   -65,   -46,   -57,    -3,    -3,   -51,   -51,   -47,   -37,   -84,   -83,    50,    40,    19,    40,    19,    -5,    15,    29,   -51,   -30,   -42,   -31,  -118,   -12,     0,   -70,   -45,   -77,   -72,   -57,   -16,   -31,     4,  -103,   -70,  -105,  -115,   -50,    -5,   -25,    10,    63,    22,     8,    27,   -29,   -41,   -52,   -65,   -65,     3,     5,    -6,     7,   -43,   -10,   -42,   -94,   -38,   -23,     2,    -5,   -32,   -14,  -143,   -38,   -49,   -97,   -58,   -34,     6,    -4,   -22,   -65,   -64,   -57,   -19,  -184,   -23,     0,    16,    -1,   -30,     2,    -5,   -50,   -53,   -42,    15,    -4,   -57,   -12,  -104,    -6,     6,   -38,    -7,   -28,   -37,   -30,   -22,   -38,   -51,   -24,   -12,  -163,   -61,    -3,    -9,   -12,   -24,    10,   -28,   -33,    -5,   -21,   -51,   -28,   -32,   -60,   -26,    31,    -1,   -33,     8,   -31,   -39,   -41,   -21,   -50,   -36,   -22,     2,   -89,   -62,    13,    -1,   -11,   -22,    -6,   -29,   -41,   -21,   -38,   -91,   -87,   -65,  -101,    14,    51,    32,   -27,   -62,   -16,   -10,    -6,   -25,   -42,   -21,    -2,   -15,     1,   -63,     3,     8,     0,   -43,    -2,   -32,   -25,     1,   -48,   -70,   -20,   -77,    -6,    37,    17,    -9,    18,   -65,     4,   -18,   -32,   -62,   -11,   -26,    15,    -9,     3,   -35,     4,   -16,   -57,   -58,    11,   -25,   -18,   -57,   -89,     0,   -24,   -37,    31,    30,     0,    51,    59,   -25,   -12,   -30,   -50,   -26,   -26,    -9,    -8,     0,   -93,   -78,     1,     9,   -20,   -11,     7,   -59,   -42,   -34,   -44,    30,    -8,   -33,   -15,   -29,   -67,     3,   -16,    38,     8,   -22,   -87,   -55,   -51,   -24,     5,   -19,   -73,    19,   -71,   -30,   -25,    -3,   -40,   -74,   -54,   -97,    -4,    61,    -4,   -75,    14,   -33,   -66,   -87,     1,    76,    14,    16,   -45,   -14,   -37,   -30,   -30,     4,   -85,    -2,   -36,   -35,   -10,   -31,   -10,   -64,   -27,   -41,   -24,    42,    34,    17,    13,   -31,   -63,   -67,    50,    46,     4,   -11,   -26,   -76,   -63,   -33,   -31,   -16,   -57,    11,     4,     8,   -28,    -6,   -29,   -55,   -48,   -35,   -54,    -2,    40,    36,   106,    32,    12,    -1,    97,     1,   -24,   -96,   -43,   -32,   -45,   -19,   -25,    -5,  -100,    10,     6,   -13,   -14,   -27,    -3,   -25,   -62,   -43,   -55,   -31,   -44,   -47,    11,    -4,    17,    19,    46,   -97,   -93,   -80,   -72,   -29,    -8,   -20,   -68,   -17,   -16,     6,    -5,    17,   -52,   -43,   -14,     3,   -30,   -62,   -58,   -56,   -55,  -139,   -17,    23,    10,    57,   -95,  -133,   -92,   -60,   -11,   -26,     2,     8,    -3,   -36,   -33,     8,    -3,     9,    18,   -16,    13,   -46,   -44,   -33,    -2,   -51,   -77,   -93,   -80,  -107,  -145,   -71,   -32,    -4,   -11,   -28,  -111,   -63,   -57,   -15,     3,    18,    -3,     8,    13,   -15,    -6,    -8,   -17,    -5,   -31,     4,   -24,   -12,   -26,     3,    12,   -45,    -5,   -11,   -53,   -67,    -1,     8,   -21,   -12,   -11,   -19,     3,   -10,    14,    14),
		    79 => (    3,     1,    15,    -1,    -7,    19,   -18,     4,     6,   -16,   -10,     4,    19,    10,    11,    10,    11,   -18,    -2,     0,     5,     1,     8,    -5,     0,    18,     8,    -9,    11,    12,    -2,     0,    14,    11,    20,    14,    20,    15,     2,   -29,   -36,   -29,    10,     8,     9,    -7,    -9,     6,   -20,     0,    11,    13,   -14,     2,    15,   -14,    -3,   -10,     9,   -12,    17,     0,   -14,    -4,    -6,   -27,   -19,   -23,    -8,   -18,   -40,   -17,   -17,   -15,   -14,   -13,    -2,    10,    12,    13,     0,    -1,    -2,     8,     3,    -4,   -13,     6,    15,   -13,   -14,   -20,   -36,   -21,   -50,   -87,   -19,   -53,   -72,   -59,   -70,    -9,    35,    61,   -39,   -23,   -43,   -21,    -6,    -1,    17,     4,     1,    14,    10,     4,     3,   -17,   -78,   -21,   -23,   -61,   -67,    69,    47,    52,     3,   -57,   -65,  -102,  -129,  -115,  -137,   -63,   -50,    14,     5,   -72,   -42,   -16,   -15,     9,     3,   -18,     1,     3,   -14,   -33,  -128,  -160,  -103,   105,    -3,    13,   -29,    45,   140,   -46,   -19,   -24,    49,   -71,   -76,   -34,   -50,   -68,   -76,   -10,     0,   -58,   -23,    -2,   -20,   -86,   -10,  -131,   -50,   -70,   -41,   -57,    41,    42,    74,    41,    21,    36,   -42,   -97,  -115,   -23,   -54,   -35,   -18,   -35,   -45,   -32,    20,   -16,   -32,    11,   -15,  -129,  -123,  -241,    89,  -148,    32,    91,    48,    39,    36,   -47,   -41,  -121,  -227,  -107,   -61,   -55,   -50,   -50,   -28,   -29,   -42,   -40,   -34,  -103,   -38,   -24,   -38,   -78,  -159,  -178,   111,   -34,    79,    95,    83,   -54,  -142,   -27,  -101,   -30,   -78,    46,   -26,   -65,   -35,   -67,   -73,   -50,  -125,    -1,     0,   -69,   -37,   -19,   -98,   -92,  -227,   -38,    97,     2,    54,     8,  -116,  -107,   -80,     7,   -23,    42,   -85,    35,   -14,   -80,    18,   -50,   -35,   -88,   -55,   -25,     7,   -23,     7,    13,   -50,   -41,   -95,    60,   106,    70,   -47,    23,   -78,    42,   150,    94,     0,    71,   104,    59,   -71,  -160,   -68,  -101,   -43,   -67,    -7,   -63,   -19,   -41,     3,   -16,   -43,   -56,   -27,    -2,    66,    18,    10,     7,    82,   103,   137,    49,    88,   113,    29,     4,   -65,   -76,  -102,   -88,   -19,   -77,     3,   -56,    20,    -8,   -30,     4,   -22,   -55,   -96,   -50,   -26,   -32,   -25,    24,     1,    73,     1,     9,    31,    38,     3,    20,   -39,   -51,    -5,  -149,  -143,   -57,   -78,   -23,    10,   -25,   -25,   -85,   -52,   -50,   -94,   -21,   -38,    22,   -87,   -29,   -15,    51,    -5,    99,    78,     1,  -158,   -61,   -78,  -105,   -27,   -58,   -73,   -48,   -75,     2,    -7,   -20,   -50,   -65,   -47,   -48,   -98,   -39,  -128,   -17,   -84,   -53,   -12,    50,   -54,   -27,    29,    20,   -65,  -110,   -73,   -20,    58,   -24,    -5,   -67,   -28,   -18,    12,    15,   -19,   -53,   -11,   -36,   -28,  -200,  -170,     5,    43,    74,    68,   -18,   -15,   -79,    38,    37,  -136,  -110,  -137,    19,    49,   -35,    17,   -40,   -33,   -44,   -10,   -13,   -37,   -26,    -4,   -41,   -42,  -101,  -235,  -204,  -118,    -2,   -26,  -126,   -84,   -75,    -9,   -72,   -63,  -179,  -114,   -29,    33,    -5,    23,   -51,     8,   -21,    -2,    -9,   -54,     5,     6,    43,    34,   -50,   -79,  -153,  -194,  -298,  -157,   -95,   -38,   -59,   -40,   -56,   -76,  -160,   -93,   -31,   -80,   -78,    45,   -19,   -30,   -22,    67,    14,   -46,   -29,   -33,   -68,   -50,   -58,   -79,   -91,  -131,  -250,  -104,   -55,   -39,   -92,   -40,   -21,   -87,  -138,  -190,   -80,   -88,  -124,   -61,    -8,   -19,   -38,    17,   -34,   -12,    -1,   -20,  -106,  -128,    77,   -72,   -98,  -116,  -161,   -48,   -47,   -26,   -49,   -62,  -105,   -48,     2,  -145,    24,    -8,   -24,   -39,   -31,   -41,    20,    -1,   -36,   -24,   -20,   -25,    24,   -87,    28,    33,   -41,     6,   -55,   -30,   -35,   -60,   -91,   -60,   -79,    -7,   -41,  -125,     2,    45,    -9,    80,    22,   -12,     4,    -2,    14,   -51,   -30,    42,    62,  -118,     3,    66,   129,    35,   -12,   -26,   -27,  -109,   -83,  -102,   -16,    -8,     4,   -35,   -61,   -16,    76,    51,    54,   -64,     2,    11,   -17,  -113,   -64,    -1,   -35,  -127,   -83,    64,    84,     4,    66,     8,    -4,   -16,   -56,    -9,   -22,    41,    16,   -12,   -51,   -41,    35,   105,   -85,   -17,   -16,    15,    19,    -7,   -49,   -10,   -70,   -72,  -100,     3,    66,    57,    93,    41,    41,    53,    38,    -8,   -21,    42,   -12,    28,   -89,    33,    24,    78,   -27,   -13,    11,   -10,     2,    -7,  -104,     1,     3,   -25,    -1,    35,    -8,    40,   -14,   -76,   -48,    -3,   -28,    24,    -3,   -80,  -103,    54,    -3,     5,    20,    -8,   -16,   -19,   -12,     1,    -7,    32,   -41,     4,    -2,    54,    91,    -4,    26,   -58,   -70,   -72,   -78,   -30,     4,    16,    79,   -88,  -114,    61,    15,    53,    52,    -4,   -11,     8,    -5,     4,    20,    -7,    46,    19,    -9,   -32,    14,  -154,   -10,    82,    33,   -13,   -11,   119,   -39,  -123,   -97,   -56,   -72,   -15,     8,   -25,    29,    33,   -10,   -17,   -11,    -2,    18,    17,   -16,   -32,   -25,    12,    19,   -34,   -44,   -18,    55,     8,   -34,     2,    57,   105,   -65,     8,     1,     9,   -25,   -14,     5,   -16,    15,    11,   -10),
		    80 => (    2,    19,   -19,    20,    -9,     7,     5,   -15,   -14,   -15,    -3,     9,   -14,    17,    10,    19,   -18,   -18,    19,    15,     1,    19,    -9,     0,    -6,   -15,   -19,     9,   -10,    17,    13,    -8,    20,    18,    -6,    20,    -7,   -15,   -17,    13,    11,    22,   -31,   -13,    11,     7,   -24,    -6,     2,     4,     0,     1,    -3,   -12,   -14,    -1,   -15,     3,   -20,   121,   111,     0,    14,    25,   -19,   -31,   -11,   -87,   -74,  -124,  -134,  -122,   -76,   -90,   -71,   -88,   -67,   -71,   -83,   -52,   -69,   -33,    -6,   -12,   -12,    -4,    17,   146,    88,    45,   -23,   -35,   -61,   -53,   -57,   -32,   -44,    55,    16,   -40,    13,   -24,   -32,    -8,    20,  -135,   -97,   -83,    -2,   -23,   -66,   -15,    -2,     7,   -13,    -6,   -33,   -43,   -60,   -66,   -61,   -37,   -41,   -53,   -92,   -42,   -25,    20,   -53,    12,    70,    26,    72,    43,   136,   -41,    -5,   -49,   -81,   -11,     2,    10,   -27,    24,    14,     8,    26,  -114,  -139,  -117,  -126,  -181,  -102,     0,   -19,   -21,   -39,    40,    43,    35,    93,    57,   146,   -25,    -9,   -55,   -73,   -34,   -18,    11,   -28,   -21,    21,    95,    14,    14,  -100,  -181,  -153,  -162,   -26,    78,    -1,    23,  -109,   -42,     3,    12,   -18,   109,    76,   -76,  -133,  -162,   -90,     0,   -14,    -8,   -14,   -34,    55,   110,    21,   -37,   -62,   -42,   -59,    21,     3,    10,   -69,   -16,   -34,   -27,    -6,    59,    32,   -65,    51,    39,   -26,   -34,  -117,    35,    46,   -38,    46,   -38,    11,    69,    48,   -49,   -56,   -84,  -130,  -118,   -47,   -43,    72,   -57,    31,   -19,    35,    23,    17,    69,    66,    43,   -84,  -111,  -120,   -23,    -6,   -12,    56,   -13,   -50,    64,   -42,   -67,   -32,  -160,   -52,  -103,   -37,   -21,    70,    39,   -73,   -15,    28,    -2,    37,   -19,    31,    82,    70,    22,   -85,    10,     7,    -4,    30,    -6,   -80,   -31,  -131,   -51,   -63,    21,   -58,   -22,    63,    -9,    15,    46,     5,   -70,  -121,   -46,   100,    67,    87,    77,    72,    29,  -148,   -17,   -15,    56,   -45,   -40,   -94,   -95,   -70,    62,    18,   -19,   -39,    13,    13,   -51,   -24,   -67,  -150,  -184,  -175,    -2,    31,    37,     2,    -7,   -23,    -5,   -81,   -11,    18,    50,   -18,   -25,   -41,   -69,   -67,   -11,   -15,   -22,    53,    62,    58,    67,    34,   -35,  -263,  -240,   -58,    47,   -79,   -21,    35,   130,   -13,   -30,   -69,     0,    18,    42,    34,   -66,   -51,   -43,     2,    21,    24,    45,    11,    58,    37,    46,     7,   -72,  -317,  -119,    62,    -8,   -69,   -86,     9,   251,    73,    55,   -64,   -16,     4,    -7,    -2,  -167,   -43,   -23,    31,    83,     1,    28,   -72,    -3,   -20,   -34,  -265,  -222,  -240,  -101,   -55,   -48,   -45,    24,    18,   110,    35,   -29,  -117,    -4,     3,    10,   -37,  -181,    26,   -60,     8,    94,    28,    34,  -106,   -41,    59,    -8,  -188,  -125,   -39,    -4,   -63,   -41,  -131,    17,    24,    70,   116,   -77,  -132,   -34,    20,    14,    -2,  -130,    34,    -4,    -4,    84,    57,   -49,   -50,     9,   -76,  -126,   -50,   -16,     6,   -34,    25,   -70,   -31,   -71,   -29,     7,    68,  -103,   -57,    10,    -2,   -21,   -57,   -63,    23,    78,    34,    88,   -42,    27,    -3,   -57,  -172,  -121,   -74,   -20,   -57,    -2,   -10,    33,    33,   -89,   -61,    21,    60,  -114,   -60,     9,   -19,     9,   -41,    -9,    37,    11,    27,    78,   108,    50,   -92,  -172,  -135,   -57,     5,    13,   -19,    -3,    32,   -64,   -11,   -26,    33,    17,    12,   -53,   -34,   -25,    20,    24,  -108,   -34,   125,    -6,     9,    57,    27,    53,   -83,  -158,   -67,   -86,    -3,    24,   -65,    17,   -50,   -33,   -97,   -26,    34,    -2,    46,   -74,   -13,    16,     5,    29,  -150,    37,   107,    23,    53,   -14,    40,    34,   -17,    29,   -32,   -41,   -21,  -108,   -24,   -28,   -28,  -105,  -117,   -40,    13,   -15,    14,   -64,    20,    20,     9,    19,  -147,    40,    21,    17,    60,    88,    21,    42,     4,    -3,   -54,   -36,     6,    45,     2,   -15,   -79,  -100,  -141,  -147,   -88,   -24,    75,   -40,    18,    27,     8,   -15,  -167,    -1,    -3,    75,    93,    38,    34,    28,    37,   -48,   -58,    13,    61,     4,  -141,  -111,   -49,   -59,  -167,   -99,   -18,   -13,    64,     8,     2,    22,    16,     0,   -26,  -119,  -133,    19,    13,     3,    18,    56,    67,    59,     6,    46,    47,   -86,  -133,   -84,  -123,  -111,  -159,   -74,    28,     4,   -93,     0,   -10,   -14,     1,    -8,   -36,   -27,   116,   149,    -8,   -34,    12,    79,   133,    86,   119,  -126,  -110,  -114,  -230,  -195,  -111,  -119,   -57,    15,   -16,    -5,    49,    12,    -7,   -17,    12,   -19,     2,    -1,   -79,  -151,  -139,  -142,  -120,   -77,  -100,  -123,  -163,  -120,   -48,  -133,  -140,  -129,  -155,  -112,    -8,   -30,   -25,   -23,    -5,    -2,   -16,     8,    18,    11,   -12,   -18,   -16,  -112,  -153,   -37,    -3,   -39,   -64,   -75,   -40,   -56,   -45,   -81,   -87,  -144,  -153,   -33,   -94,   -39,   -39,   -22,     0,    10,   -17,    11,   -17,   -20,    19,    15,     3,    10,    14,   -17,    -6,    -3,     5,    13,    14,    -8,     3,    -3,    -8,     8,    -2,   -26,   -16,   -26,   -26,   -20,     2,     1,    17,   -15),
		    81 => (  -17,     8,    17,    18,   -12,   -12,     3,   -16,   -18,    10,    -8,    18,     3,    -6,    18,    -5,     7,    -3,    11,    -2,    13,    -5,    15,    -3,   -19,    14,   -14,    15,    -9,     5,    12,     1,     2,   -17,     2,    -4,     4,    19,    -1,   -12,    -3,   -31,    21,    26,   -11,   -28,     2,   -15,    -6,    -2,   -11,    10,    11,    -5,    10,   -11,   -12,    10,   -14,    18,    -4,    14,    -2,   -20,   -23,   -22,   -23,   -17,     0,     4,   101,   124,   264,   196,    98,   -65,    16,   -87,   -65,   -50,    -7,    14,    15,   -10,    -5,     0,    45,    36,   -20,   -67,  -138,   -46,    89,    28,   -56,  -101,   -85,   -21,    41,   146,   164,    32,     5,   -70,     4,    91,   -20,    -4,   -68,    -3,     9,    -8,    12,    19,    50,    44,    94,    41,   -29,   -37,   138,   106,    64,   -12,   -10,   -59,   -14,    37,    47,    25,   -32,   -33,    70,    92,    42,    67,   -12,   -50,   -47,   -64,    -4,   -18,   -11,   -14,   108,   209,    90,    78,    55,    21,    15,  -105,  -106,    20,    67,    17,   -34,    19,     6,    37,    69,    71,    62,    21,    11,   -24,   -58,   -58,    14,     8,  -134,     9,    17,    44,    90,    29,   -61,   -77,    41,   -22,    -2,   -17,   -11,   -22,   -78,    57,    29,    98,    56,   -16,    25,    -9,    -8,   -12,   -30,   -14,   -20,    14,  -150,  -132,  -130,    -7,    51,    61,  -101,    20,    70,   -59,   -12,   -85,   -18,    56,   -17,    21,    54,   107,    17,   -10,    36,   -31,   -34,     2,   -62,   -34,    -6,   -13,  -169,  -102,  -124,   -22,    24,     4,   -27,    47,    26,    20,    44,   -81,   -87,    18,    61,     7,    63,   -87,   -52,   -42,    21,   -53,    -6,    -5,   -65,   -12,     9,    -8,  -164,   -67,   -81,   -88,     3,    45,    71,    10,    16,   123,    97,   -60,  -110,   -32,   -58,   -60,   -62,   -44,   -37,   -45,   -61,     0,   -23,    13,    11,   -21,     3,    -7,  -129,   -21,  -145,   -72,  -130,    13,    55,    84,    36,   135,    35,   -35,   -56,   -35,   -84,   -67,   -25,  -120,   -76,   -87,    -6,   -11,   -24,   -17,    23,     3,    -3,    26,   -29,   -12,  -119,   -65,  -113,     3,   -55,    37,     9,    72,    29,   -27,   -15,   -83,     9,   -88,   -80,  -106,   -67,   -52,    13,     1,   -17,   -15,   -12,    20,    -9,    -8,   -17,   -44,   -84,   -85,    38,    74,    16,     6,   -38,    11,    -7,   -67,   -86,   -23,   -27,   -93,   -35,  -109,  -159,   -71,   -38,   -37,   -20,   -25,    11,    35,     0,    -5,   -23,   -18,  -112,    45,    74,    76,   104,   -42,   -59,    -4,   -22,   -89,   -38,    54,   -28,   -65,   -73,  -230,  -106,   -90,   -75,   -65,   -58,    -6,    -7,    -5,    -9,     1,    13,    -4,   -96,    84,    71,   -17,   -31,  -132,  -173,   -98,   -61,   -53,    26,    36,    -5,   -57,   -94,  -152,  -136,  -158,  -103,   -68,   -39,   -62,     5,    12,   -17,    11,    -7,    30,   -19,   -78,   -47,   -47,   -89,  -116,  -146,  -152,  -175,   -14,    76,    15,   -22,   -65,   -90,  -202,  -115,  -121,   -95,  -100,  -231,   -33,   -11,   -27,    11,    -6,    26,   -49,   -43,   -45,   -70,   -68,  -153,   -84,   -92,  -161,  -140,   -13,   100,    74,   -24,   -88,   -73,  -157,  -135,  -165,   -59,  -113,   -78,   -30,   -20,   -32,   -10,    -9,    -9,   -84,   -22,   -38,   -66,  -118,  -119,  -113,  -129,  -277,  -153,  -125,    46,   -44,   -39,   -49,     7,   -60,   -81,   -60,     0,   -67,  -122,  -129,   -10,   -46,   -24,    10,    12,   -22,   -23,   -99,  -195,  -113,  -193,  -128,  -139,  -353,  -307,  -171,     0,   -60,   -27,    25,   -31,   -26,    68,    45,   102,   -46,  -231,   -52,   -52,   -42,    -7,     0,   -23,   -43,   -67,  -179,  -103,   -24,    -9,   -70,   -97,  -167,  -109,   -85,   -59,    42,    83,    11,   -73,    -5,    35,     1,    -9,    44,   -13,    -8,   -78,   -24,    12,   -19,   -50,    66,    -6,  -134,   -56,    22,    27,    58,   116,    16,   -28,    10,    42,    39,   110,    67,   159,   119,    99,    -6,    39,    47,    25,    15,   -59,    13,    43,    20,   -67,    71,    86,    31,    91,    80,    99,    99,    55,    55,    -6,    37,    39,    88,    23,    92,   150,    45,    55,   -12,   -74,   -40,    32,    66,   -75,    16,    44,     9,  -190,  -115,    57,   139,    46,    11,    24,    40,    41,    32,    22,    36,   -13,    30,   -35,    36,    20,    83,    87,    45,  -147,   -94,    21,   -14,    -7,     4,    19,    10,   -19,   -55,    29,   -29,    47,   -22,   -10,   -36,   -53,     9,     8,    59,   -70,  -110,  -150,  -122,   -40,    24,    70,    82,   -34,   -82,   -81,  -101,    50,    11,     1,    -1,   -15,     2,   -34,   -56,   -78,   -16,    24,    46,   -24,   -16,  -140,   -92,  -181,  -150,  -137,   -84,   -54,   -17,    19,    35,   -47,   -62,   -89,   -14,     1,    16,     1,    -8,    18,   -23,    -7,   -11,   -39,   -14,   -11,   -89,   -39,   -57,   -80,   -94,   -61,  -121,   -90,  -103,  -124,  -103,  -124,  -102,   -80,   -35,     1,    10,     4,   -15,   -15,    18,   -12,     5,   -29,   -33,   -39,   -31,   -24,   -86,     4,   -15,   -42,   -67,   -46,   -83,   -22,   -87,   -50,   -71,   -53,   -42,   -29,     7,   -16,   -10,    13,    -8,     9,   -11,    -7,   -16,    -1,    18,     5,    -6,    -4,   -11,   -31,   -30,    -3,   -24,   -20,   -24,   -25,   -19,   -16,    -3,     1,     1,    -8,    -2,     9,    12,    -7,    20),
		    82 => (    4,     5,   -15,   -12,     0,    -9,     7,   -19,    19,     0,    -2,     4,   -18,    -2,    24,    19,    -5,     4,   -13,    10,    -7,   -20,    15,    -6,   -20,     9,    -3,    -4,     1,    17,    18,    -4,   -16,    19,    11,   -47,   -75,   -30,   -69,   -65,   -76,  -136,   -58,     8,    66,     9,   -77,  -148,   -98,   -52,   -74,   -24,    -6,   -12,    -5,     6,    11,    19,    -1,  -105,  -110,    16,    -5,   -18,     0,   124,   106,    48,    28,    34,    15,    49,    -3,   -11,   -57,   -95,   -58,   -45,   -34,    -4,    17,    22,    -1,     3,    -4,   -11,    -6,  -117,  -150,   -19,    -5,    40,   -44,    51,    22,    18,   -35,    39,    86,    46,    46,    10,   -51,   -65,   -43,    17,   -78,  -190,    20,    26,     9,     3,    -2,    12,   -31,    32,    30,   -50,    13,   -20,  -100,    48,   100,    15,    15,    59,    76,    26,    45,    23,   103,    12,    -5,   -35,   -90,   -43,   -61,   -21,   -43,    -2,     1,   -17,    29,    -8,   -11,    26,    29,   -94,    -9,    26,   -64,   -45,    24,     0,     0,   -18,    69,   -29,    18,   -47,   -30,   -28,   -59,   -32,  -129,    -4,   -51,   -42,    -7,     6,    10,   -46,   -50,     8,     5,    75,   -66,   -56,    22,   -38,   -87,    79,    -5,    22,    92,    14,    28,   -77,   -43,    -8,   -48,   -69,  -159,    64,   -31,   -22,   -15,     9,   -16,   -43,   -48,   -21,    45,     0,   -66,   -57,    55,    14,    -3,   -62,     5,    44,    -5,    13,  -107,   -23,    46,    72,   -14,  -158,   -59,    19,   -78,   -36,   -32,    30,   -31,   -67,   -39,   -98,   -58,     4,    40,    32,    78,    44,   -91,   -56,  -111,    -7,    -2,    20,    35,    76,     6,    13,     7,   -74,  -131,  -159,   -59,   -25,    -4,   -31,   -16,   -56,   -35,  -132,  -113,  -142,  -173,   -46,     5,   -90,  -137,    -7,   -16,   -81,   -21,    29,    55,   -58,   -24,    88,    -4,   -72,   -70,   -85,   -55,   -48,   -17,     7,   -17,   -90,   -93,  -127,  -144,  -276,  -392,  -354,  -285,  -230,   -70,   -85,   -16,   -93,     7,   -37,    39,     7,    -7,   -30,    -7,   -36,  -119,   -97,   -45,   -20,    -5,   -54,   -53,  -107,  -105,  -131,  -196,  -237,  -314,  -268,  -225,  -124,   -94,  -130,   -29,   -88,   -61,  -141,  -138,     5,    -3,    10,    45,   -38,  -118,   -14,   -48,   -35,    19,   -63,  -133,   -99,  -167,  -122,  -113,  -147,   -40,   -35,   -22,    26,   -18,   -25,    17,   -59,  -103,  -123,   -91,   -48,   -26,    39,    87,   -98,   -98,   114,    14,   -27,   -19,   -57,     8,   -35,   -80,   -57,    18,   150,    65,   -16,   -39,    30,   144,    98,    39,    22,    -3,     3,   -53,   -68,   -11,    53,   115,    -8,   -21,    50,    -7,    -2,    -1,   -60,   -83,   100,    63,   -14,   101,   152,   126,    87,   125,    96,    80,   129,   114,   -15,    61,  -106,   -57,   -20,    46,    -9,    22,    21,   -23,    70,    61,    55,     2,   -37,    20,   232,   100,   124,    75,    70,    60,    63,   108,    37,    60,    33,   -54,    39,   -19,    18,   -45,    -3,   -57,   -36,   -23,    65,   -14,    95,   179,   110,    -4,     5,    20,    94,   -35,   122,   186,    86,    38,    58,    71,    11,   -67,    41,    42,    34,    27,    33,   -10,     5,   -58,   -69,   -39,   -28,   -79,   134,   177,    71,    14,   -28,    11,   -52,    52,    36,   122,   -33,    57,   -45,   -63,    29,     1,   -22,    89,    59,    60,     9,    -4,   -59,   -12,  -137,   -95,  -113,  -145,    20,    40,   117,    11,   -15,   -72,    23,    -7,    90,    95,     1,    -1,   -41,   -62,   -33,    -4,    25,   -21,    -5,    64,    17,    57,    83,    44,   -38,   -63,   -56,    22,    91,    51,   112,     7,   -67,   -67,   -28,    56,    53,    67,    57,    32,    17,   -54,    14,     5,   -22,   -58,   -13,    18,    -3,    69,    81,    12,    66,    70,    30,   107,   100,    81,    58,   -12,   -78,     6,   -10,    40,   125,    42,     7,   -19,   -71,   -43,   -81,  -107,   -92,   -94,   -18,    -3,   -76,   -52,   -13,   -25,    -1,   -30,    24,   122,   -18,    35,    -5,   -20,    51,    -1,    31,    53,    38,    33,    31,    51,   -64,   -76,   -19,   -24,   -95,   -68,   -62,   -71,   -24,   -64,    -5,    47,    80,    34,    68,    37,   -66,   -43,    -9,   -18,   -12,    -9,    25,    59,   -60,   -54,   -25,   -19,   -59,   -19,    16,   -35,   -86,  -115,   -42,   -73,   -84,  -110,   -19,     8,    18,   -27,   -38,   -46,  -116,  -126,   -15,   -15,   -19,    30,   102,    93,    16,  -102,   -22,   -66,  -120,   -35,   -73,   -10,  -148,   -80,  -135,   -51,   -69,   -90,  -154,   -74,    -4,    61,   -95,   -89,   -67,   -84,    13,     7,    15,   -53,   -38,   -38,   -16,   -36,   -79,   -93,  -159,  -185,  -137,  -110,  -178,  -136,  -115,  -112,   -48,   -71,  -154,  -188,  -109,  -172,  -105,    29,    51,    52,     5,     2,     5,   -27,     3,   -39,   -33,   -25,   -54,  -108,  -142,   -50,   -32,   -47,  -127,  -101,   -64,   -97,  -120,   -76,  -159,  -121,   -73,   -93,   -33,   -37,    33,    68,     0,     7,    13,    -8,     8,   -35,   -54,   -48,   -35,   -43,   -18,   -14,   -11,     0,    -4,   -53,   -26,  -129,   -98,   -80,   -54,   -31,   -26,   -17,   -39,    18,     1,    -8,     1,    17,    20,    -2,    -5,   -12,     1,     3,   -17,     6,    16,   -37,   -16,   -17,   -36,    -7,   -12,   -10,     0,   -26,   -27,   -47,   -59,   -37,   -14,    -2,    -4,   -12,   -14),
		    83 => (   18,     4,    10,    12,    -8,    -8,   -17,   -18,   -13,    -2,    -7,   -15,    -5,    -3,   -30,   -27,    -7,    -7,    11,     2,    15,    -1,    12,    19,     7,   -17,    12,    17,     0,    10,     4,   -11,    12,   -16,     5,   -16,   -20,    -4,   -34,   -23,   -29,   -87,   -67,   -65,   -34,   -98,   -48,   -51,   -28,   -21,   -21,    -5,    20,    10,   -16,   -18,    -6,     7,    -4,    -3,   -43,   -39,   -48,   -51,   -98,  -126,    48,    -6,   -43,   -77,  -104,  -101,   -71,   -11,    13,   -89,  -120,  -158,  -143,  -119,   -21,    19,   -15,     6,   -12,    14,   -22,   -25,   -21,    45,    84,   227,   216,    83,    94,    91,    69,    29,   -16,   109,   142,    93,    82,   187,   330,    33,  -206,  -214,  -108,   -59,     5,     6,    17,    -9,  -130,     7,    44,    67,    26,   138,   176,    -1,    98,    46,    53,   -16,    39,     3,    62,    99,    79,    83,    35,  -111,  -113,  -422,  -325,  -121,   -86,     9,     6,    17,   -19,   -11,   -14,    70,   157,   196,    20,    47,    75,   -34,   -65,    10,   -38,   -11,    91,   -50,   -19,    56,    16,   -24,   -31,    28,    33,  -158,   -72,     9,    10,    24,    44,    -7,   -21,   137,   212,   176,    85,    88,    40,     6,   -55,    29,    -8,    59,    49,    19,    22,   -13,     9,   -26,    -5,    20,    68,  -185,   -87,   -31,    -6,    11,     4,    38,   -18,    29,   197,   254,   132,     8,    18,   119,    18,   -68,    20,    -5,    49,   -35,   -64,    36,   -32,   -36,   -54,   -24,    57,  -167,  -105,   -47,   -58,   -21,   -78,    -6,    34,   141,    25,    67,    17,   -30,   -24,   -92,  -111,   -66,   -28,   106,    52,    65,   -81,    55,    16,   -72,    49,     7,   -51,  -109,  -101,    -7,    -1,   -43,  -194,   -43,   205,   197,    85,    88,   101,   -47,    40,   -63,   -53,   -32,   -51,   -48,    11,   111,    54,   -19,    37,   -44,   117,    93,  -227,   -97,   -71,    12,   -19,    -7,  -213,    13,    44,   101,   122,   155,    -1,   -43,  -101,  -119,   -64,  -103,   -31,   -54,    -9,    68,    81,    31,   -88,   -69,    39,   147,  -102,  -107,   -84,     2,   -18,   -76,   -98,   111,   174,   164,   101,    40,    75,   -41,   -17,   -92,   -95,   -29,    -7,   -87,    14,    20,    45,   -79,  -106,   -53,     7,   -43,  -272,  -190,   -91,   -20,   -19,   -24,  -101,    43,   113,   164,   115,    61,    18,   -69,    31,   -41,   -56,   -60,   -68,    15,    20,    -7,    18,    37,   -57,  -122,   -51,     9,  -171,  -118,   -41,   -12,    18,   -27,   -86,     7,   175,   123,    77,    59,   135,   -11,    52,   -42,   -58,   -21,   -37,    73,  -187,   -52,    85,    72,   -63,   -68,   -87,    53,   -30,  -189,   -46,   -16,    -5,    47,   -19,    41,    77,   130,   129,   -15,    55,     4,   -40,   -24,    -2,   -50,    36,   -87,   -89,   -23,    50,    55,    38,    25,   -35,    52,   -30,  -260,  -114,    14,   -23,    53,   -46,    24,    60,   163,    98,   -91,   -49,  -102,   -10,   -70,   -30,   -74,   -59,   -32,   -87,   -97,   -32,   103,    11,    32,    59,   116,   131,  -266,    47,   -53,    15,     5,    23,   171,   159,   136,    21,    53,  -120,     5,    12,   -98,  -158,   -27,    15,   -42,   -96,   -72,    83,   127,    21,   -51,    59,    14,    88,  -299,  -126,   -68,     1,    28,   -35,    83,   106,    27,   -36,    19,   -45,   -30,   -72,   -71,     2,     0,   -96,   -62,    28,    28,    61,   119,   -19,    12,   -61,   -45,   -61,  -241,   -73,   -35,   -41,    26,   -13,    53,   135,    94,     0,    -7,   -38,   -95,    -2,   -31,   -76,    76,    -1,    73,    -7,    49,   122,   -61,    38,   -48,   -31,  -150,   -43,  -237,   -13,   -62,   -13,   -38,    41,    28,    53,    89,   -48,   -66,   -83,  -146,   -73,   -85,   -17,    25,    89,    80,     6,    76,    63,   -33,    37,   -19,   -37,   -57,    36,  -121,   -96,   -72,   -10,    34,   -98,    23,    49,    62,     0,   -27,   -87,    -4,   -71,   -61,   -30,     2,    80,    54,   153,   106,   -21,   -27,    66,    54,    64,    70,   -10,  -168,   -75,    -7,   -21,   -22,    40,   -10,    18,   -86,    64,   112,    -3,   -31,   -57,     0,    35,    74,   115,   124,    85,    38,    54,   112,   -10,    57,    93,   -27,  -133,  -164,   -87,   -16,   -20,     1,    87,    64,   -90,    51,   111,   129,   -25,    22,    65,    32,   -41,    26,    71,    37,   -55,    45,   -28,    86,    13,    76,   171,    36,  -102,  -114,   -69,   -16,    14,    15,    37,     9,   -50,   -26,    49,   113,    41,    33,    22,    58,    -7,   -37,   -33,    55,    41,   -11,   -43,   -74,     6,   173,   165,    80,   145,    59,   -90,    16,     6,     4,    97,   162,   142,    -2,   110,   101,    71,   124,    43,   -39,   -35,    15,    42,   -37,    -7,    14,   -73,    37,   223,   142,    80,    93,  -145,   -86,   -28,    -6,    17,     1,    23,   -47,     3,   135,   107,   -19,    44,    49,   -61,   -27,    46,   139,    11,   -19,   -19,    25,    63,    73,   -62,  -173,  -198,  -193,  -153,   -46,   -32,   -19,    -1,    15,    -1,   -25,  -194,    88,    45,    13,    59,   -45,   -37,   -88,   -88,   -50,   -68,     5,   173,   187,   171,    32,   -38,   -73,  -209,  -100,   -11,   -12,     7,    17,    -2,   -13,    13,     8,   -32,   -59,   -55,   -26,   -44,  -123,  -108,   -89,   -72,  -119,  -105,   -66,    -9,   -26,   -10,   -89,  -112,   -34,   -37,   -24,    16,    11,    12,     8),
		    84 => (    1,    -4,    19,    11,     9,     3,     8,     6,    16,    -1,     3,     0,   -66,   -35,   -23,   -33,     1,     6,     9,   -14,    12,     2,     9,    -4,    -7,    11,    -2,   -12,    10,   -14,     6,    -8,   -12,   -39,   -64,   -87,   -51,   -84,   -77,   -74,   -92,  -102,   -22,   -92,   -84,   -15,   -49,   -47,   -86,   -56,   -37,   -75,     1,     9,    13,   -16,    16,    10,   -43,   -73,   -99,  -122,  -108,  -112,  -181,  -156,  -222,  -240,    22,    48,    -6,  -120,  -110,  -140,  -207,  -115,  -234,  -107,  -112,   -74,   -40,   -52,    19,     9,    15,    -5,   -12,  -215,  -138,  -150,   -85,  -127,   -99,  -195,  -170,  -178,  -108,  -237,   -28,   -16,  -118,   -70,   -65,   -12,    84,    -2,  -108,  -126,   -71,   -45,   -21,     1,     9,    20,   -92,  -206,   -20,    -2,    42,     3,  -101,     7,   -29,  -143,   -14,   -30,   -68,   -90,   -43,   -11,   -25,    12,    -1,   -64,    24,    33,    49,   -37,  -138,   -22,   -20,   -18,  -106,   -15,     5,   -28,    -9,   -24,    52,   -31,    75,     3,    87,   -68,   -40,   -98,   -66,    55,   -18,    12,   -91,   -37,    16,    -9,   -49,    49,   -55,    -6,    -8,    12,   -56,   -86,    42,   106,    68,   -94,   -32,  -106,   -11,    32,    -6,   -67,  -159,  -166,  -127,   -94,  -132,   -74,  -163,    -6,   -11,   -12,   -38,   -17,    -3,   -70,    16,  -190,   -70,     2,    46,    80,   -80,  -101,  -147,   -67,   -33,   -12,  -108,   -86,  -115,  -146,  -125,   -38,   -73,   -91,   -83,   -60,   -66,   -49,    24,    95,    86,  -119,   -64,  -163,   111,    31,    85,    33,  -139,  -151,  -164,   -69,  -140,   -94,   -68,   -17,  -196,  -113,  -112,   -28,   -46,   -23,   -79,   -91,   -60,   -17,    76,    87,     1,   -40,    -3,  -129,    92,    24,   -72,    -5,  -101,   -65,   -83,   -87,  -131,   -36,     2,   -49,  -113,   -44,   -69,   -29,     5,    50,    39,    91,    48,    62,    98,   -71,  -121,   -40,    20,   -81,    65,    16,   -53,    59,   -40,   -98,   -48,    -9,    -5,     4,    74,   -27,   -55,    78,    64,   128,   -31,     6,    54,    38,    32,   -10,   -14,    19,   -64,   -27,   -13,   -96,   -15,     1,     5,   115,     1,     8,    35,   125,    98,    60,   121,   -34,    11,    82,   128,    26,   -52,   -24,    -2,    20,    55,    52,   -21,   -25,  -136,  -121,    -5,    -8,    57,    64,   -20,    87,    69,    51,    77,    96,    93,    87,   111,    45,   -36,   -10,    11,   -21,   -65,   -12,   -22,    50,    90,    49,   138,    79,    67,  -138,    14,   -21,   -11,   114,    51,   101,    41,    75,     5,    53,    59,   147,   130,    75,     2,   -41,    65,    43,   -80,    15,    20,    94,    68,    87,    70,   184,   168,   -82,    13,    26,  -177,    49,   167,   117,    58,    48,   100,    69,    56,    46,    89,    -1,   -29,   -51,    73,   123,   -67,   102,   -47,   118,    58,   -51,    -5,   107,   107,   -20,    -9,    30,   178,    83,    -4,    95,    34,   -43,    23,    47,    59,    46,    29,    20,   -22,    70,   108,    21,    -4,    90,   -12,    -6,   109,    62,   -45,    73,   204,   -28,     1,     9,   -39,   114,    37,    86,   112,    84,    59,    24,   -10,   -30,    37,     3,   -23,   123,    41,    56,   117,   154,    45,    23,    -1,     4,   -13,    63,   129,   -48,   -15,   -31,    51,   -43,   142,   104,    45,    66,     9,    17,     6,    -4,     8,    41,    37,    38,    60,    17,    10,    71,   -57,     1,    26,    28,    27,    18,    82,    -6,  -111,     1,   105,    46,   109,    -2,   -25,   -27,    35,    72,     7,    55,    18,    82,    91,    13,    14,    25,    46,   -39,   -33,     6,   -21,   -59,   -31,  -117,   -37,   -42,     6,   -76,   -57,   147,    -9,   112,    17,   -94,    48,    15,   -56,    14,     6,   -34,    71,     8,   -42,   -51,   -67,  -124,   -88,   -74,  -131,  -144,   -37,   -88,   -44,   -41,    -5,   -20,  -101,    99,    56,    -3,    10,     4,    22,   -81,  -186,  -104,  -136,   -64,   -28,   -82,   -39,  -102,  -123,  -105,  -186,  -140,  -104,  -130,   -44,  -205,   -36,     1,    -6,   -32,  -159,    48,    64,    23,   -89,  -147,   -47,   -86,  -127,   -76,  -108,   -81,  -128,   -58,    -3,   -50,   -81,  -131,   -46,  -108,   -55,   -89,    24,  -122,  -135,    -9,   -22,     2,     0,  -118,  -184,   -31,    -1,  -145,  -158,  -140,   -27,   -42,   -99,  -110,   -62,   -35,   -74,   -89,   -71,   -30,   -98,    22,    15,    60,   -63,   -46,   -23,   -35,   -15,    -6,    -6,  -158,   -74,  -186,     1,    49,    12,  -112,    54,   -55,   -41,   -47,   -59,   -39,   -50,     5,   -59,   -21,   -57,    24,   -39,  -100,  -134,    12,    -7,    17,    -7,     5,     1,   -20,  -146,   -12,    42,    63,    57,    38,   -72,   -24,  -130,    44,    67,   -64,    -4,   -71,  -160,  -103,   -18,    47,   -24,   -77,  -227,   -36,   -56,     9,     4,   -13,   -45,   -26,    29,  -109,    26,     2,   -48,  -104,   -38,   -42,  -136,  -112,   -52,  -167,   -25,   -59,   -80,  -128,   -36,    -8,    54,   -19,  -143,   -68,   -47,    -5,     9,    14,    -2,  -119,   -56,   -31,  -122,  -138,   -59,   -65,  -200,  -143,  -100,  -209,  -187,  -134,  -183,   -72,   -44,  -198,  -271,  -260,  -232,   -65,   -59,   -19,   -15,   -12,    16,     2,    14,   -14,   -10,   -27,   -22,   -27,   -43,   -49,  -157,  -173,   -94,  -129,  -165,   -53,   -87,  -179,  -111,  -126,  -153,  -114,  -105,   -29,    12,   -12,     9,   -17),
		    85 => (    5,    -3,    17,   -20,     0,     1,     5,   -20,    -5,   -15,   -17,   -15,   -12,   -28,    -3,    11,    10,   -13,     8,     0,   -11,   -17,     2,     7,    20,    -4,   -15,   -15,   -11,    18,    -3,   -12,   -20,   -11,   -17,    16,     5,    14,   -32,   -74,   -70,   -83,   -61,   -58,   -85,   -78,   -98,  -122,   -69,   -64,   -30,   -14,   -19,     6,    -7,    -5,     4,    19,   -36,   -36,   -27,   -25,   -55,   -38,  -191,  -149,  -225,  -198,  -156,  -162,  -163,   -27,   -19,    31,    41,   -38,    46,    20,   -19,    44,   -73,   -37,    13,    11,     4,    13,   -60,    66,    94,   -61,  -213,  -169,   -31,    18,    66,  -112,  -134,   -23,   -73,   112,    82,    41,   156,   121,   134,   257,   203,   144,   -61,    64,    48,     2,    -7,    -5,   -71,    71,  -219,  -194,  -107,   -65,  -212,   -58,    68,   -55,   -51,   -99,    28,    98,    94,   158,   294,   137,   148,   177,   307,   142,  -100,    21,   -69,   -54,     7,    16,   -99,    99,  -237,   -78,   -69,   -61,    -2,    70,    88,    12,   -63,  -105,    41,    40,   102,   141,   174,   183,   229,    45,   142,    45,   -57,   -71,  -104,  -115,     6,     7,   -22,  -224,   -35,   115,   114,    49,    99,    47,    45,     0,     2,   -99,   -11,     8,    26,    -6,   127,   204,   126,     2,   110,    94,   152,   150,    24,    30,    -6,   -33,   -17,  -249,  -137,   -55,    54,    23,    11,     0,     2,    89,   -76,   -42,   -48,  -153,   -37,   -52,    91,   157,    53,    72,   239,   197,   180,    45,    80,   142,   -65,   -75,  -106,  -263,   -82,   -95,    39,    64,   -19,    -5,   -86,    38,    59,    -5,   -57,  -114,  -151,   -24,   -49,   148,   107,   109,   203,   175,   114,    19,    61,    89,    13,     1,  -107,  -141,   -68,   -59,   -35,    41,    25,   -59,    22,    12,   -15,    -8,   -90,  -155,  -154,  -116,   -26,   127,    13,    34,   105,   141,   143,    74,    10,    -4,   -10,   -25,   -72,  -225,    43,    -3,   -92,  -101,     3,    55,   -91,    71,    65,   -55,   -91,   -67,  -177,  -143,    44,    20,    25,   110,   100,   157,   186,    34,   -52,   -55,   -11,   -19,     5,  -160,    36,   -77,     5,   -77,    23,   -31,   -44,    -7,    21,   -48,  -119,   -65,    69,    36,    -4,    17,   -86,   -30,    78,   134,   171,   114,   -61,   -44,     5,    -1,   -30,  -119,   141,   -23,   -28,    59,    50,    76,   154,    12,   115,   -32,   -30,   -97,   -23,   -44,   -23,   -91,  -100,   -80,     3,    34,    46,   134,   200,   -66,    16,   -12,   -15,  -141,    14,    22,   -28,    97,     2,    -3,    51,    68,    88,   -29,   -72,   -19,   -32,   -75,  -114,    30,   -34,    76,   -87,  -125,  -130,   -85,   142,   -62,     3,     5,   -45,  -153,    83,    42,   126,   -17,    -1,    76,    75,    68,   -41,    13,    27,   -12,    -5,   -50,    24,    -7,    77,   -23,    61,    -2,   -27,  -153,  -156,   -65,    34,    -7,   -93,   -29,   108,   149,    13,    65,   -28,    33,    62,   -18,   -25,     9,   -29,  -148,   -49,    21,   -27,   -22,   -39,   -23,    12,    46,    37,   -68,  -122,   -36,    -1,   -22,  -109,   -37,    41,   132,   169,    61,    20,    28,   -44,   -53,   -79,     4,   -37,   -80,  -128,     8,    78,    19,   -58,    62,    93,   -10,   -97,  -199,  -176,   -51,     6,   -30,  -137,   -25,    93,   171,    64,   212,   117,     5,   -13,   -37,  -152,   -29,    25,   -78,   -43,   -64,    22,    17,    67,    16,    77,     5,   -63,  -202,  -304,  -186,   -38,   -23,  -139,    -7,    25,    50,   182,   148,   136,    62,   -95,   -33,  -132,  -146,    49,    26,   -30,  -105,   -37,   -33,    81,   -19,   -14,    13,   -89,  -200,  -173,  -153,    15,   -51,    76,   112,    11,   105,   162,    74,     1,    19,    22,    27,   -64,  -106,    26,    67,    32,    28,   -46,    -1,   -79,    44,    -8,    59,    70,   -38,  -202,  -116,    -9,   -36,   130,    95,   119,   221,    93,     6,    43,    96,    16,    47,   -38,    40,     7,   106,    29,    25,    25,    28,   -38,    -2,    -7,    70,   -87,    39,  -248,    11,    -7,   -25,  -110,   -14,    72,   140,   216,    47,   -42,    14,   -34,   -55,    21,     9,   -19,   -54,    -3,    -5,    40,   -11,    18,    42,    37,    14,   -55,    35,    30,     1,     7,   -10,  -199,  -104,   -21,    20,   -24,    90,     3,    29,   -17,    50,   -37,   -40,    78,    42,    47,    84,   -19,    90,    43,   -19,   -67,    17,    20,    65,   150,   -10,    -8,    -9,    60,   -29,    25,     7,    51,    34,   -35,   -29,   110,    53,    65,    98,    67,    63,    47,    30,  -167,   -61,    18,   -38,   -90,   -17,    94,    81,   181,   -19,    -4,   -19,  -108,   -71,  -136,   -16,     1,    -1,    66,    84,    29,    37,    71,   103,    92,    65,    97,    38,    44,     4,   -35,   -29,   -39,  -111,    30,  -183,   -82,   -11,    -7,   -17,   -25,    92,  -199,  -187,    -3,   -38,    10,   -39,   -13,   -15,    -4,    33,   -65,   100,   111,    96,    32,   106,    98,    99,   183,   165,   125,   -48,    -8,   -19,    -5,    20,     8,   -69,  -113,  -139,  -180,  -249,  -121,   -48,   -31,    51,   102,   248,   130,   176,    49,    13,   -51,    46,     5,     7,    -3,  -136,   -53,    -6,    -1,     6,   -14,   -14,   -20,    -7,    17,    33,   -23,   -28,   -41,   -36,    12,    -5,    22,   -19,  -201,   -97,   -29,   -20,   -60,   -50,  -127,  -163,  -114,   -93,   -19,    12,   -13,    20),
		    86 => (    2,     5,   -19,    14,    17,     0,     8,   -12,     1,     3,    12,    11,    68,    50,   -11,    -1,     6,    -7,   -11,     2,     8,   -11,     3,   -14,    12,    -9,   -19,     0,   -18,    -8,   -13,   -19,     7,     3,    61,    76,    68,    78,    83,    30,    94,    66,  -105,     6,   -14,    60,    49,    75,    99,    32,    21,   -10,   -18,    13,     7,    -8,    -4,   -18,    33,   -10,    46,    15,    75,    51,    84,   108,    62,    46,    90,    49,    37,     5,    62,    61,    93,   104,   170,   145,   105,    48,    18,    52,   -19,   -17,   -19,   -10,   -67,   -10,    15,    71,   135,   153,   140,   140,   163,   130,    77,   118,    82,   -28,    12,   106,    98,    -2,    36,   133,   151,   141,   102,   -36,    -6,    -8,     2,    14,  -138,   -66,    61,   135,   168,   114,    41,    99,   151,    82,   117,   -14,    34,   -49,    60,    82,    22,    51,   122,   -52,     5,    67,    60,    67,   -23,    43,   -10,    -4,   -88,   -80,    72,    90,    66,    83,   101,   119,   138,    46,    73,    -8,    20,    -6,    76,    38,   -73,   -53,    13,   -34,    61,    69,    75,   121,    44,    28,   -13,     3,    -1,   -30,    75,    23,   101,    36,    19,   116,   151,    41,   -42,   -47,   -43,   -30,    14,   -25,    36,    24,    24,   100,    32,    49,    52,    48,   -10,   -36,     4,    12,    -9,   -59,    35,    38,    15,   112,    75,   135,    64,    14,    -3,   -58,   -10,   -52,     0,    32,   127,    26,    86,    37,   -26,   -65,    38,    -9,   -50,   -92,    -8,   -10,   -62,   -92,    91,    32,   -27,    36,    62,    65,    63,     1,    31,   -58,    31,   -41,   -72,   125,   -62,    35,    69,   126,   -98,  -124,  -133,  -185,  -116,  -157,     8,   -17,   -93,  -102,    33,   -17,   -38,    11,    48,    -6,     5,    40,    24,   -22,    -2,   -50,   -81,  -133,   -84,    50,    58,   -37,  -117,   -98,   -32,  -157,   -59,  -138,     7,     4,   -76,  -119,    24,   -54,   -49,   -49,   -35,    11,    16,   -50,    35,     9,    16,   -99,  -120,  -138,   -80,    45,     0,   -65,  -135,  -128,  -132,   -44,   -65,  -198,    -1,    -6,   -72,  -152,   -14,   -11,    -5,   -74,  -122,   -49,   -23,    37,    49,   -31,   -79,   -64,   -48,   -41,    45,    47,    -2,   -54,   -92,   -55,   -77,   -46,  -148,   -57,    -8,     3,   -15,   -98,   -24,    15,   -35,   -86,  -191,   -14,    -8,    18,    -2,   -24,   -40,    -5,    55,   151,   125,    34,   -46,    25,   -69,   114,    41,   -52,  -149,   -54,    -9,     1,   -25,   -99,   -21,   -50,   -61,  -189,  -237,   -86,   -28,   -20,   -46,    24,   -46,    24,    80,   -41,   -19,    42,   -43,    38,    -7,   150,   -72,   -83,  -125,    -9,   -17,     2,   -20,  -109,   -97,   -42,  -121,  -114,  -146,   -80,    -9,    -1,    -3,   -21,     4,    39,    12,   -51,   -93,   -49,   -51,    -1,    49,   108,   -15,   -16,   -18,     2,    15,   -18,   -31,  -101,  -143,   -84,   -83,   -33,  -212,  -179,   -76,     3,   -21,   -33,   -53,    47,    35,   -81,   -67,    19,   -26,     5,    15,    -7,     1,    45,  -103,  -157,    15,   -21,   -50,  -181,   -29,    47,   -78,   -21,  -154,   -73,   -34,   -15,   -52,   -97,   -47,     8,    29,    -4,    28,   -13,   -20,    21,    13,    14,    36,    31,  -102,  -138,    -1,     0,   -45,  -156,    31,   -50,    -3,    27,   -14,    17,    38,    64,   -52,  -118,   -72,   -35,    18,   -15,    46,    11,   -15,   -39,    -7,    81,    95,    67,   -73,  -176,     3,   -15,   -30,  -195,   -28,   -61,   -20,    13,    19,    88,   125,   106,    60,   -31,   -17,    27,    30,    82,    84,    31,    66,    64,   -29,    49,    69,   104,   -75,   -83,    14,   -53,  -163,  -147,     0,   -47,    59,    75,    93,    16,   179,   162,   119,    27,    51,    -4,    -2,   -25,   -11,    35,    34,     5,   -11,   -19,     8,     0,   -56,   -34,    13,   -45,   -43,  -118,   -44,   -55,   -63,   156,   129,   135,   208,   168,   169,    93,   129,   134,    -8,   -73,   -19,   -86,    18,   -11,   -35,   -48,  -115,   -24,  -123,    -5,    19,    -2,  -111,   -54,   -59,  -109,   -62,   100,   293,   175,   139,    65,    97,    96,   116,    31,   -23,   -35,   -40,    62,    38,   -19,   -24,   -29,  -186,  -152,  -106,   -20,   -14,   -15,   -26,   -71,  -122,  -178,  -126,    12,    79,   135,   103,    84,    61,    11,    14,   -17,   -63,   -47,   -42,    -2,    51,    47,   -21,   -61,  -241,  -142,   -87,    -6,    20,     0,    -7,  -101,   -65,   -89,   -98,   -98,  -104,    -5,   -10,   -19,     4,   -18,   -18,    39,    39,  -103,   -35,    97,    61,   -29,  -102,  -165,  -194,   -67,   -71,   -20,    -3,    14,     8,     1,   -48,   -41,   -20,  -109,  -198,  -199,  -198,  -251,  -128,  -174,  -118,     3,   100,   130,    88,   -73,   -42,  -164,   -90,   -93,   -55,   -21,     9,    14,    13,     9,    -9,    12,   -19,   -61,   -83,  -140,  -100,   -73,   -86,     3,    65,    26,   -51,   -70,   -82,   -74,   -75,   -31,  -144,   -74,   -87,  -118,   -36,     4,    19,    -8,   -19,    -9,    -6,     0,   -36,   -48,    -8,     6,     1,    11,   -35,   -48,   -13,    19,   -28,   -37,    -1,    17,    -5,    -2,   -45,   -21,   -25,   -33,   -14,    -3,   -13,     3,    -8,   -11,    -2,    17,   -12,   -10,     8,     7,   -15,    -3,   -17,    22,   -12,     4,     1,     1,    -6,    15,   -23,    -3,   -14,   -24,    -7,    15,    13,   -11,    -9,    11),
		    87 => (    9,    -7,    12,     5,    11,   -10,   -16,     2,    15,   -15,    12,     4,    16,     2,    -4,     4,    14,    14,   -10,    10,     8,     8,     5,    11,    20,   -12,     5,   -19,    13,    -1,    -9,    15,     3,     6,   -17,   -14,     8,    -2,    -3,   -44,   -68,   -50,    -5,   -87,  -162,  -142,    -7,    -9,    -5,    11,    -5,   -21,     4,    17,   -14,    -7,     1,   -11,    10,     7,   -26,    -4,    11,   -15,   -18,   -27,   -97,  -174,   -26,   -20,    -3,  -125,   -46,   -58,   -46,   -26,    -2,   -14,    -7,    -6,    -4,    13,    14,    17,     9,    -2,    15,   -31,   -20,   -39,   -86,  -151,  -109,   -95,   -54,   -74,  -112,   -93,   -69,   -90,   -92,   -70,   -50,  -112,   -39,   -41,   -57,   -11,    -7,   -21,     3,    13,    13,    14,     1,     8,  -109,   -72,   -49,  -192,  -190,  -168,  -342,  -126,   -65,   -12,   -24,   -54,  -152,  -117,  -112,  -118,  -122,   102,     8,  -104,  -127,   -68,   -27,   -11,    17,   -18,     9,  -161,   -66,   150,    20,    95,    49,    72,   -69,  -180,  -199,    -4,   -74,  -123,   -66,  -122,  -155,   -80,   -62,   -47,   -74,  -182,   -75,  -112,   -11,     3,    16,    -9,    82,   112,    91,   146,   100,   103,    59,    75,   163,   -13,    11,  -100,   -93,  -105,   -49,   -22,   -81,     6,    -8,     4,    51,  -150,   -27,  -104,   -52,   -40,    -1,    28,   112,     2,   175,   163,   193,   229,    34,   205,   187,    84,    75,    50,    29,   -34,   -59,    -7,    28,     7,    22,    -6,   169,    38,   -29,  -109,   -28,   -56,   -68,   -25,     5,    18,    20,    75,    35,   152,    30,    99,    97,    81,   134,    29,    54,    49,     5,   -16,   -30,    16,   -11,   -14,   130,    -1,   -91,  -161,   -98,   -75,   -17,     4,   143,    67,    55,    10,     5,    53,    49,     6,     7,    31,   151,    83,   129,    60,    16,     5,   -22,     5,    37,     2,    81,    37,  -163,    23,   122,   240,   -12,   -66,    58,   -18,   -61,   -45,   -34,   -56,    37,     4,   -33,   -80,   -80,    12,   -22,   -11,    13,    73,    54,   -35,    45,   -62,   -50,   -50,   -59,    88,   120,   223,    14,   -41,    47,   -50,   -61,  -113,   -60,   -48,   -54,   -29,  -127,   -28,  -114,  -161,   -49,    -9,   -27,   -17,   -68,   -38,    15,   -94,     5,    36,  -122,  -157,  -115,    30,     4,    45,   -71,   -88,   -69,  -123,  -118,  -135,  -159,  -207,  -244,   -97,  -127,   -93,   -69,    35,    41,    -4,    21,    26,    18,   -28,   -67,   -77,  -280,   -36,  -137,    24,     3,     1,    37,  -105,  -191,   -75,   -67,  -102,  -114,   -88,  -112,   -85,   -43,   -82,   -35,    95,   -25,    37,    43,    -4,  -116,    67,   -52,   -11,  -143,   -88,  -112,   -61,   -23,    16,   -19,   -38,   -58,   -40,    -1,     0,   -66,   -56,    35,    15,    48,    30,    51,    40,   -66,   104,    51,    95,   -10,    66,   -12,    43,    13,   -93,   -80,   -10,    13,   -10,   -20,     2,   -18,     1,    -5,   -31,   -95,   -17,   -58,   -31,    -5,    27,    13,    28,   -72,    59,    76,     5,  -100,   128,    -2,    56,   -18,   -85,   -27,   -70,    19,   -29,    -3,   -65,   -20,   -20,   -39,   -21,   -46,     2,    60,   -32,    43,    79,     0,   -16,   -13,   -14,    33,    12,    39,    13,   -34,   -68,    20,  -189,  -143,   -22,    -3,    18,  -115,  -109,  -123,   -79,    65,    76,    14,    80,    92,    28,    48,     1,    -1,   -28,    42,   -24,   -92,   -40,    36,     5,    15,   -21,    12,   -77,    33,   -87,    21,     8,   -17,   -63,   -84,   -11,   -61,    82,    11,    15,    18,    -7,     0,   -12,   -50,   -59,   -74,   -34,   -88,   -43,   -16,  -103,   -33,   -31,   -48,   -92,    73,   -85,    -4,    16,   -19,   -14,   -76,  -125,   -36,    14,    13,   -16,   -77,    16,   -13,    23,    12,   -40,   -90,   -61,  -163,   -90,  -112,  -171,   -71,   -20,   101,   -19,  -107,   -46,   -17,    74,   -25,   -62,  -205,  -175,   -89,    -1,    22,   -21,   -71,    28,   -18,     5,   -26,   -68,   -42,  -179,  -205,  -130,  -120,  -133,  -174,    10,    18,  -136,  -114,   -17,   -14,   -18,   -45,  -137,   -79,   -92,  -106,  -178,  -133,  -108,   -44,   -49,     6,    14,   -48,   -53,   -67,  -128,  -157,  -116,  -143,   -99,  -140,     1,   -18,   -62,   -24,     8,   -27,   -14,   -31,  -179,     9,   -38,   -56,   -28,  -145,  -118,   -26,   -18,   -20,   -48,   -86,     7,   -26,     7,   -69,   -52,   -98,  -291,  -232,  -154,   -82,   -21,  -114,   -18,   -15,    -9,   -62,  -219,   -26,    -7,    30,    44,  -146,   -59,    -3,   -13,    13,    -3,    -5,    13,   -42,   -16,  -136,   -46,   -89,  -119,  -217,   -94,   -88,   -46,  -112,    11,    -2,     3,    43,   -19,    59,    63,   -24,   -33,   -27,   -58,  -103,    -1,   -22,    12,   -10,   -34,   -70,    81,   -92,   -38,    35,    46,  -119,   -91,   -79,   -30,   -23,     5,     9,    11,   -57,    56,   -52,   -71,   -59,   135,    62,   -41,   -89,   -59,   -39,   -23,   -14,   -83,     1,    -7,   -30,     6,   -62,   -29,   -35,   -35,  -118,   -23,   -39,    20,    13,    15,   -19,   -73,  -257,  -191,  -222,   -61,    -7,   -52,   -78,  -132,   -94,   -34,     9,   106,     0,   -53,    -3,  -109,    14,   -18,   -41,   -73,   -13,     7,     3,    12,   -13,    14,    15,     2,     8,    18,    -2,   -44,    32,   101,   125,    85,   -26,   -51,   -71,    82,    96,   133,   113,   -27,   -13,   -12,   -55,     5,    -8,   -13,     2,   -15),
		    88 => (   -8,    -9,     6,    -8,   -13,     4,   -20,    19,   -11,    -6,    18,    14,    15,    11,     9,    11,   -14,     6,    12,     7,   -15,    18,    -9,    -3,    13,    18,    -1,    -6,   -10,    -6,   -19,    -5,   -10,    -1,   -16,     4,   -13,   -17,   -17,   -35,   -55,   -49,   -82,  -202,  -217,  -180,   -36,   -32,   -39,   -24,   -35,    -8,     7,    10,   -19,   -16,     3,    17,    -5,    -2,     3,    -1,   -38,   -13,   -80,   -77,  -106,  -125,   -83,   -44,    -5,  -102,  -133,    41,    60,    -5,   -85,  -123,  -133,   -15,   -24,   -32,   -11,    -4,     4,    10,   -15,   -45,   -37,  -162,  -134,  -169,  -109,   -60,    39,    54,    68,    14,   -21,   -99,  -142,  -196,   -92,   -31,    32,    79,     9,    45,    48,   -50,   -22,    13,   -17,     9,    25,    -7,   -83,  -177,  -125,  -126,    67,    38,   141,   140,    24,  -134,    -3,   -63,   -61,    18,    -6,   -83,   -65,    18,   -81,    26,    53,    49,    31,   -36,     1,   -12,   -61,   -53,  -159,  -138,  -149,     9,   -50,    46,   105,    85,    23,    68,    14,    77,    85,   111,    45,     2,    -6,   -40,  -120,  -101,    60,    24,   -54,   -74,    14,    18,  -127,  -119,    33,  -108,  -145,   -88,   -13,   -23,    38,    23,   -39,    -7,    53,    80,    74,    29,    45,   -70,   -32,    -2,    46,    39,    14,    56,    -6,   -22,     5,  -121,   -68,    30,    65,   -54,   -84,   -10,    31,    47,    12,    -4,   -29,   -18,     5,   118,   119,    39,   -15,   -48,    41,    41,    92,   115,    46,    26,    14,   -82,   -64,   -83,   -66,   162,    85,     5,    40,    45,   -89,    19,    45,     0,   -17,    20,    24,    57,    51,    32,    36,   -25,   -24,   -53,    -4,    62,   -35,    39,    61,    16,    13,   -59,   -92,    92,   177,     1,    10,   -54,   -36,    20,    14,   -65,   -33,   -43,    10,    49,   -19,   -62,   -16,    25,     6,    -7,   -50,    11,   -16,   118,   168,  -124,   -20,   -58,  -124,   -77,    88,   -10,   -24,    -2,   -70,   -89,   -83,   -96,   -50,    64,    72,   -32,  -146,  -105,   -83,   -62,   -12,   -60,    36,    40,    57,    44,   121,  -104,    18,   -32,   -91,   -44,    62,    -9,    56,   -33,   -53,   -36,  -125,   -63,   -12,    57,     0,  -173,  -162,   -98,   -71,   -22,   -39,   -28,   -38,    95,    32,   -80,    68,   -93,     6,   -12,   -18,    22,   -87,    -8,  -114,  -141,   -81,   -89,   -26,    64,    68,    44,    49,     4,   -61,   -95,   -38,   -50,    22,     8,    45,    -3,   -70,  -211,  -233,  -129,   -15,    -5,     4,   -48,  -105,   -57,   -98,   -82,   -49,   114,   113,    96,   139,    72,     3,    39,    -6,   -46,    16,   -38,    43,    99,    55,    15,  -138,  -186,  -175,    13,   -32,   -16,   -31,   -73,   -98,    -8,    37,   -46,    49,   133,   136,   161,   125,    83,    14,    44,   -12,   -35,     1,    71,    85,    81,   -27,   -83,   -75,    14,   -95,   -45,   -24,    -7,   -47,   -21,  -117,   -21,    99,    98,   108,   172,   200,   104,    85,   115,    43,    19,    28,     6,    58,    57,    73,    36,    39,   -97,   -84,   137,  -156,   -51,   -16,     0,   -59,   -58,   -88,   -59,   -28,    81,    39,   132,   158,   141,    48,   -13,   -12,    -7,    71,   148,   134,    31,    91,    58,     2,    -9,    -1,    66,  -202,   -72,   -16,   -24,   -95,   -55,    16,   -96,  -112,     1,    13,    15,    55,    17,   -36,   -63,   -25,    87,     6,    25,    52,    46,    17,   -22,   -25,    31,    41,   -49,   -22,   -89,   -17,   -37,  -100,  -152,   -75,  -101,   -38,   -70,   -61,    -8,   -39,   -76,   -75,   -23,    68,   -17,    -1,   -74,    16,   -41,  -125,  -111,   -39,    61,   -29,  -121,   -12,   -37,     8,     8,   -52,  -182,   -89,  -153,  -133,  -137,  -122,  -106,   -65,   -74,    11,    74,    87,    31,    72,   -37,   -38,   -82,   -69,    -7,    47,    19,   -61,  -150,   -87,   -60,   -18,    -2,   -83,  -171,   -95,   -86,   -81,   -19,     5,   -97,   -52,   -53,    63,    80,   135,    90,    45,    23,   -63,     7,    38,    24,     9,    -3,  -137,  -118,  -112,    -8,   -41,   -44,  -103,   -32,   -77,    -1,    15,   -14,    -2,    -7,   -54,    92,   219,    89,    65,   122,    80,    71,   -12,     4,    30,   -75,   -47,    -4,   -77,   -61,  -115,   -17,   -40,   -35,   -50,     5,    84,    41,   -16,   -50,   -60,    11,    18,   107,    58,    37,   163,   133,    44,   -17,   -16,   -68,    41,   -51,    36,    53,   -49,  -112,  -110,   -29,   -15,    -8,   -29,   -11,    44,    21,   -45,   -93,   -54,    83,   100,    10,    71,   163,   115,    85,    48,   -62,   -20,    -1,    71,    12,    54,    72,  -159,  -131,   -71,    -3,     3,    12,   -56,   -45,   -32,   -66,   -72,  -101,   -70,    12,   -17,    34,   136,   180,   121,    12,   -29,   -71,    23,   153,   121,    27,  -111,   -57,  -184,   -91,   -43,    -4,    -7,     0,   -55,   -10,  -200,  -137,    -7,   -59,  -128,  -131,   -19,    89,    81,   111,    40,    25,  -124,   -47,    11,    25,   -69,  -181,  -175,  -111,   -97,   -38,   -69,   -15,    14,    -1,     9,   -81,   -71,   -78,  -130,   -95,   103,    62,   -72,   -37,   -23,    44,   -15,  -165,   -80,   -55,  -109,  -113,  -216,  -170,   -87,   -64,   -19,    -5,     6,   -12,     1,    -8,     6,     4,     0,   -31,   -25,    -3,  -105,  -145,   -79,   -23,   -26,   -91,  -171,  -122,  -128,  -107,   -63,   -37,   -13,    -6,   -32,   -13,    16,    16,    -2,   -11),
		    89 => (    2,   -17,    11,    13,   -14,     3,    16,    -9,     8,     0,     3,     3,   -14,     7,     9,   -15,    19,   -18,     1,     4,    -3,     1,     1,    14,     7,    18,     8,    -8,    12,    10,    20,    14,    12,    -6,     2,    -9,    -3,    13,    -4,   -49,   -98,   -65,    -4,    -8,   -27,   -10,   -71,   -57,     7,   -30,   -23,    -1,    19,     0,    12,     9,    13,     8,   -14,   -82,   -38,    -1,    -6,   -33,   -25,    -4,   -23,   -74,    -3,   -23,  -110,   -46,   -34,   -27,   -41,   -43,   -57,   -28,   -29,    -7,   -24,    -1,     0,   -18,    -2,    20,    17,   -46,   -78,   -93,   -78,   -95,   -25,   -39,   -10,   -59,   -53,   -81,  -112,   -95,   -80,   -83,  -132,   -84,   -55,   -52,   -47,   -14,   -14,   -19,     4,    16,    -5,    18,   -12,   -17,   -51,   -20,  -107,    18,   -64,   -31,   -38,   -91,  -153,  -120,   -75,   -69,   -32,   -33,   -74,  -128,  -148,   -72,   -41,   -35,   -11,   -98,   -19,    15,   -10,     7,    10,   -43,     5,   -12,   -25,   -41,   -44,   -61,  -142,   -52,   -54,   -52,    -4,   -17,     9,   -56,   -32,   -69,    -8,   -24,   -81,   -51,   -11,   -37,   -44,   -12,     6,    -2,   -20,   -57,    -1,   -24,   -84,   -79,  -184,   -87,   -65,   -73,   -39,    44,   133,    78,    43,    56,     1,    10,    41,    -2,   -63,   -72,   -37,   -66,   -28,   -39,     7,    -1,   -43,    -2,   -56,  -109,  -142,  -131,  -191,   -10,   -37,    50,    54,    -4,   -37,    57,    -7,    -2,   -40,    -9,   -13,   -22,   -67,   -59,  -109,   -45,    -7,   -32,   -61,   -50,   -21,   -66,   -20,  -123,   -93,  -193,   -66,   -84,    44,    -2,   -51,    -4,    -2,  -165,   -63,    -8,   -19,   -20,    13,   -69,   -50,  -103,  -156,   -42,   -29,    -1,     9,    -8,   -30,   -52,  -121,  -147,   -92,  -140,     3,    39,   -10,    50,   -27,   -32,    25,   -80,   -81,   -30,    89,    33,    25,   -79,   -61,   -32,   -62,  -148,   -12,   -64,    16,   -37,   -66,     4,   -21,   -45,   -73,    40,    36,    15,   -93,   -62,  -144,  -111,   -60,   -75,  -139,   -88,    86,     8,   -22,  -112,   -45,     5,   -73,   -16,   -21,   -51,     4,  -133,   -13,    57,   -13,   -55,   -51,   -13,    34,   -27,   -65,  -175,  -103,   -18,   -41,   -69,   -78,     3,   -52,     0,    -8,   -42,   -24,    57,   -89,   -38,   -18,   -57,   -18,   -24,    16,    47,    26,    27,    17,   -11,    70,   -40,   -71,  -146,   -37,   -94,  -152,   -94,   -56,   -42,  -110,   -19,     3,    51,    -5,    21,  -173,   -70,   -17,   -27,   -16,   -85,   -65,    87,    79,    37,    19,     3,   -23,  -118,   -67,   -79,  -133,  -105,   -41,   -27,    34,  -101,  -107,   -16,   -16,    58,     2,   -57,  -121,   -74,   -27,   -12,   -20,   -65,   -95,   -10,    48,    30,    29,    20,    87,  -111,   -51,  -172,  -124,   -80,   -55,    36,    14,   -61,    51,    50,     3,    13,    29,  -136,   -84,   -49,    26,   -14,    -2,   -12,   -86,   -26,     8,     6,    61,    42,    46,   -90,   -40,  -165,  -141,  -134,   -72,   -59,   -69,  -107,    41,    37,    85,    31,    16,  -202,  -144,   -37,    16,    -8,    17,    -8,   -95,   -70,    46,   -58,    92,    -6,    11,   -41,    50,   -36,     3,   -36,   -75,   -99,  -119,   -60,   101,    39,    57,   -45,   -28,  -158,   -66,   -73,   -10,     7,     7,   -11,   -73,   -65,    67,   -67,    -1,    78,   -72,    -3,   -17,   -18,   -23,  -101,   -41,    -7,     7,     1,    38,    27,    42,   -46,   -31,   -91,   -23,   -30,   -62,   -25,     2,    13,   -77,   -40,    67,    55,    48,   -12,   -49,   -13,   101,    40,    65,    14,    32,   -40,   -56,    48,    66,    23,   -39,    25,    43,   -71,  -145,    -3,   -75,   -58,   -13,    -4,   -48,   -27,    29,   132,   100,   157,   -46,    14,    94,   198,    47,   -22,   -59,   -13,   -14,     9,    86,   -60,   -20,   -41,   -20,   -79,   -50,    37,   -81,   -11,     9,   -23,   -30,   -37,    -8,    56,    30,   -19,    20,    36,   -12,    -2,   -12,   -60,  -134,   -61,   -44,    36,    98,   -45,   -32,     8,   -21,   -30,   108,    42,   -76,    -1,    10,    14,   -76,   -49,  -111,   -33,    18,    71,    42,     9,    -6,   -23,   -56,   -53,   -46,    -2,    14,    -7,    48,    16,    28,   -74,     2,     9,   131,   -28,  -152,    19,   -12,    12,   -28,   -40,   -68,   -65,   -81,   -81,    -7,   -14,   -51,   -84,   -34,   -96,    59,    21,   -25,   -21,    -3,    12,    27,   -13,    45,   -24,   104,    26,  -118,     4,    -6,    -6,   -17,    24,   -68,   -77,   -69,   -98,   -97,  -169,  -182,  -164,  -136,   -29,    35,    84,   -66,   -28,   -73,    58,    16,    45,   134,   -11,   116,    40,   -72,    -5,     8,     2,   -36,    10,    -8,   -15,   -38,   -24,   -60,   -80,  -156,  -142,   -32,   111,   -24,    -5,    -2,   -38,    18,    48,    79,    94,   127,    88,    97,    36,    -6,    12,    -8,   -13,    67,   -47,   -44,    19,   -17,   -53,   -49,   -78,    -2,    25,    76,   106,   -10,   -63,   -80,  -102,   -28,   124,   152,    98,   156,    72,    61,   -31,   -36,     9,     3,    10,     9,    23,    44,     8,    -2,    14,    -7,   -10,    -6,   -12,   -36,   -76,   -42,  -138,  -175,   -91,   -19,    16,   115,    68,    49,    58,   -10,    -2,    16,    19,    -4,   -11,    -2,    17,   -33,   -10,    -4,     3,     3,     6,    16,    15,   -11,    -7,   -52,   -23,   -67,  -113,   -79,   -77,   -47,   -66,     8,   -26,     9,     0,     3,    11),
		    90 => (  -19,     6,   -11,     8,     8,    -8,   -15,     7,    -3,    -9,    11,     8,     3,    16,     3,   -15,   -13,    17,   -20,    15,     3,    -4,     6,     2,   -15,    16,     7,   -18,   -15,    -1,   -11,    19,    -2,     8,   -14,   -11,   -13,     2,   -15,   -16,    18,    15,   -26,   -15,    -2,    11,     3,    13,    -3,     2,   -20,    -2,    19,     5,    -2,   -10,    11,   -15,     3,    21,    -4,     6,   -42,   -22,   -30,   -44,   -41,   -25,   -37,   -52,   -37,   -18,    -8,    12,    -6,   -21,    -8,     1,   -10,   -28,   -22,     8,     2,     0,     0,   -16,     2,    18,   -24,     4,   -23,    -1,    12,   -18,   -25,   -41,   -71,   -32,   -22,   -23,    18,    43,    40,     2,     1,     4,   -20,   -34,    21,    15,    -3,    -2,    16,    -7,    16,   -29,   -25,   -73,   -51,    29,    14,     6,    -9,   -57,   -37,   -38,   -29,   -25,    52,    68,    29,    61,    58,     2,   -11,   -22,    -4,   -17,   -23,    12,    20,    10,   -17,    13,    -6,   -19,    18,   -65,   -24,   -36,   -37,   -18,     8,    12,   -29,   -25,     4,   -27,     6,    80,    79,     9,   -23,   -22,   -20,   -19,   -15,   -56,    20,    -6,   -32,   -29,   -18,   -48,    18,    30,    11,   -39,   -32,   -11,   -25,   -43,   -21,   -37,    43,    17,     5,    34,    56,    37,   -24,   -25,   -29,   -84,   -19,     3,     7,   -25,   -40,   -43,    -8,    24,    63,    12,   -33,    31,    27,    14,    29,    18,     1,    74,    20,    45,    93,    26,     4,    21,    57,    -3,   -15,    -1,   -49,     6,     4,   -16,    44,   -39,    33,    37,    25,    51,    25,   -50,   -34,    12,    45,   -39,   -12,   -33,     5,    34,    14,    29,    71,    64,    37,    40,   -28,   -21,   -42,   -30,   -18,     2,    21,    -9,    93,    13,   -25,    -5,    28,    33,   -25,   -97,  -106,   -83,   -77,   -81,   -38,   -18,    -8,     1,     6,    84,    49,   -18,    24,   -29,    -4,   -14,    11,     9,     9,     2,    -7,    75,    69,    62,    52,     8,   -93,   -77,   -89,   -62,   -44,     7,   -87,   -58,   -59,   -32,   -39,   -47,    60,    14,   -18,   -30,   -43,    -5,    16,    60,    10,   -20,    48,    80,    34,   -45,     9,   -82,   -97,  -132,  -103,     5,    21,    26,   -49,   -55,   -86,  -125,  -105,   -61,     5,    10,    68,     3,    -8,    -9,   -11,    -6,    13,   -20,    55,    38,    22,   -31,   -12,   -68,  -111,  -133,   -85,     5,   -17,   -33,  -123,  -143,   -87,   -92,   -95,   -39,    -4,   -23,    39,    32,   -15,    19,    19,   -13,     6,    10,    93,    14,    82,   -41,   -48,  -100,  -148,  -151,   -73,   -40,   -16,   -51,  -113,   -90,  -109,  -104,  -101,   -50,     8,    44,    44,    14,     3,   -30,    11,    -5,    -6,   -61,   104,    65,   -23,   -78,  -109,  -126,  -109,   -95,   -92,   -74,   -44,  -105,   -93,   -81,   -88,   -94,   -91,   -45,   -62,   -22,   -48,    30,   -30,   -13,   -15,    14,    -3,     9,    92,    42,   -16,   -56,   -73,  -109,   -88,   -94,   -51,   -50,   -53,   -17,   -42,   -78,   -68,   -81,   -88,   -41,    10,    -5,   -31,     9,   -25,    -1,    13,     7,   -36,    -6,    53,    72,    50,   -11,   -36,   -53,   -62,   -55,   -69,   -54,    46,   -41,   -40,  -121,  -118,  -113,   -46,   -81,   -21,    80,     2,    32,   -48,    22,    10,   -11,   -36,    44,    81,    61,    64,    64,   -42,   -54,    13,    -5,   -41,   -49,   -34,   -64,  -122,  -120,  -119,  -105,   -68,     4,    47,   -10,   -16,    30,  -109,    18,     9,    -7,   -19,    -9,   118,    36,    34,    61,   -15,   -17,    -4,   -44,   -21,   -36,   -98,   -44,   -95,   -99,  -139,   -82,   -41,    40,     6,    24,     8,   -18,   -23,   -12,    18,     5,    18,    -5,    75,     7,    17,    33,   -16,     6,    22,   -18,     1,   -30,   -32,   -49,   -72,   -28,   -31,   -10,    46,    -1,     6,   -36,     9,   -66,   -34,     8,   -19,     1,    16,    -1,    58,   -28,    57,    32,    11,   -50,   -33,    19,   -36,     6,    22,    -6,    41,    49,   -57,   -15,    12,   -12,    33,   -25,    -7,   -49,    -9,     0,     9,     4,   -25,     0,     3,   -65,     7,    78,     5,     6,   -17,    35,   -35,     1,    -9,    -4,   -38,    14,     7,    38,    26,    14,   -44,    -2,   -38,    -3,    18,    22,    18,    -8,   -11,   -33,   -42,   -25,   -57,    60,    22,   -22,    12,    28,   -29,     9,   -20,   -42,    40,    46,    -7,    17,    17,   -33,   -21,   -29,   -49,     5,    22,    24,    20,    -6,    -6,   -38,   -24,   -30,    26,    52,   -19,   -38,   -12,     0,    18,   -44,   -18,    -8,   -47,    -9,   -33,    19,    -4,     2,    -2,   -47,   -65,   -51,   -47,    -9,   -11,   -12,   -20,   -17,   -32,   -16,    72,    54,    37,   -42,    -6,   -13,   -38,    20,    44,    34,    11,    23,    34,   -29,   -35,     2,   -11,   -23,    -1,     1,   -11,    15,   -15,     6,     9,     0,   -22,   -15,    44,    82,    82,    19,     4,    -2,   -33,   -29,   -56,     5,    -3,   -34,   -89,  -117,  -103,   -72,   -67,   -43,   -10,   -14,    -8,    -5,    11,    18,    12,    -2,    -6,   -45,   -69,    -1,   -20,    -2,   -22,    -6,     8,   -45,   -43,   -32,   -53,  -154,   -85,   -83,   -87,   -58,   -24,   -63,    -1,   -15,    12,   -12,    16,     1,   -13,    -1,     8,    -7,    -2,    -8,     3,   -17,     0,    -7,    17,   -28,   -24,    -8,    -5,    -4,     0,   -19,     8,   -40,   -53,   -49,    -2,    -6,     0,   -19),
		    91 => (   -8,    -2,    12,    -7,    12,    -8,   -14,    -6,    13,     6,    -4,     8,    18,   -10,    -6,    19,    20,    15,    18,    -8,   -15,    -6,     9,    14,     9,    14,    17,   -13,    -6,     8,    -3,    10,    -6,    20,    -4,    -1,    10,    -4,    -7,   -10,    -8,   -36,   103,    51,    60,   -66,   -19,    -3,   -12,    -9,   -14,     1,   -13,     5,    -1,    13,   -10,    17,   -13,    11,    15,   -19,     7,    17,   -64,   -68,   -49,   -56,   -19,    37,    36,    73,   167,   101,    90,    33,    51,  -109,   -82,  -102,    -9,    -1,   -19,    -2,    -1,   -13,   126,    61,   -12,   -64,  -115,    70,    19,    17,   -88,  -144,   -63,    -5,   -13,     9,    31,     4,    14,   -89,   -28,   -65,   -56,   -67,   -53,   -10,    -3,    -9,    11,    -7,   122,   115,   100,     7,   -33,    42,    83,    72,    41,    11,   -93,    19,   -31,    35,   -19,    -7,    -7,   -92,   -98,   -47,    90,    73,    65,   -44,   -34,   -51,    -5,   -18,    47,    34,   137,   114,    19,    22,    79,    12,   -21,   -16,   -39,   -45,   -92,   -23,   -24,   -30,   -46,   -35,  -108,    36,    93,   121,    96,   -80,   -43,   -67,   -19,   -15,   -59,     5,   137,    53,    42,   -10,   -84,   -65,   -22,   -31,    38,   -46,   -28,   -66,   -86,   -60,   -44,  -156,   -47,    58,   105,    94,    31,    -6,   -28,   -28,    14,    -5,   -69,   -79,   -71,   -57,   -82,    48,  -152,   -33,   141,   104,    87,   -22,    25,   -56,  -124,   -62,   -30,  -105,   -30,    75,   104,   117,    23,   -55,   -77,   -27,   -18,     3,   -88,   -61,   -71,   -73,   -68,    94,  -126,   -33,   127,    -9,    84,    -5,   -35,   -45,   -60,  -102,   -90,   -91,    49,    55,    55,    18,    17,   -41,   -87,   -35,     2,    -4,   -81,     1,   -60,   -78,   -49,   114,   -40,    19,    55,    -6,   -66,   -85,   -66,   -50,   -87,  -160,   -93,  -132,    15,     9,    49,    40,    13,   -19,   -76,   -40,   -13,   -12,   -55,    -4,   -55,   -38,   -78,    41,    30,   -52,    86,    12,     9,    -4,   -21,   -54,  -130,  -116,   -27,   -33,    -1,     7,    49,    75,   -47,    -9,    17,    38,   -18,    10,    -8,    -1,     3,   -59,  -110,    48,   -78,   -30,    -9,   -48,   -23,   -52,    56,     3,  -104,   -37,   -26,   -33,   -27,   -54,    68,    39,   -46,    10,     1,    94,   -19,    15,   -58,    -1,    17,   -38,   -46,   -55,  -104,   -86,     6,     0,   -30,   -59,    27,   -32,   -34,   -24,   -16,   -33,   -38,   -59,     5,    23,   -75,    29,    56,   107,    10,    -9,   -43,    -5,   -23,   -43,   -11,   -17,     7,   -24,   -31,   -47,    20,   -44,     4,    11,   -56,   -35,   -91,   -39,   -63,   -80,   -70,  -159,   -77,    71,    20,    17,    -4,    17,    23,    24,   -33,   -66,    20,   -33,   -41,   -68,  -136,  -185,   -63,    57,    41,    42,     5,   -20,   -28,  -123,   -93,  -108,  -122,   -67,   -45,   -87,    -5,     5,    14,     7,    -9,    -7,   -42,  -136,   -68,   -67,   -92,  -140,  -209,  -177,   -63,    35,    76,   -62,   -82,    30,    11,  -100,  -115,   -56,  -113,   -62,  -145,  -126,  -105,   -26,     9,   -17,    -1,    -7,   -44,   -30,   -63,   -70,   -95,   -18,   -82,   -57,   -90,   -28,    95,    23,   -43,    28,    21,   -34,   -29,   -11,     0,   -51,    91,  -132,  -100,   -26,    20,    -4,   -10,   -27,   -15,   -15,   -27,   -44,    15,     5,    48,    18,   -68,   -26,    61,   -15,    46,   -41,    34,    16,    64,    55,    51,   -16,     1,   -99,   -70,   -68,    12,   -20,   -12,   -71,   -45,     7,   -82,    -5,    53,   103,    60,   -90,  -108,   -75,    33,    15,    18,    69,    15,    27,   -62,   -25,    30,     3,    23,    -6,   -64,     3,   -19,     2,    42,   -69,   -42,   -12,   117,   130,   163,   149,   119,    18,  -119,    -6,   -18,    53,    81,    10,    26,   -55,    -8,     6,    75,   173,    56,    51,   -66,   -27,    17,     5,    -7,   -37,    41,    81,   118,   136,    89,    81,    67,    -4,   -46,   -14,    43,     0,    49,     6,    12,    24,   107,    97,   120,    67,    40,     4,   -47,   -11,    32,    39,   -17,   -13,   -41,   -85,   -48,    -3,   -12,   -42,   -46,   -91,   -25,    17,   -65,     7,   -80,   -50,     9,    44,    42,   -15,    58,    21,    -6,    62,   -31,    -5,    58,    25,   -53,   -35,   -36,    67,   -11,   -41,  -108,   -91,   -85,  -109,    18,    14,    -6,    33,   -82,   -31,   -13,    -8,     9,    -2,   -91,   -62,   -19,    -1,    21,   -15,   -18,   -15,   -18,   -42,    18,    83,   104,    44,   -11,   -15,    22,     6,    87,    22,   -68,   -67,   -65,    46,   -38,   -29,    75,     9,   -41,   -58,   -53,   -72,    93,     0,    20,     6,    15,   -25,     2,    -2,    -1,   -34,   -34,   -36,    19,    19,   -23,     6,   -65,  -136,   -59,   -74,   -44,  -116,   -10,  -106,   -41,   -42,   -93,    61,    84,    11,   -16,    -3,    -2,   -38,   -30,   -47,   -13,   -42,   -57,   -33,   -60,   -21,    -3,    70,    75,   -49,  -108,   -74,   -75,   -79,  -141,   -97,   -44,   -31,    13,     5,    -9,     2,   -12,    -7,     6,   -33,   -33,   -88,   -83,   -58,   -31,   -29,   -21,    -3,   -25,   -60,   -80,   -59,   -51,   -75,   -13,   -16,   -29,   -34,   -20,   -14,    15,    14,     9,     8,     7,   -16,     4,    12,   -17,     5,   -16,     0,   -11,    15,   -34,   -61,    15,   -15,   -19,     6,   -10,    13,   -11,   -17,    -2,     0,    -2,    -5,    -2,     7,     5,    -7),
		    92 => (   15,    19,    19,    14,     7,    -1,   -11,   -14,    -6,   -14,    19,   -18,   -20,   -24,    37,    35,    19,   -13,   -16,    -7,     3,     0,   -16,   -10,     7,     3,   -11,     6,   -13,    13,    -6,     9,    -8,    16,   -20,    23,   -31,   -65,   -89,  -128,   -26,   -36,   -15,    53,    72,     5,   -55,  -157,  -100,  -107,   -74,   -16,    19,   -16,    -1,    14,    10,   -14,   -10,   -48,   -53,     4,    20,     8,    10,   131,   128,   149,    12,    42,   112,   183,   152,    67,   -67,  -141,   -76,   -32,   -75,   -22,    -8,     2,    19,    17,   -13,    -3,     8,  -102,  -126,    57,    79,   104,    -3,   -90,  -136,  -177,  -228,     1,   -26,     1,    13,   -71,  -171,  -113,   -98,   -22,     6,  -109,  -119,    -9,   -20,     2,   -10,    -6,   -30,   -85,    -2,    43,   186,   147,   110,   182,    52,   -44,   -63,   -66,   -45,    26,   -55,   -17,    25,   -36,   -28,   -85,    10,   -86,  -144,   -11,   -96,   -31,     6,   -11,   -78,   -46,     0,   -79,   -66,    16,   112,    34,    87,     1,    27,    27,    44,    17,    -8,    17,    48,    63,    32,   101,   -36,   -61,  -125,    40,  -170,   -44,    -8,    -9,    14,     4,    40,   -19,   -16,   -24,    79,   -13,    22,   -85,    19,   -68,     5,    -1,    49,    30,    72,    30,    -9,    36,   -18,   -53,  -215,   -26,  -156,   -38,   -19,   -15,    61,     3,    76,   173,    50,    23,    51,   -16,  -116,   -59,    -7,    25,   -36,    27,    62,   -54,    18,   -26,    20,    97,    85,  -151,    32,    92,  -100,   -67,   -90,   104,    66,    24,   -15,   143,    54,   -32,    43,    31,   -35,    35,    33,     7,   -11,   -82,   -52,   -19,   -70,    18,     7,   -64,     5,    89,   -27,   -56,  -165,   -49,    12,   -71,    19,    78,  -100,    11,     8,   -48,     5,   -42,     1,    49,    59,    52,   -39,     0,   -34,   -15,     0,   -35,    -7,   -28,    82,   -15,   -74,  -219,   -29,   -36,    20,     9,   -41,    42,   -47,   101,   157,    22,    21,   -53,    93,   -34,     6,     8,   -28,     5,   -41,   105,   -56,   -65,   -15,    23,   -44,  -143,   -82,   -66,   -53,   -66,    -8,   -80,    13,    10,   -31,    45,    76,    57,    22,    49,    58,   -19,   -76,  -103,   -23,   -83,   -18,   -62,    -4,    29,    33,   -13,  -105,   -82,    37,    42,   -50,   -94,    -7,   -45,  -152,    -1,   -53,    13,   142,    70,    -3,    95,   -20,  -103,   -59,   -46,  -107,   -82,   -86,   -51,    59,   114,   -41,    94,    83,   -84,    99,    25,    -2,   -25,   -14,   -87,   -54,   -18,   -20,    65,   233,    74,   -37,    10,   -25,   -14,   -28,    25,   -91,   -66,   -83,   -27,    42,    74,   -18,    23,    85,   177,   134,   144,   152,   -23,    13,    -8,   -33,    16,    68,    82,   145,   158,   -86,    54,    14,  -130,   -61,   -86,   -64,   -40,   -33,    -8,   -12,    62,  -116,    52,   150,   263,   217,   112,    97,    45,    -2,   -59,   115,   130,    -5,    34,    72,    63,    94,    20,   -42,   -26,   -33,   -71,   -21,    -3,   -26,   -66,   -22,   -55,    33,    86,    83,    75,   -17,    84,   178,   142,    -7,    -8,   148,   136,   -86,   -66,    15,   141,    62,   143,    62,    13,    56,   -12,   -39,   -31,   -20,   -62,   -40,    29,   -36,   280,   227,   141,    30,   158,   192,   107,     1,   -26,   136,    94,   -29,   -50,    30,   -23,   -25,   -22,    16,     5,    10,    -6,    41,   -24,   -44,    -8,   -15,   -21,    82,   294,   163,    64,    47,    74,    75,    69,   -10,     2,    21,    51,   -33,   -23,    12,   -59,    33,   -37,   -55,     8,    25,    -8,   -92,   -49,   -71,   -95,   -12,    71,   255,   223,   172,   124,    97,    83,   -24,    37,     9,   -79,    30,   -35,    -6,    -7,   -48,     0,    43,    31,    49,    70,   -40,   -48,    16,    58,   -43,  -108,    44,   142,   161,   215,   150,    61,    -4,   -48,    31,   107,   -20,   -45,   134,   -68,   -24,    -6,    -8,     3,    -2,    58,    91,   104,     3,     0,   -79,    12,   -87,   -25,    51,   170,   211,   261,   106,    82,    39,    20,    17,   -16,   -13,    -9,   127,   -50,    81,   -22,    25,     0,    92,   147,    83,     2,    43,    41,   -85,    -2,   -21,   -84,   185,   295,   218,   190,   243,    35,   -38,    24,   -27,   -14,    -2,     1,   -42,   -92,   -31,    36,   -68,    -3,    80,    74,    30,    41,   -56,    -5,   -56,   -34,    10,    65,   248,   248,   225,   175,   168,    71,   -94,    40,   -15,   -11,   -18,    13,     4,  -120,    -7,    39,    61,    23,    33,   141,    63,    38,    26,    22,   -49,   -41,   161,   299,   240,   173,   237,   216,   158,    98,   -81,     5,     5,   -17,    12,    -1,  -100,   -40,   -77,  -138,    59,   -55,    -3,    70,    77,    35,  -124,  -197,   -31,    24,   185,   256,   339,   239,   140,   189,   141,   -37,    47,    14,    47,    -2,    17,    -5,   -39,   -19,  -115,  -218,    77,   -63,   -63,   -84,  -122,  -114,  -152,  -151,    23,    35,    27,   130,   214,    57,    12,    34,   -85,   -79,   -45,     1,    35,   -15,    19,    16,    15,   -17,   -30,   -60,  -137,  -204,   -98,  -225,  -266,  -202,  -184,  -270,  -268,  -213,  -213,  -200,  -163,  -259,   -77,   -45,   -95,    10,     6,    -1,     8,     5,     8,    16,   -18,    15,   -32,   -27,   -37,   -32,   -23,   -26,   -99,  -120,   -87,  -105,  -116,   -54,   -60,   -52,   -34,   -43,   -30,   -34,   -42,     6,   -17,     9,    12,    16),
		    93 => (   -4,    -2,   -10,    10,   -12,   -18,     9,     7,    12,    -9,     9,    -6,   -10,   -24,     5,   -10,    12,   -10,   -18,    16,    16,    19,     4,   -12,     9,   -16,    -4,    13,    18,   -19,    -2,    -3,    16,     6,    -4,    -9,    17,   -21,   -19,    -6,   -14,   -22,   -32,   -31,   -40,   -47,   -11,    -4,   -18,     3,     4,   -20,    10,    13,   -19,     8,     1,   -19,     1,    -2,    -7,   -19,    -4,     1,   -82,  -100,   118,    29,   -39,   -77,  -126,   -75,   -75,   -53,   -68,   -45,  -137,  -106,  -127,   -77,   -11,    -2,     8,   -18,    -6,    -4,    -9,   -11,     1,   -33,    18,    52,   -73,  -117,  -156,  -125,  -149,  -188,  -238,  -124,   -98,  -118,  -156,  -105,   -98,   -71,   -41,   -98,   -34,   -26,     7,     5,   -17,     5,    11,     3,    39,   113,   131,   -52,   -31,  -157,   -26,   -38,   -43,  -115,  -188,  -177,  -175,  -160,  -152,  -160,  -120,   -37,   -57,   -48,   -36,   -77,    -2,    19,    17,   -13,     4,    24,    53,   110,     9,   -42,   -16,    49,    96,    74,    72,   -37,   -58,   -34,   -57,   -49,  -117,  -165,  -105,   -95,  -100,   -40,   -24,  -102,   -34,    20,     7,    -3,     7,    69,    37,   -67,    31,    85,     2,    68,   -35,    50,    23,   -52,   -72,   -87,  -115,  -103,   -73,  -145,  -118,   -92,   -95,   -94,   -71,   -10,   -61,     7,    -7,    38,   -12,    62,    13,   -16,    86,    30,    56,   -15,   -21,   -89,    -7,    12,   -27,    50,   -83,  -122,  -170,  -190,  -118,  -112,   -82,   -95,   -67,   -14,   -47,   -23,    14,    15,   -63,    36,     1,    -8,   -28,   -81,   -22,   -18,   -97,    -1,   107,   115,   127,    84,   -24,  -166,  -197,  -204,  -155,   -68,   -84,   -96,   -64,   -35,   -36,    11,   -12,   -53,   -52,    11,   -27,    37,   -63,   -45,   -81,   -27,   -41,    77,   102,   112,   133,    11,   -84,  -229,  -212,  -210,  -140,   -78,   -60,   -28,   -49,   -64,   -53,   -16,    -3,   -88,   -37,   106,    13,    56,    -1,   -45,   -76,     4,    10,    50,    82,    69,    18,   -73,  -111,  -236,  -256,  -201,  -162,  -148,   -80,    -3,   -36,   -43,   -25,    -1,    -9,  -129,    -6,   138,    80,    17,   -22,    -5,   -27,    39,    61,    35,    62,    -3,   -66,   -78,   -85,  -111,   -94,  -133,  -102,  -139,  -110,   -39,    -9,   -94,   -58,     0,     5,   -98,  -117,    95,   -30,    -8,   -94,   -62,    48,    34,   104,    85,    76,    15,    13,    10,   -82,   -82,    31,     2,    -7,    55,   107,    74,   -76,   -60,   -38,   -16,     5,   -37,   -91,   105,    65,    21,    -9,   -40,    45,    75,    76,    65,    63,    53,    23,   -46,   -12,   -14,    32,    -9,   -28,    32,    60,    95,    91,   -81,   -53,     3,   -22,    40,   -10,    49,   -90,   -61,   -58,   -41,    22,    69,    35,   -16,   -18,     5,   -49,   -18,    27,   -50,    -9,    86,   -10,    13,    12,   171,    63,  -102,   -39,   -24,    -7,    48,     7,    26,  -100,   -83,   -64,   -10,    43,    11,   -38,   -75,   -63,   -65,   -13,   -68,     9,     8,    -4,    61,   111,    75,    67,    64,    16,   -85,   -14,    -4,    16,    16,    -2,     7,  -102,  -157,   -65,  -105,    22,    88,   -71,   -83,   -79,  -142,  -174,   -55,   -72,   -69,    -2,    31,    94,    97,    93,     8,   -15,   -67,   -64,   -32,    17,     3,   -21,    74,   -31,   -75,   -59,  -123,   -53,   -59,  -149,   -81,   -82,   -88,  -161,  -158,   -81,   -83,  -126,    54,    45,   140,    71,    49,   -12,   -56,   -27,   -11,   -16,   -10,    17,     8,     8,   -44,   -99,   -66,    -3,   -47,  -162,   -68,   -33,   -80,   -69,  -128,   -64,    -8,   -27,     7,    48,    69,    49,     5,    25,   -50,   -29,   -62,    19,     1,   -29,   -41,   -53,   -38,   -45,    38,   -10,   -29,   -72,   -43,    19,    44,    17,   -33,    18,    61,   -28,     0,    13,    35,    18,   -42,    31,   -13,   -84,   -45,    20,     3,   -40,   -83,   -59,   -73,   -97,    -2,    35,    41,   -31,    24,    29,    48,    68,    73,    95,    -5,   -43,   -27,    57,    57,    19,   -10,    44,   -34,   -25,   -16,   -18,    -7,     1,     7,    49,   -17,  -123,   -90,   -53,   -33,   -60,   -52,   -77,   -34,    18,     6,    11,   -33,   -69,    -7,    -1,   -81,   -29,    27,   -43,    -4,   -41,   -10,     5,    -6,     1,    -6,     4,   -17,  -111,  -107,  -107,   -96,   -62,   -84,     0,    -8,   -80,   -29,   -81,   -81,   -32,   -29,   -29,   -34,   -18,    32,   -55,   -42,     7,    13,    14,     9,    27,   -56,   -15,   -26,   -18,    -2,   -45,   -44,   -60,     2,    38,   -27,   -58,   -25,   -63,   -47,  -103,   -43,   -53,   -51,   -41,   -85,   -23,   -36,    -1,    -3,    12,     6,    41,   -29,   -57,   -44,    44,    64,    36,    -1,     3,   142,    25,   -55,   -16,   -27,   -73,  -104,   -62,   -23,   -67,     7,   -21,  -107,   -52,   -35,     8,     3,    17,     2,     9,   -79,    -7,   -31,    12,    39,    17,    -5,   -32,   -40,   -25,    52,    33,   -36,   -66,   -55,     6,   -20,  -141,   -92,   -87,  -125,    -5,    -7,     9,    17,     4,    17,    -3,   -40,   -38,   -49,   -43,   -53,  -101,   -92,   -35,   -84,   -61,     1,  -109,   -46,     8,     3,   -58,   -50,   -52,   -19,   -92,   -12,    16,     4,    -3,    14,     1,    -8,    -7,   -10,     7,   -11,   -13,    -4,   -14,   -44,   -29,   -48,   -46,   -72,   -51,   -97,   -11,    10,     3,   -73,   -37,   -46,   -27,    14,     3,    -4,    19,     7),
		    94 => (   -8,   -20,     8,    -9,     7,    16,     3,    -6,     9,    13,    20,   -14,   -33,   -13,   -35,   -25,    -6,   -12,   -10,   -18,    12,     8,     0,    16,   -13,     6,    -3,   -20,    17,    17,    -1,    13,     5,     1,   -37,   -77,   -17,   -72,   -72,   -79,   -82,   -70,   -17,  -100,   -94,   -49,     3,    -1,   -84,   -24,   -35,    -9,   -20,    -6,    -2,     5,     8,    -9,     7,  -104,  -156,   -36,   -77,  -110,   -58,   -81,  -140,  -221,  -148,   -96,  -139,   -61,   -17,   -49,   -98,   -93,  -101,   -17,   -74,   -66,   -98,   -48,   -20,     1,    -5,   -14,    -4,  -116,  -194,   -43,  -142,  -138,   -72,  -108,  -130,   -60,   -78,  -168,  -110,   -77,    57,   -74,  -114,    -1,   -23,    13,    21,    38,  -105,   -70,     9,    19,    16,    11,   -52,   -94,    14,   -57,  -118,    10,    12,   -39,  -117,   -13,    56,   -63,   -58,  -160,   -55,   -89,   -88,    92,    66,    53,    -7,   -59,  -111,    23,   -35,    -3,    -7,     2,   -53,  -107,  -111,   -57,   -80,   -10,    37,    24,   116,   -37,   -31,   -67,  -119,  -155,   -60,    24,   188,    37,    13,    32,   -65,   -68,  -110,    45,   -72,    11,     7,     0,   -20,   -20,   -61,   -58,   -18,    11,   -29,   -22,  -135,   -60,   -66,   -18,  -177,  -281,   -49,    14,    80,   109,   168,   163,   -78,   -48,   -81,   -64,   -19,   -57,    19,   -41,   -78,    -1,   -68,   -11,   -24,   103,   -24,   -73,  -109,    21,    74,   -49,  -220,  -196,   -28,    43,    77,    59,    49,    47,   -56,   -59,  -116,   -95,   -36,   -58,   -79,   -90,    74,    -7,   -42,    -2,    37,    54,   -65,  -101,   -81,    41,     6,   -88,  -135,  -103,  -101,   160,    20,    57,     2,   -93,   -98,  -133,  -110,   -47,   -92,   -45,    -4,   -83,    55,   -39,   -53,   -72,    12,   -16,   -46,   -30,  -123,   -11,   -37,   -29,   -82,  -142,   -10,    98,    45,   -25,     5,    76,    23,  -103,   -98,   -28,   -26,   -40,    -3,   -61,    68,    95,   -12,   -67,   -95,     8,    17,   -64,    44,     1,   -30,   -17,   -98,  -199,   -50,    68,    19,   -27,   -51,    66,   -75,  -165,  -146,   -24,    -5,   -35,    11,  -128,   -39,    75,   -85,     0,   -25,   -38,    52,    -4,    38,    60,    27,   -49,  -191,  -148,    11,    75,     8,   -12,   -67,  -142,  -134,  -135,  -211,   -85,   -22,   -90,    13,   -63,    31,    -9,   -74,     1,    88,    29,     5,   -16,    93,    37,    50,  -140,  -147,  -143,     3,    15,    23,   -24,   -87,  -119,  -124,    14,    45,    28,   -58,   -85,     4,   -64,   -22,   -23,   -31,     7,    96,    22,     4,    27,    58,    56,   -29,  -134,  -155,  -122,   -47,    40,    50,   -59,   -93,    21,    74,    66,   -64,   -42,   -98,    17,     9,     4,  -116,   -28,   128,    76,     2,    44,   -28,   102,   125,    91,   -15,   -40,   -41,   -90,    -7,    12,    30,    24,    26,    76,    -9,    15,   -33,   -91,   -79,    -6,     6,   -11,   172,    -5,   102,    30,   -24,   -27,    12,    23,    86,    57,    57,    12,   -63,  -100,   -33,   -12,   -22,    56,   -14,    54,   144,   -41,  -129,  -146,   -57,    15,    -3,   -16,     8,   -97,   -53,   -88,    32,     3,   -45,   -14,   -20,  -138,   -79,   -49,   -82,   -31,   -22,    12,    37,   -31,    75,    25,   -11,  -153,   -40,   -76,   -99,   -44,   -14,    17,    42,  -140,     4,   -20,     5,    50,    62,   -22,    -2,   -20,  -146,   -20,     6,    54,   -16,    30,    43,   -41,    19,    56,   -75,   -52,  -104,    59,   -17,   -63,   -44,    14,    44,   -81,    28,    58,    43,    80,    -2,   -22,   -45,   -56,  -145,   -26,    38,    95,   -15,    38,    22,    39,    84,    12,  -119,   -25,   -98,   -77,   -33,   -12,     9,   -15,   -85,     8,   -25,    20,    92,     2,    16,    17,   -11,  -164,  -162,   -47,   -25,   103,    15,   -65,    73,    46,    49,    76,   -75,   -55,   -93,  -127,    -3,   -16,    -8,     9,   -45,   -22,    20,   -51,     5,    34,    -5,   -64,  -116,   -30,   -16,    -1,     7,    19,     5,    48,    64,    64,    57,    81,   -87,   -27,    -8,   -44,    -7,    -3,   -14,     8,  -102,   -20,    15,   -27,    22,    38,    33,   -93,   -87,   -93,   -20,    -3,    -2,    24,   -44,    59,    42,    17,    61,    74,    64,   -50,    69,   -16,   -61,   -12,    16,    17,    -7,  -103,  -152,    58,    24,   -24,  -101,  -152,  -230,  -108,   -75,     1,   -18,   -32,   -43,   -69,    27,    57,    76,    93,    27,   -31,   -13,   124,    35,   -10,     0,     2,   -10,   -65,  -107,   -81,   -16,   -41,   -20,  -152,  -200,  -106,   -89,   -66,   -16,    -4,    52,   -83,     1,    53,    91,   145,   -84,   -59,    10,    36,    27,   -10,    17,    14,   -12,   -21,   -49,   -13,     0,   -18,   -59,   -96,  -118,  -107,   -58,   -18,   -96,   -53,     8,   -36,     4,   -33,    18,   -22,  -107,   -13,   -90,   -59,   -41,     6,   -11,    16,   -52,   -17,   -56,    -7,   -24,     6,   -42,  -100,  -140,   -54,     5,   -58,  -174,    -5,    24,   -26,   -99,  -183,   -91,  -126,  -155,   -74,  -105,   -76,   -50,    12,     0,   -13,    -2,   -19,   -78,     6,   -12,   -23,   -31,   -94,  -171,   -18,   -55,  -112,  -175,  -110,  -185,  -139,  -137,  -126,  -193,  -144,  -159,   -21,   -17,    14,    -9,    11,    16,   -16,    17,    12,   -20,     9,   -20,   -48,   -32,   -57,   -99,   -83,   -80,   -46,   -74,    11,  -107,  -142,   -94,   -74,   -82,   -54,   -90,   -33,    14,     2,     9,   -13),
		    95 => (   -8,     9,    11,    -5,    -9,     8,    14,     1,    15,    18,    -7,   -14,    12,   -10,    -4,     2,    -5,   -15,     0,     9,   -10,   -19,   -12,     6,   -16,    15,     5,   -17,    19,    -1,   -12,     7,    -8,    17,    -3,    12,    -7,    16,   -21,   -14,    -3,     6,   -16,   -27,   -36,   -49,   -12,    -8,    -8,    -8,    16,    12,    -7,   -20,     2,    14,    -5,    -3,   -12,    13,    14,   -16,   -26,   -42,   -49,   -77,   -69,   -64,   -84,   -53,   -37,    42,   -13,   -13,   -11,    40,    59,    27,    24,    80,   -23,   -14,    -1,   -12,     0,     2,   -35,    20,    -8,   -21,   -80,  -113,   -30,     4,    76,    20,    77,   113,   151,    52,   -40,   -81,   115,   -30,   -27,    34,   -43,   -54,   -60,    16,    31,    -8,    12,   -12,   -47,     3,   -60,   -64,    61,    -5,  -109,    88,     2,    67,    75,   -74,   -82,   -30,    25,   -46,    27,    89,   -70,    22,    78,    95,   174,   163,    50,   -44,    10,    16,   -35,    11,     1,    16,   -47,   -90,    12,   121,   117,     7,   -92,  -102,   -67,   -30,    52,     7,    37,    11,    30,    78,    82,    79,   122,   103,    97,   -37,    -8,   -22,   -22,   -25,    46,    29,   -72,   -28,   109,    20,    36,  -101,   -88,   -17,    39,   113,    46,    99,    72,   -29,    29,    59,   110,   -22,    62,    57,    99,     3,     1,    -3,    -3,   -67,    -7,   -15,   -49,    59,    67,    88,    73,    -8,  -101,   -47,   105,    94,   152,   115,    40,    30,    35,    27,   -35,   -71,   -51,    72,    72,    28,    -1,   -14,  -112,   -86,   -96,   -49,    -3,    29,   135,    97,    89,   -66,   -43,   -94,   -19,    28,   -37,    16,    32,   -61,   -24,  -102,   -57,   -58,   -53,   -72,   116,    21,   -11,   -27,  -110,  -105,   -57,   -30,     8,    17,    69,    74,    44,    70,  -140,  -176,  -207,  -249,  -274,  -356,  -196,  -263,  -255,  -240,  -158,  -118,  -113,   -72,   116,    60,    15,   -11,   -36,   -82,   -35,   -14,   -46,    10,    56,    54,    26,   -34,  -133,  -171,  -204,  -147,  -145,  -300,  -327,  -287,  -346,  -330,  -303,  -138,   -77,   -43,    36,    71,   -11,    -8,   -11,   -16,    -9,   -43,    -4,   -20,    43,    28,   -65,   -27,   -45,   -59,    -2,    43,    53,     4,   -83,   -94,  -168,  -188,  -222,  -181,  -139,   -33,     6,    21,    -2,    -8,     3,    59,     6,    57,    67,    25,    93,    14,    74,    12,   -38,   -49,   -50,    36,    40,    33,    38,   -37,    10,    19,   -84,   -51,   -90,   -71,    -5,     8,   -10,    12,     3,    29,    73,    32,   -52,   -47,   -21,    37,     4,    46,   -46,   -54,   -79,   -86,    -7,    -8,    21,    13,     5,     5,    17,    63,   -23,   -44,   -56,   -93,     5,   -33,   -27,     6,   102,    40,    88,     3,   -22,    61,    -1,   -32,   -33,   -87,   -66,    13,   -18,   -69,   -40,   -80,   -10,   -25,    57,    26,   160,   -78,  -105,   -56,     4,    35,   -23,  -130,   -83,  -114,    44,   -93,    -1,   -28,    63,    57,   -36,   -47,   -54,   -68,   -32,  -140,   -75,     4,    18,   -43,   -13,   -15,   135,    -1,   -83,   -89,   -20,   -19,   -13,   -71,  -141,  -111,   -65,   -33,   -53,    20,    46,     1,   -28,   -75,   -15,   -22,   -20,   -60,  -140,   -62,   -28,    19,    30,    18,    -5,   -75,  -152,  -136,   -10,   -30,   -57,    75,     2,   -73,    35,    16,   -57,   -24,    12,    10,    -6,   -51,   -97,  -131,   -63,   -76,   -33,    50,    30,    33,    40,    11,    10,   -13,  -147,  -141,   -12,     4,    62,   102,   -46,    29,   -27,    -4,   -15,   -94,     7,   -34,   -70,  -112,  -206,  -111,   -93,   -89,   -21,     6,     0,    79,   -64,   -71,   -16,    -7,  -160,  -135,    15,     3,   115,   103,    47,     6,   -53,  -110,  -172,   -94,   -53,  -126,   -59,  -209,  -107,  -141,  -117,    25,    33,    59,    89,    41,    13,   -56,   102,     4,   -30,   -97,    -8,   -11,    59,    77,    74,   -22,   -72,   -64,   -53,   -14,   -38,   -39,   -42,    22,   -36,    53,    19,    72,    49,    43,     0,    18,     3,   -23,   -48,   -18,  -107,    13,   -17,   -11,   -31,    38,    70,   -11,    18,     5,   -71,  -127,     4,   -35,   -24,    -4,   -71,    84,    34,   105,    22,   -29,     1,    51,    64,   100,    34,   107,   -18,     3,   -15,     9,   -75,    34,   -27,    32,     3,   -23,   -31,   -66,   -82,   -28,   -38,   -35,   -62,    74,    76,    19,    19,   -14,    15,     7,    25,   168,    36,   164,   153,    -4,     2,   -18,    57,    57,    -4,     9,   -18,   -45,    64,    14,   -37,    -8,   -25,    -7,    21,   -46,   -43,   -42,   -47,   -67,    82,    23,    84,    77,    47,   115,   187,   -19,   -10,   -11,     5,    76,   106,    52,    82,   -46,   -27,    63,   -28,   -74,   -10,    56,    35,    93,   -80,   -14,   -10,    17,    17,    41,   -33,  -112,   -23,   -43,   -21,     5,   -19,     7,    18,    97,   -86,   -50,   123,    66,   111,   130,    90,   -19,   126,    87,    93,    73,   -66,    -3,    70,   108,    98,    78,   150,    90,    65,   -18,    12,     2,   -17,   -18,   -10,   -10,   -18,   -30,   -27,   -18,     4,    10,    -1,    25,     9,   108,    58,    18,  -162,   -73,   -36,    19,   -95,   -61,    21,   -46,   -30,    13,    18,   -11,     8,    -9,     6,    10,    12,   -14,     0,     4,   -18,    17,     5,    -8,    -8,     7,   -39,   -29,   -16,    -3,    -6,   -34,   -78,   -99,   -84,     0,     4,    10,    -7,   -11),
		    96 => (  -10,    11,   -13,     7,   -15,    -5,   -14,   -16,    15,     7,   -12,   -19,    80,    84,   -19,    -1,    15,   -18,     0,    14,     7,     2,     8,     8,     6,    15,    11,   -13,     3,    18,    -3,     7,    13,    40,    39,    78,   118,    75,    60,    39,   114,   175,   -55,    35,    77,   106,   100,    28,    87,    44,    44,    28,    12,     7,    11,   -15,    -4,     9,     7,    -7,   113,   125,    85,    87,    47,    54,    93,   130,   203,   143,    74,    70,    88,    99,    33,     6,    25,   -26,   -23,   -27,    33,    24,    15,     4,   -10,    11,   -15,   160,     3,    19,   139,   168,    90,    61,    98,    17,    45,   153,   101,    60,   -27,   -90,   -64,   -11,    40,   -64,   -29,   -28,   -14,   -25,     1,    15,    -9,     2,   -30,   189,    12,   144,   111,    -2,   -10,    26,    27,    25,    78,    16,    -4,   -51,   -77,   -20,   -35,   -52,  -161,   -88,  -120,  -123,  -119,   -90,   -11,    28,     1,     4,   -26,   -36,    57,    44,    -8,   -49,   -68,    19,    35,     5,    94,    11,  -127,    -8,  -136,   -43,   -49,  -104,  -176,  -181,  -210,  -144,   -82,   -55,    35,    33,    13,   -20,   -17,   -98,    45,   -28,   -60,  -127,  -111,   100,    43,    73,    57,    10,   -45,  -141,  -101,  -115,  -235,  -236,  -159,  -237,  -216,  -202,  -101,   -30,    15,   -71,    -9,    -1,   -13,  -120,    55,    26,  -101,  -137,    -7,    -8,    54,    49,    23,     5,   -81,  -155,  -217,  -223,  -279,  -189,  -132,   -36,  -224,  -223,  -163,   -64,    33,   -90,   -12,     6,     9,  -106,    76,     2,   -47,   -40,    68,    47,    13,    -5,   -36,     0,  -196,  -323,  -233,  -132,  -140,     3,    11,    47,   -67,  -118,  -157,  -141,    11,  -101,     1,   -23,     1,   -31,    84,   -19,   -80,   -24,    49,   -16,   -21,    28,    -1,  -214,  -139,  -106,   -34,   -10,   -15,   111,   128,   105,    60,    32,    -6,  -120,   -91,   -46,    -9,   -27,    -8,   -36,    39,    35,   -53,    -5,    51,   -55,    24,   -24,   -31,  -239,  -150,     8,    31,   106,    89,    48,    58,    40,   -20,   -14,    37,   -48,  -124,  -145,    11,    20,   -21,   -64,    72,    61,   -80,    27,    15,   -38,   -45,   -59,  -100,  -208,  -107,    -2,    65,    53,    52,    55,    67,    -4,    -2,   -24,    17,    10,   -58,   -74,    -8,     1,   -39,  -111,    24,   -13,   -24,    -1,    27,   -25,   -46,   -45,  -111,   -59,    67,   -62,    75,   -32,    53,    71,    73,    38,    80,    80,    92,    44,   -92,   -87,    -7,    -4,   -38,  -107,   -34,    68,    35,   -49,    -2,   -24,    22,  -103,  -146,   -41,   -11,    -4,    51,    -5,   -93,    57,     8,    54,    58,   126,    99,    32,   -76,    17,     9,    -5,   -26,   -92,   -65,    30,    94,   -34,    70,   -20,    32,    13,   -72,    -3,    12,    49,    18,     4,    83,   -61,    38,    24,    84,   107,    22,   180,   -21,     3,   -14,     6,   -36,   -63,   -80,   -26,    80,   -13,     7,    15,     0,   -10,   -23,    62,    59,    21,   -24,   -32,    21,   -52,    34,    55,   -19,   -14,    37,   129,    -2,  -116,     6,    -5,   -43,   -89,   -40,    15,    65,    12,   -32,     8,    52,    89,   -51,   -15,    51,    -2,    21,    -9,  -102,    28,   -46,   -14,   -53,    20,    87,   125,    -2,   -70,   -15,     7,    15,   -81,   -53,   -43,    -3,   -19,    57,   -54,     0,   -51,   -31,    25,    78,    55,   -36,   -72,   -62,     1,  -109,   -23,   -45,     6,   136,   121,   -13,   -66,    19,    16,    -7,   -82,    49,   -47,  -105,    47,    -2,   -52,  -148,   -88,   -62,    -3,    38,   -25,   -24,    11,   -19,   -30,   -18,   -37,    19,    74,    74,    20,   -46,   -39,     4,   -20,    -5,   -32,    81,   -70,   -54,    25,    38,     3,    -3,  -104,  -100,   -49,    87,    73,    62,   -31,  -108,   -44,     2,   -27,   -33,    -3,     4,    66,   -53,     7,     9,   -19,     5,   -54,    79,     2,  -112,   -30,   -95,   -26,    18,   -71,  -103,   -45,    44,   165,    85,    35,    82,   -51,    58,   -46,   -77,   -87,   -46,    53,    12,    -2,    11,   -10,   -15,   -34,    22,   -15,    -8,    37,   -72,   -36,   -46,   -77,   -97,    25,    64,    53,    21,    47,   -61,  -105,    18,   -70,   -39,   -85,   -99,   -13,    24,    11,    17,     4,   -22,   -30,   -34,    -5,    35,  -104,  -180,  -118,   -86,  -148,   -77,    14,   -13,   -60,   -86,   -41,   -73,  -108,   -57,  -152,  -165,  -173,  -180,   -44,    36,     2,     0,   -15,     3,   -24,   -45,   -13,   -20,   -55,   -77,  -149,  -205,  -156,  -117,   -26,   -26,  -137,  -254,  -266,  -224,  -136,   -35,  -124,  -135,   -87,  -153,    -5,   -12,   -13,    13,   -14,    -9,    -2,   -19,    -3,     2,   -30,   -30,    -8,    -7,    34,     6,   -69,  -115,  -113,  -160,   -80,  -130,  -158,   -47,   -37,   -41,     0,   -12,   -15,    -3,     2,    15,    17,   -20,    -7,    10,     2,   -25,   -39,   -36,   -27,   -21,     3,   -14,     2,    -9,   -20,     2,   -10,   -17,   -45,  -112,   -48,   -75,   -62,   -19,    18,    -8,    11,     9,    20,     1,   -12,   -12,     1,    14,   -25,   -20,   -18,   -21,   -54,   -25,   -10,   -42,   -28,   -19,   -20,   -24,     7,   -31,    -7,     9,    -8,     8,     3,    -4,   -14,     4,     2,     8,   -15,   -20,     5,    16,     1,    20,   -14,   -41,   -10,    16,     9,    -7,     4,    -3,    -3,     7,   -15,   -10,     8,     9,    12,   -18,   -15,     0,   -20),
		    97 => (   -3,     8,    18,   -18,    19,    -8,    20,     8,   -14,    -6,     1,    -2,    -2,     8,   -19,    -5,    12,    20,     5,    15,     6,    -6,   -19,    11,   -14,     5,    -2,    -5,     7,    11,     5,    17,   -14,   -15,   -20,    15,   -14,    -3,   -13,   -74,   -41,   -45,    14,   -37,   -91,  -130,    -4,   -29,    -4,   -11,    -5,     3,   -17,    -2,   -11,    -9,    20,    -6,   -16,   -20,   -39,    -8,   -15,   -33,   -20,   -74,   -80,  -156,   -24,   -12,   -31,   -63,   -38,     0,    -8,    -1,   -37,   -31,   -51,   -56,    -5,    -6,     2,     1,    -2,   -10,    15,   -34,   -11,  -100,   -91,  -204,  -179,  -153,  -179,  -219,  -193,  -219,  -114,   -50,   -45,   -41,     0,   -64,   -87,   -92,  -152,   -40,   -30,   -42,   -11,     6,     6,    -5,   -23,   -30,  -111,  -147,  -158,  -171,  -264,  -276,  -256,  -141,  -143,  -139,  -131,   -90,  -189,  -144,  -102,   -91,  -106,   -58,  -117,  -215,  -217,  -120,   -41,    17,     4,     3,    13,  -134,  -226,    43,  -105,   -35,    27,    44,   -72,   -49,     9,    64,    88,   -15,    84,    30,     4,  -101,  -180,  -113,   -73,  -243,  -167,  -208,  -100,    -5,    -3,    -2,    79,    80,    67,   -60,   -50,   -46,   -61,     6,   -22,     5,    38,    11,    36,    75,   -20,   -47,   -22,    23,   101,    70,    73,   -91,  -166,  -128,  -122,   -75,   -17,    94,    99,    37,    77,   -87,   -42,    20,   -25,    -3,   -34,    27,    45,    23,    36,   -46,   -44,   147,     8,   -35,     9,    -9,   -21,   -35,    -6,  -135,  -174,   -89,   -92,   201,    47,   -15,    46,    -2,   -60,    29,    42,    82,    73,    43,     7,   -33,   -53,    -3,   -26,    54,    93,    26,    61,     2,   -51,   -57,   -68,  -201,  -234,   -71,    20,   100,   -32,    20,    62,    47,    57,    17,    63,   123,   115,    20,   -92,   -43,    44,    40,     7,    61,    72,    -4,    78,    -3,    43,   -51,   -92,   -17,    -9,   205,    10,    81,    55,     0,    59,    55,   -14,    67,   110,    57,    60,   -75,  -131,   -34,    60,   133,    62,    -2,    49,    31,    92,    -1,   -28,   -77,   -75,    52,     4,   176,   -14,    15,   132,    33,   -38,   -12,   -14,    37,    65,    46,   -65,   -66,    51,   101,   178,   118,    81,     2,    65,   -43,    36,   -54,     3,    46,    29,  -147,   -83,   111,     1,    57,   126,    32,   -62,   -57,   -12,   -12,    48,    13,    34,   100,    83,    89,   176,   160,   101,    55,     9,   -93,   -29,    -3,   131,     5,    43,    91,    71,   102,     3,    30,   123,     0,  -101,   -60,    30,   -14,     5,    33,     6,    68,    87,    62,   203,   129,    86,    35,   -83,   -75,  -139,   -47,    20,   -41,     8,    91,   -28,   -78,   -23,    48,    52,   -83,  -128,   -14,   -25,   -71,    -9,    16,   -44,    29,    13,    28,   117,    25,    32,    52,   -41,   -42,   -63,  -120,   -38,    23,    80,   -84,  -102,    -3,   -11,    -2,    26,   -79,  -100,   -21,    11,   -35,  -140,  -124,   -52,   -32,   -51,    10,   -33,   -59,    -2,    47,   118,   -26,    18,    15,   109,    75,    71,    30,   -44,   -60,     5,   -28,    -8,   -64,   -31,    -9,     2,   -19,    -1,    78,    57,   -51,  -126,   -72,   -66,   -25,   -38,   139,   214,   166,    45,   136,    84,   126,    97,   -89,   -83,   -72,     7,   -29,   -24,   -42,    -2,    17,     3,   -68,    -5,    -3,    -1,   -90,  -150,   -53,     3,     4,    99,   146,   184,    34,    98,    63,   123,   103,    13,    62,   -23,  -108,    26,    10,    39,   -38,   -10,    72,    69,   -39,   -67,   -88,   -38,   -75,   -83,   -55,   -36,    13,    29,   208,   116,    62,    34,    19,    70,    27,     7,    22,     8,   -72,   -18,    39,    10,   -13,    29,    42,    42,    20,    45,   -81,   -43,   -44,   -78,  -107,   -49,   -55,   114,   215,    76,    69,    11,    36,    12,    -9,    62,   -20,   -80,   -24,     8,    50,   -20,   -51,  -132,    25,     7,    48,    41,    12,   -30,   -34,   -51,     2,     1,    38,     7,    45,   -13,    -8,    -9,   -10,   -52,   -47,    51,   -52,   -91,    10,    -2,    10,   -15,   -43,   -86,    74,    64,    72,    45,    86,    79,    12,    25,    22,   -38,    44,    13,   -67,  -102,   -78,   -44,    31,   -39,   -29,   -87,   -71,   -25,    14,    -7,    -7,   -51,   -88,   -94,    44,   125,    58,    11,    12,    41,   -22,    40,    29,   -25,   -86,    -9,  -109,   -84,   -94,  -104,   -77,  -146,  -141,   -90,    13,   -93,   -15,   -15,    18,   -38,  -158,   -81,    63,   116,    75,    42,    -7,    87,    -6,   -34,    -5,  -156,  -129,   -56,  -119,  -144,  -118,   -82,   -81,  -166,  -151,   -54,    13,   -73,    12,    -1,    10,    -1,   -24,    -9,    84,    39,    73,    -3,     6,    -1,    23,   -12,     3,   -91,  -109,   -72,   -59,  -166,  -151,  -128,   -35,  -140,  -157,   -89,   -78,   -12,    17,   -11,   -16,   -51,    97,    -8,    -4,    10,    25,   -68,    39,    35,   -19,   -29,    20,  -143,  -125,     6,   -92,  -122,  -168,  -106,   -27,    -7,  -107,   -42,   -21,   -12,    -5,   -17,    -8,   -11,  -105,   -71,  -102,   -56,   -51,    16,   112,   -17,   -33,    -9,    -9,     7,    20,   -26,   -99,   -26,   -25,     0,    45,    -8,    -3,   -16,    -2,    16,    10,    -2,    19,   -17,     3,    44,    55,     1,   -51,   -36,     1,    -2,   -81,   -25,   -47,   -86,    25,     8,   113,    45,   -47,     1,    58,    -7,    77,   -13,    -1,    -8,   -16),
		    98 => (   12,   -13,   -12,    -5,    11,    -8,     4,    20,     4,    -6,     7,   -11,    11,   -15,     2,   -19,   -18,    -8,     8,    11,     4,   -16,    -8,    -9,    -2,     5,     0,     2,     4,    16,     9,    20,   -15,     3,    19,    14,     9,    10,     1,    12,   -16,   -30,   -28,   -72,   -68,   -73,   -28,    19,   -24,   -17,     0,   -19,   -10,   -13,   -11,    10,     8,    20,   -19,    -4,    -1,    -4,    10,    -7,   -41,  -113,  -155,  -145,   -54,    -9,   -33,   -99,   -99,   -38,   -16,     3,   -23,   -35,   -56,   -38,    -1,    -2,     1,     3,    16,    20,   -23,   -12,   -24,   -59,   -46,  -193,    64,    92,   121,    49,   117,   135,    87,    47,    12,    43,   -36,   -89,   -72,  -116,   -69,    -7,   -25,   -31,   -21,   -10,     6,   -26,    18,   -21,  -122,  -141,   -28,    30,    41,    54,   -38,   -89,    12,   -35,   -21,   -34,   -14,     7,   -15,    38,     6,    31,  -125,   -68,   -28,    -4,     9,   -28,    -4,   -12,    -2,  -101,  -123,  -218,   -65,    39,    53,   -51,    -6,    19,  -112,   -63,    51,   -12,    25,    75,    44,     2,    59,    -5,   -50,   -78,   -64,   -24,    26,   -21,    16,    -8,  -116,   -57,   -49,   -65,     6,   167,    86,    52,    55,    25,     7,    28,    40,    69,    50,     3,   -64,    55,   -46,   -15,   -64,   -22,   -59,   -54,     5,    -7,   -18,   -74,   -43,   -96,   -31,    -8,    95,   138,   -81,   -32,    30,   -66,   -18,   -68,   -49,   -47,   -69,   -16,     2,    35,   -23,   -90,   -50,   -77,   -34,   -40,   -25,   -26,   -23,   -44,   -80,   -51,  -124,  -116,    37,   145,   -52,   -36,    77,    45,   -46,   -96,  -101,   -45,  -151,    18,     1,    20,   -29,   -39,   -19,  -100,     3,    41,    49,    -6,    13,   -10,   -32,   -25,  -152,  -114,   -20,   -43,   -50,    12,    92,   109,    47,   -55,   -71,   -39,   -16,    73,   -86,   -17,     2,    46,   -21,   -46,   -26,    22,  -128,  -120,    12,   -31,   -58,   -65,   -72,  -147,    41,   -66,  -188,   -42,    58,   202,   186,   125,    45,   -14,    12,    27,    28,  -100,    87,    48,    12,   -78,  -137,  -161,  -133,  -132,    -4,   -20,   -19,   -87,   -55,   -57,     7,   -15,   -70,   -14,  -144,     9,    98,   154,   110,    -1,   -36,   -83,   -29,   -34,   -23,   -25,   -65,   -64,  -150,  -109,   -34,   -48,     5,     9,   -36,   -19,   -33,   -75,   -40,  -107,  -159,  -163,  -193,  -190,    13,    12,    39,   123,    27,    -9,    39,    45,    12,    32,    28,   -13,   -21,   -84,   -60,   -43,   -14,    -6,   -41,   -13,   -51,   -29,   -17,   -91,  -156,  -222,  -171,  -127,   -98,    -7,    -5,    78,    31,   -31,   -14,   -52,  -106,     6,    31,  -112,  -103,   -79,   -71,   -21,   -11,   -14,     4,   -98,   -56,    18,    -5,   -60,   -80,  -115,   -20,    53,    24,    22,   -19,   -64,     1,    11,     4,   -87,   -45,    51,   -33,  -111,  -112,   -64,  -129,   -64,   -20,    16,   -60,   -71,   -90,   -45,   -59,     3,   -29,    20,    -1,    44,   -25,   -79,   -51,   -23,    60,   -41,   -81,     6,    -5,    47,   -98,   -71,   -78,   -67,  -143,   -53,    -3,   -21,   -38,   -37,   -71,    -9,    74,    57,    18,    98,    19,     4,   -79,   -20,  -125,     4,  -125,    84,   -64,    75,    74,    38,   -46,   -22,   -45,   -37,  -176,   -69,    15,    -8,   -54,  -137,    41,    18,   -40,    72,    64,    13,   -47,   -14,   -34,  -149,  -130,   -35,   -95,   -30,    30,    95,    25,   110,    88,    -2,   -73,   -59,   -34,   -82,   -21,   -11,   -27,   -46,   125,     0,    37,    88,   -20,   -78,   -52,    30,   -55,  -136,   -55,   -46,  -172,   -60,    36,    61,    56,    53,    46,    32,  -118,   -63,    -4,   -52,    -2,   -39,   -78,    84,    91,   122,    91,    42,   -93,   -51,    11,    31,  -131,   -82,   -91,   -25,   -55,    -9,   -50,     1,    34,    53,     8,   -72,  -106,   -43,  -151,   -51,   -17,    -8,   -65,    14,    81,    43,    61,    41,   -36,  -115,   -22,    21,   -94,   -22,   -17,    25,    55,   -52,   -56,   -41,    63,    52,    27,   -64,   -55,   -11,  -132,   -18,   -51,   -29,   -75,   -75,    18,    -7,     7,   -14,   -59,     4,   -48,    -9,    20,   -51,    58,   -36,   -41,   -78,  -123,    25,    58,    70,   -22,   -52,   -75,   -45,  -111,   -21,   -54,   -38,   -67,   -89,   -76,    10,   113,    82,   -69,   -43,    18,    33,    56,   -79,   -18,  -101,   -65,   -31,   -59,   -31,    15,   -40,  -117,   -42,     8,   -12,   -70,    -7,   -18,    17,   -19,   -35,  -111,    71,    22,    89,    23,   -76,   -40,   -73,    15,   -12,    -4,   -31,   -40,   -84,   -34,    -6,   -54,  -154,   -68,   -29,     6,    57,  -105,   -11,   -19,   -14,   -42,   -29,   -87,   -90,    43,    36,    24,    -4,   -71,   -61,   -12,     3,    48,    61,    95,   -58,    10,    -9,    -4,   -58,   -58,   -15,   -85,   -13,   -27,    -6,     6,    13,   -10,    -8,   -20,   -59,    -2,   -35,   -88,   -58,   -95,  -107,   -91,  -111,  -110,  -121,   -89,   -54,   -24,    -6,    -1,   -47,   -20,   -22,   -22,    -7,   -20,    16,    -6,   -19,   -14,   -42,   -33,   -21,   -12,   -26,   -27,   -28,   -38,   -21,   -79,   -94,  -116,   -64,   -52,   -39,   -37,   -78,  -130,  -126,   -70,     9,    -2,   -15,    19,    -3,   -16,    -7,    16,     1,   -30,   -23,   -41,   -22,   -26,   -29,   -13,   -15,     1,   -71,   -24,   -16,   -30,   -31,   -33,   -22,     6,   -14,    17,   -12,    -9,   -12,   -16,     5),
		    99 => (    4,    10,    -4,    -3,   -20,   -16,   -15,   -16,   -17,   -16,    -3,    -7,     4,   -12,     8,     6,    -2,   -14,    16,     8,     0,    19,    -6,   -20,   -14,     7,     5,   -12,   -15,     0,   -20,     6,     7,    18,    12,     5,   -10,    -7,   -30,   -41,   -57,   -57,    13,   -15,     7,   -11,   -29,    -1,     0,    -7,   -29,   -13,    -5,    -3,     8,    -8,    -2,    13,   -11,   -15,   -13,     6,    -9,   -15,    -4,   -23,    -1,   -31,    -2,    11,   -43,     6,     7,     6,   -16,     3,   -28,   -33,   -40,    -6,     4,     5,   -18,    -5,    12,    -2,     3,   -44,   -20,   -33,   -30,   -21,   -69,   -55,   -32,    -5,    14,   -23,   -24,     6,   -11,   -27,   -31,   -35,   -69,   -17,   -58,   -34,   -67,   -45,    -8,   -18,    -1,     3,    -8,   -19,   -26,   -28,  -105,    -8,     8,     4,     4,   -29,   -85,   -79,   -39,   -89,   -50,   -88,   -43,  -108,  -152,   -16,   -15,    -9,     6,   -95,   -31,   -10,    18,    14,   -15,   -41,   -14,     8,    -5,   -27,   -27,   -43,   -24,   -63,   -84,  -110,  -130,  -151,   -93,   -27,   -15,    42,   -58,   -49,   -51,   -26,   -13,   -29,   -43,    14,   -13,    14,    -7,   -45,   -11,   -44,   -62,   -56,   -96,   -29,   -57,    -4,   -15,   -10,    -5,     2,   -56,  -104,   -37,   -63,   -82,   -61,   -58,   -36,   -25,    -3,   -37,   -52,     9,   -13,   -22,   -39,   -37,   -63,  -117,  -147,  -149,   -75,   -58,    19,    -1,    47,    10,    28,    49,   -76,   -29,   -78,   -70,  -124,   -65,    43,   -46,   -14,   -17,   -36,   -71,   -60,   -27,   -40,   -80,  -101,  -117,  -161,  -105,   -82,     4,    22,    23,   -30,    14,     2,    74,   -72,   -27,    24,   -15,    -2,   -74,    -1,   -11,   -88,   -21,    -1,     0,   -73,   -56,   -71,   -93,   -58,  -107,   -31,    17,   -35,     6,    34,    45,    28,    31,   122,    31,   -39,    16,    80,    17,    -1,    -1,   -16,   -40,   -63,   -42,   -37,   -18,   -87,   -59,     2,   -46,   -69,   -98,   -45,    19,   -67,   -97,    45,    47,    27,    81,    11,    55,   -41,    79,    58,   -20,     9,   -18,   -74,   -69,   -68,   -28,   -53,    -3,  -160,   103,     2,   -29,   -41,   -49,    -6,    -1,   -44,  -121,     4,    24,    66,    39,   -10,   -58,   -82,    -5,    14,    13,   -26,     1,   -39,  -103,   -95,   -19,   -31,    -5,   -74,    35,    89,    75,     7,    42,     0,   -52,  -158,  -103,   -18,   -33,   -49,     7,    -5,   -27,    -5,   -20,    41,     1,    56,   -12,   -20,  -101,   -51,   -74,    -9,    14,   -79,   -29,    51,    46,    25,    49,   -13,   -57,  -189,   -52,   -25,  -132,  -123,   -74,    14,    -5,   -73,    14,    11,   -41,    71,    21,   -43,  -120,   -73,   -38,     6,    -6,   -54,   -68,    65,    56,    55,    -8,   -16,  -129,  -113,   -36,   -25,   -85,   -91,  -105,   -24,   -28,   -63,    -3,    18,    42,    48,   -33,   -88,  -100,   -56,     3,    -4,   -13,     9,   -98,    61,    91,    25,    30,     2,   -74,  -134,   -28,   -63,   -83,   -16,   -11,     7,     1,  -110,    14,   -14,   -22,    35,    37,   -98,  -115,   -62,     3,   -35,     7,   -29,   -60,    61,   116,    74,   134,    45,    17,    27,    20,   -80,    13,     3,    13,    -1,  -119,   -79,   -57,   -80,     3,   -17,    79,    53,   -97,   -11,   -53,   -18,     6,   -22,  -155,   -10,   -14,    -4,    48,    76,   113,    85,    68,    94,    59,   -13,   -25,   -72,   -92,  -105,   -14,   -56,   -41,   -17,    69,   -23,   -96,   -35,   -68,   -64,   -16,     2,  -151,    44,   -43,   -75,   -16,    35,    -9,   -15,    95,    20,    -9,  -116,   -32,     0,   -37,   -32,    -8,  -101,   -18,   -42,    59,    54,   -46,   -14,   -84,   -44,   -17,   -23,   -85,    66,     2,   -87,   -76,   -51,  -111,   -96,   -37,   -36,     9,  -124,    37,     1,   -56,   -56,   -40,  -128,     3,   -77,   -22,    75,    87,    58,   -71,   -11,   -19,     0,   -31,    64,    49,   -18,   -58,   -77,  -114,   -68,   -92,   -50,  -144,  -102,    44,    38,   -59,  -109,   -40,   -59,    20,    -3,   -24,    77,    89,   160,   -81,   -14,     3,    15,   -55,    24,    28,   -14,   -49,   -52,   -63,  -106,   -70,   -25,   -21,   -66,    61,   -46,  -201,   -55,   -20,   -40,   -29,    60,   -63,     4,    38,    97,  -100,   -11,    -8,    14,   -64,   -48,   -86,   -31,   -44,   -71,   -42,   -63,   -37,   -65,   -14,   -13,    98,  -115,  -133,   -18,    -2,   -35,     2,     9,   -16,    15,   -35,   -93,   -23,    -9,     3,    -6,   -53,   -48,   -46,   -15,   -24,   -34,   -35,   -14,   -48,   -12,    -1,     5,    34,   -54,    15,    37,    -9,   -41,    78,    -4,    98,    39,    -2,   -40,   -25,   -10,     7,   -15,   -42,   -10,   -70,   -38,     4,    29,   -75,   -82,   -46,   -24,     8,   -21,    27,    33,    61,   -37,   -12,   -10,    69,    43,    59,    39,     7,   -20,   -20,    10,    -1,   -17,   107,   -77,     0,    55,    22,    -1,   -99,   -39,   -34,    -4,   -34,   -72,    61,    49,    28,   -18,   -34,    39,    81,    53,    62,    10,   -30,   -24,   -12,   -17,     1,     7,    16,   118,    61,    50,    53,    -8,    11,    69,   -58,   -20,   -29,   -87,     5,    29,   -10,   -15,   -10,    52,    83,   129,    68,     3,    30,    12,    19,    -7,    -4,    -9,   -17,    -1,   -42,   -23,    37,    84,    68,    60,     1,    17,   -23,   -66,   -11,   -22,   -20,   -14,   -53,   -34,   -28,   -15,    38,   -45,    20,   -16,    -2,     0)
        );

 ---------------------------------INFO-
 -- COEF =172.55234

 -- MIN =-511.99997
 -- MAX =339.14417

 -- SUMMIN =-36377.68
 -- SUMMAX =26448.615
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
