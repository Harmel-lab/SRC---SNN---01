----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (   -1,     0,     0,    -1,    -1,     2,     0,     0,     1,    -2,     0,     2,     0,    -4,    -4,     1,    -2,     2,     1,     1,    -2,    -2,    -1,     1,     2,     2,    -1,    -2,    -2,    -2,     0,     1,     0,    -2,     2,     1,     0,     0,    -1,     2,     3,     2,    -3,     2,     7,     3,    -1,    -2,    -2,     2,    -1,     1,     1,     0,     1,    -2,     2,     2,     0,     2,     7,     0,    -3,     0,    -4,   -11,    -1,    -2,    -1,    -6,    -6,    -9,    -1,    -2,    -4,    -1,    -1,    -2,    -6,    -4,    -4,    -5,     1,    -1,     1,    -2,    -1,     5,    -1,     4,     3,    -8,    -5,    -4,    -7,    -5,   -10,    -6,    -9,   -10,    -3,     6,     0,    -8,    -6,    -4,    -6,    -3,     2,     2,    -1,     1,    -2,     1,     1,    -1,    -4,    -9,     2,    -6,   -13,    -6,    -6,   -10,   -17,    -1,     0,    -5,    -2,    -9,    -6,    -6,    -1,    -3,    -5,    -3,     1,    -3,    -5,     1,     1,     2,    -5,    -1,     0,    -3,    -2,    -1,    -4,    -2,    -8,   -15,    -9,   -13,     2,     6,    -1,    -6,     1,    -9,   -11,     0,    -2,    -2,    -3,   -11,    -3,    -3,    -2,     2,    -5,    -3,    -3,     0,    -3,    -2,    -5,    -5,    -4,   -16,   -11,    -5,    -1,    -5,     7,     5,     1,   -10,    -9,    -5,     1,   -11,    -5,   -10,    -3,     6,     0,    -5,    -4,    -4,     1,    -2,    -3,     2,    -4,    -4,   -10,   -16,   -16,    -6,    -1,     0,    11,     6,   -10,     0,    -9,    -8,     3,    -6,    -9,    -4,   -10,     6,     8,   -13,     7,     5,    -2,    -2,    -3,     0,    -2,    -9,    -6,   -16,    -3,    -3,     4,    -6,     2,    12,    -5,     2,   -10,   -13,    -3,    -7,    -4,   -13,    -4,    -3,    -3,    -2,    12,    -1,    -1,    -1,    -8,    -1,    -6,   -15,    -6,    -2,    -3,     4,    -3,    -4,     8,     2,     0,    -8,   -19,    -2,    -1,    -4,    -6,   -10,     0,     2,    -3,    -2,     3,     5,    -5,    -6,    -3,     4,     0,    -1,    -5,    -3,    -2,    -1,   -12,   -13,    -4,    -9,     3,    -8,    -9,    -3,    -8,    -9,    -4,    -3,    -9,     1,     1,    11,    -5,     2,    -6,    -1,    -2,    -1,    -4,    -3,    -8,     1,     5,    -4,    -5,     1,    -6,     2,    15,   -11,    -9,     1,    -8,   -12,    -4,    -7,    -5,    -2,    -1,     3,     2,     0,    -1,     2,     1,     0,   -12,     0,     2,    -3,     6,    -2,    -5,   -13,     1,     7,    13,    -2,     0,     8,     0,   -13,    -8,    -8,    -7,     2,    -1,     6,     6,    -2,     0,     1,     6,    -7,    -7,     1,    -3,    -9,     3,    -9,   -23,   -18,    -1,     6,    11,     3,    -2,     9,    -4,    -7,    -6,    -3,   -10,     0,    -1,     0,     0,    -3,    -2,     4,    -6,    -8,    -6,    -2,     3,     4,    10,    -1,   -16,   -17,    -1,     2,     5,     4,    -9,     1,    -1,    -5,    -6,     2,    -8,    -1,     0,    -2,    -5,    -4,     2,    -8,     0,   -13,    -6,   -10,    -2,     4,    14,     3,   -21,    -7,    -2,     3,    -1,    -3,    -9,     7,    -7,    -5,     1,    -5,    -6,    -1,    -2,     0,    -2,    -6,     2,     1,   -15,    -4,    -9,   -11,    -6,     6,     6,    -7,   -25,    -1,    -2,    17,    -5,    -3,    -7,    -6,     0,    -6,    -7,    -5,   -14,     6,     0,     1,    -8,    -4,   -11,    -3,    -7,    -7,    -8,   -20,     2,     3,     8,    -6,   -18,    -7,     0,     8,     3,     0,     5,    -6,    -3,     3,    -6,    -8,   -14,     5,     0,     1,    -4,     3,    -4,    -6,    -3,    -1,    -6,   -10,     7,     7,    -6,   -10,   -21,    -2,    -1,     1,    -3,     0,     0,    -2,     2,    -5,     0,    -1,    -6,    -3,     2,     4,     1,     3,     1,    -6,    -3,   -10,    -7,     2,     6,     6,     0,   -11,   -12,     8,     2,    -7,    -5,     0,   -10,    -4,    -4,    -4,     1,   -18,    -4,    -2,    -1,     0,    -2,    -4,     2,    -2,    -6,   -13,   -10,     3,     1,    -7,    -8,    -2,    -3,     2,     3,    -6,     0,   -11,    -7,    -8,    -2,    -2,    -3,    -4,     2,     3,     1,    -1,    -6,    -6,    -3,    -3,     0,    -8,    -5,    -3,     2,    -3,     0,    -2,    -2,     5,    -2,    -2,    -7,   -10,   -10,    -5,     2,     1,    -9,     1,     4,     3,     0,     1,    -5,   -15,     1,     1,     3,     1,    -5,     3,     1,     5,    -2,   -11,     8,     7,     7,   -15,    -6,    -8,    -7,    -5,     2,    -2,    -1,    -2,     4,     1,     1,     1,    -5,   -11,    -5,     2,    -4,    -1,    -5,   -11,     6,     3,     5,     7,    -8,    -7,    -8,   -18,     0,   -11,    -7,    -3,     5,    -1,    -4,   -10,    -5,    -2,     2,    -2,    -3,     0,    -6,     6,     3,     2,   -11,   -13,    -8,    -8,     2,    13,     3,     2,   -11,    -4,    -2,    -8,    -7,     4,    -5,    -6,     0,    -2,    -2,     1,     0,     2,     1,    -2,   -18,    -7,    -7,    -6,    -3,    -6,   -11,   -12,   -18,   -17,   -21,    -9,    -5,    -6,    -7,    -5,    -9,    -3,    -6,    -5,     0,     0,    -1,     0,     0,     2,    -2,    -1,    -2,    -8,   -13,     1,    -1,    -8,    -5,    -2,    -7,    -5,    -6,    -6,    -3,    -9,   -14,    -6,   -10,    -6,    -3,     0,    -2,    -1,    -2,     0,     1,    -2,     0,    -2,     0,     1,     1,    -1,    -1,    -2,     1,    -1,     1,    -6,     1,     0,    -4,     0,     2,     0,    -1,    -3,    -3,    -5,    -1,     0,    -3,     2),
		     1 => (    0,    -1,    -1,     2,     0,    -1,     0,    -1,     2,    -2,     1,    -2,    -1,    -2,     1,     2,     0,     1,    -2,     1,    -2,    -1,     2,    -1,     0,     1,    -2,     2,     2,     2,     2,     2,    -2,     2,     1,     1,    -2,    -1,    -1,    -2,    -4,    -3,     8,     6,     0,    -4,    -3,     2,    -2,    -2,     0,    -1,    -2,     2,    -1,     2,     1,     0,     0,     2,     1,    -1,     2,     1,    -7,    -7,     0,    -2,    -2,    -2,    -4,    -8,   -10,   -11,   -14,     1,     5,   -12,    -4,    -1,    -2,    -3,     1,     2,     2,    -2,    15,    11,    -1,     2,     2,    12,    10,     6,     7,     4,     1,   -19,   -19,   -19,   -17,    -5,    -5,    -2,     2,   -10,     5,     1,    -7,    -1,     2,     2,     0,     0,    10,     9,     5,    -3,    -2,     0,     0,    -2,    -7,   -18,   -17,   -21,     2,     8,     1,     2,     3,     4,     2,     4,    -5,   -21,   -11,   -17,   -10,   -10,     1,    -2,    10,    14,     4,     1,    -5,    -5,   -24,   -11,    -9,   -15,   -20,   -11,    -1,    14,    -1,    -1,     0,     5,     6,    -6,    -9,   -20,   -15,   -11,   -10,    -9,    -1,    -1,     0,     6,     5,    -4,     0,     2,   -20,     1,     2,   -15,   -15,    -8,   -11,    -4,    -1,     5,    -1,     6,    -6,    -7,    -3,   -21,   -15,    -6,    -1,    -3,    -2,    -1,    -4,     4,     3,     0,    -4,    -8,   -22,    -5,   -11,   -18,   -13,    -2,     8,     4,     4,    -1,    10,    -2,    -8,    -5,     0,   -13,   -14,    -6,    -6,    -4,     0,    -3,    -3,    -3,    -2,    -3,    -7,    -8,   -15,   -13,    -6,   -24,   -23,     0,     6,     5,     9,     5,     3,    -5,    -8,    -4,    -7,   -12,   -15,    -8,    -8,    -2,     2,     0,    -3,     4,    -3,     0,   -11,    -6,    -4,    -7,   -17,   -32,    -8,    -2,    -4,     0,    10,     2,   -10,    -7,   -14,    -6,    -4,    -8,   -13,    -7,     0,    -8,     0,     3,    -1,    -3,    -1,    -1,   -10,   -13,    -9,   -11,    -2,   -16,   -13,    -6,     2,    12,    10,    -2,   -10,    -9,   -13,    -5,    -5,    -6,   -14,   -16,    -1,    16,     1,     0,     2,     4,     5,     1,    -6,    -8,   -13,   -21,   -11,   -18,    -5,    -7,     0,    15,     1,   -13,    -8,    -4,    -5,     2,    -4,    -8,   -15,   -14,    -1,    14,     0,     1,    -5,    11,     3,    -3,    -4,    -3,   -20,   -17,   -10,   -10,     1,    -4,    10,    -2,     6,   -20,   -22,    -7,    10,    13,    13,     9,    -4,     0,    -2,     9,     1,    -2,    -1,     3,     5,    -4,    -5,    -2,   -10,   -23,   -10,    -5,    -4,     3,    12,    -5,     4,   -19,   -22,     2,     9,     1,    -1,   -17,    -9,     1,     5,     2,    -2,     2,     5,     5,     7,   -12,    -7,    -5,    -3,   -15,   -10,     4,    -2,    -8,    12,     0,    -9,   -19,    -1,    11,    13,    16,     9,    -5,    -7,    16,    15,     0,     2,     1,     6,    15,     6,    -2,    -4,    -2,     9,     1,    -4,     9,     1,    -5,    -4,   -12,    -9,   -15,    -5,   -12,    -2,    17,     7,    -9,   -21,     5,     3,    -2,     1,     2,     2,    -6,    -5,    -1,     3,     1,     9,     5,     5,    10,     4,     5,    -8,    -4,    -3,   -18,   -15,   -16,    -2,    13,     9,    16,    20,    -5,    -4,    -1,     1,    -1,     3,    -7,     3,     1,     8,     3,     6,     2,     3,     4,    -1,     3,     3,    -4,    -8,    -6,     3,     7,     9,    15,    17,    19,    11,    -1,    -3,    -7,    -6,    -1,     0,    -4,    -5,    -6,    -7,    -3,     3,    -8,     2,    -4,    -2,     6,    -9,   -19,   -15,     3,    10,    11,     7,     1,     1,     0,     5,    10,     2,     7,    -1,    -2,     8,     8,    -9,     8,    10,     3,     1,    -8,    -2,     4,     4,     5,   -11,   -14,   -21,    -4,     7,    -2,    -2,    -4,   -11,     1,    10,    14,     3,     7,    -1,    -2,     8,     3,     0,    13,     6,    -8,     0,    -3,    -9,     3,     0,     5,    -6,   -16,   -18,    -4,    -5,    -2,    10,   -11,    -7,     0,     5,     5,     6,     0,    10,     7,    -3,    -1,     0,   -11,   -18,    -6,     1,    -4,     1,    -3,     5,    -7,     0,    -4,   -15,   -16,   -14,    -5,     6,     4,     4,     5,     7,     7,     2,     1,     8,     9,     1,     0,     1,    -9,   -21,    -4,    -1,    -6,     4,    -6,    -2,    -2,     6,    -7,    -5,   -13,     1,     9,    15,     5,    10,     7,     9,    13,    20,     2,    -2,    -2,    -2,     1,    -7,    -2,    -7,    -9,     8,    -5,    -2,     5,     0,     1,     4,    -2,     2,     3,     5,    12,    15,     1,    -1,    -3,     6,    10,    20,    -1,     0,     1,    -2,    -3,    -6,   -11,    -3,   -10,    -6,   -10,   -17,    -5,    -8,   -19,     7,     6,    -2,     3,     2,    25,    17,     3,    -1,     3,    -4,     3,     5,    -1,     2,     2,     0,    -1,     0,    -1,    -2,    -2,    -8,     5,   -17,    -9,   -13,   -11,   -11,   -18,    -7,   -11,    -7,    -8,   -10,    -8,    -5,    -4,    -3,     1,    -2,     2,    -1,    -2,    -1,    -2,    -4,    -8,   -11,    -5,    -7,    -8,     3,    -2,   -13,   -13,   -17,   -17,   -14,   -10,    -2,    -5,    -3,    -2,    -1,     1,    -2,     1,    -2,     1,    -1,    -1,    -2,     1,     2,     1,    -1,    -1,    -1,    -2,    -2,    -3,     2,     2,     3,    -1,    -2,    -1,    -2,    -2,     0,     1,    -2,     2,     2,     1,     1,     2),
		     2 => (    0,    -2,     1,    -2,    -2,     1,     1,     1,     0,     2,     1,    -2,     0,     1,     0,     1,     0,    -2,    -1,     0,     0,     1,     0,     1,     1,    -2,    -1,    -1,     0,     1,     0,     0,     2,     2,    -2,     2,    -5,    -7,    -5,    -4,    -2,   -11,    -8,    -3,     0,     3,    -1,    -2,    -3,    -2,    -2,    -4,     1,     1,     2,     2,     1,    -2,     0,    -7,    -7,     0,     2,   -13,    -3,    -5,    -6,    -9,    -5,   -25,    -7,    -1,    -4,    -6,   -10,   -13,   -10,    -2,    -6,     1,     3,     5,     2,     2,    -1,     2,    -4,   -10,   -10,     0,    11,    -5,    -2,    10,    11,     1,   -11,   -14,    -8,   -14,   -13,    -5,     7,    -4,   -14,    -8,    -2,    -6,    -7,     3,    -2,    -2,    -2,     2,    -1,     6,    -3,    -7,    -1,    11,     2,    -1,   -11,    -8,    -7,   -16,   -16,   -10,     4,     4,     1,    -5,     5,     8,    -2,   -12,     2,     1,    -7,    -3,     0,     2,    -4,     2,    13,     3,    -1,    -1,    -2,    -4,   -12,   -17,   -18,   -17,   -14,    -6,    -2,     1,     8,     9,     6,    11,     3,    -9,    -7,     1,    -7,    -2,     2,     2,     4,     1,     2,    -3,    -3,     6,     3,    -4,    -4,    -7,    -3,   -17,   -13,   -12,    -7,    11,     4,     7,    -3,     3,     2,   -14,   -12,    12,    -7,    -1,     1,     2,    10,     1,    -1,    -6,    -1,     7,    -1,     3,     0,     5,     4,     8,    -6,    -7,    -5,    -4,   -13,    -3,     4,     3,     1,   -23,    -3,    17,    -9,    -1,   -13,    12,    11,    -7,    -5,     4,     0,    -4,    -7,   -14,     1,     9,     0,     4,     6,   -16,   -20,    -7,    -9,     2,     5,    -2,    -1,     2,     3,     8,   -12,    -3,     0,    -6,    13,    -6,   -11,    -2,    -2,     0,    -9,    -6,     4,    -5,    -8,     1,     4,     2,    -6,    -5,    -2,    10,     3,     5,     4,    -2,    -2,   -12,     9,    -4,    -2,    -4,    10,   -13,    -7,     7,     6,     9,    -1,     0,     3,     1,     6,    13,    24,     8,    -9,    -5,     1,    11,     4,     6,     2,   -11,    -6,    -9,     6,    -6,     2,   -10,    -7,    -9,     6,     2,     6,    13,    11,     6,    -7,    -5,   -14,    -4,     1,     1,     0,   -11,    -1,     7,     0,     3,     2,   -11,     0,    -4,     4,   -10,    -2,     1,   -20,    -6,    11,     8,     7,     7,     0,     3,     1,   -15,   -17,    -9,    -7,    -7,    -9,    -8,    -7,     3,     5,     1,    -1,   -18,    -3,     3,    15,    -1,    -1,     1,    -1,     8,    -3,    -9,   -13,   -13,   -24,    -7,    -6,     0,    -9,   -16,   -10,   -13,    -7,    -1,    -1,    -2,    -5,   -10,    -4,    -4,     6,     9,    22,     3,    -2,    -1,    -4,     1,   -13,   -18,    -6,    -8,   -15,   -17,   -13,     4,     6,   -11,   -17,    -6,     6,     4,    -3,    -6,   -16,   -11,     2,     4,     0,     9,    17,     6,     2,    -3,     2,     3,     4,    -4,    -9,   -20,   -10,   -12,     4,     2,     9,     5,     0,     5,    -5,     5,     5,     0,    -3,     0,     1,     3,     4,     4,     6,    10,    -1,     1,     1,     6,     9,     4,    -6,     1,    -4,    -3,     2,     3,     6,     0,    11,    13,    11,    17,    -1,   -12,   -22,   -12,    -5,    -3,    -5,     3,    11,     9,     2,    -3,     7,     8,     1,     7,    -1,    -7,    -1,    -4,     6,    -4,    12,    -1,     1,     1,     4,    -2,    -6,   -10,    -5,    -2,     2,    -3,     1,    -1,    10,    15,     1,     0,    -8,    16,     9,    17,    11,    -1,    -7,    -3,    -2,    -8,    -3,     5,     4,    10,     5,    -1,    -3,    -4,     0,    -4,     0,    -1,    14,     2,    13,    23,     2,    -2,    -2,    14,    18,     8,     7,     3,    -2,    -4,    12,     6,     6,    -2,    -2,     4,     7,     6,    -1,   -10,    -6,    -1,     8,     5,    16,     9,    17,    18,    -1,     2,     3,     7,    10,    10,    11,     8,     3,     1,    -1,     0,    -8,     0,     0,    10,     6,    -4,    -3,    -1,    -6,     0,    -4,     8,    15,     4,    17,    -2,    -1,     4,     2,    -1,     9,    14,    -3,    -5,    -3,    -3,    -5,    -8,    -8,   -19,    -9,     3,     2,     7,    16,    12,     7,   -11,    -1,    10,    11,    10,    14,     0,     0,    -2,     7,     4,    12,     0,   -10,   -11,    -8,    -7,   -10,   -13,   -15,   -20,    -8,     1,    -3,     7,     7,     3,    -7,    -3,    -2,     3,    10,    -7,    -9,     0,    -2,     0,     4,     5,     6,     2,    -1,    -4,    -2,   -10,   -13,   -12,   -18,   -14,   -11,     2,   -16,   -29,   -10,     1,    -1,     2,    -8,    -9,    -2,     5,    -3,    -2,     2,     2,    -6,     4,    -7,   -10,    -2,    -6,    -2,   -19,   -20,   -18,   -17,   -20,    -9,    -8,   -22,   -33,   -17,     5,     2,     5,    -7,    -4,     7,     0,    -1,    -2,     0,     1,    -1,    -5,   -10,   -14,   -14,   -11,   -14,   -16,   -17,    -9,    -6,   -16,     3,    -5,   -13,   -12,   -25,   -22,   -11,     1,    -8,   -10,    -4,     2,     2,     0,     1,    -2,    -1,     1,    -8,    -8,    -8,    -9,    -6,   -20,   -10,    -4,    -5,    -8,    -4,   -12,   -11,   -15,   -19,   -21,   -15,   -13,   -13,     0,    -2,     2,     2,     0,     2,     2,     1,     1,     0,    -2,     0,     0,    -2,    -2,    -9,    -6,    -1,    -7,    -5,    -6,    -5,    -4,    -4,    -5,   -15,   -16,    -6,     0,     1,    -1,     2,    -1),
		     3 => (    0,    -2,     0,     2,     0,    -2,     2,     2,     2,     0,    -2,    -2,    -1,    -3,     0,     0,     2,     2,     2,     1,    -1,     0,     1,     2,     2,     2,    -1,    -2,     1,     1,     2,     1,     2,    -1,    -2,    -1,    -2,    -1,     1,    -2,    -4,    -1,    -2,    -5,    -6,    -5,     1,     1,     2,     2,     0,     0,     0,    -2,    -2,    -2,    -1,     2,    -2,     2,    -1,     2,    -3,    -3,    -2,    -9,   -10,    -3,    -9,   -11,    -7,    -8,   -14,   -17,   -15,    -8,   -21,   -18,   -20,    -6,    -2,     0,     0,     2,     2,    -2,     2,    -3,    -2,    -6,    -3,    -7,    -7,    -7,   -11,    -8,    -1,    -2,    -9,   -10,     2,    11,     7,    -5,    -3,    -5,   -15,   -19,    -9,    -2,    -1,    -1,     1,     3,    -2,     4,    11,     5,     0,     7,     9,    14,    11,    -1,     0,     5,     9,     2,    -9,    -3,     7,     1,    -2,   -17,    -8,   -32,   -21,    -1,    -6,     1,     1,     0,     1,    -4,     4,    -6,    -7,   -10,     3,    -8,     5,     4,     1,    -1,    -2,     0,     0,     4,     8,     3,     3,     8,     3,    -5,    -7,    -6,    -6,     0,     2,     2,     1,    -2,    -6,    -3,    -2,     0,     6,     0,     2,    -2,     4,    16,     6,     0,    -2,     0,     1,     9,   -10,    -6,     2,     0,     0,    -9,   -11,    -1,     1,     4,     0,    -9,    -5,    13,     1,    -1,     2,     0,     6,    10,     2,    -5,     3,     7,    10,    -1,    -2,     1,    10,    -3,    -8,   -16,   -10,   -14,   -10,    -2,     2,    -1,     2,    15,     7,     4,    -7,     8,    -2,   -12,     8,     5,    11,     3,     0,    -5,    -3,     4,    -1,     1,     6,     7,    -3,   -25,   -29,    -8,   -12,    -2,    -2,    -7,    19,    15,     3,   -17,    -5,    -2,    -7,    -2,   -11,    -8,   -19,   -24,   -37,   -16,     4,     1,     4,     6,     7,     3,     2,   -18,   -37,   -15,   -16,     1,     1,    -4,    24,    11,    -9,   -18,   -21,   -30,   -25,   -27,   -25,   -44,   -36,   -33,   -13,    -4,     1,    -5,    -3,     2,     2,     9,     5,    -7,   -33,    -9,    -9,    -3,     1,    -3,    -3,    -6,   -14,   -19,   -29,   -21,   -29,   -39,   -27,   -23,   -11,     9,    13,    13,     1,     5,     0,     7,    16,    11,     7,   -18,   -17,   -14,    -6,     0,    -2,    -1,    -9,   -13,     4,    -5,    -4,   -13,    -6,   -12,    -5,     2,    14,    12,     9,    -4,     1,    -4,     7,   -12,    -3,    -1,    -4,    -6,     1,    -2,    -3,    -2,     1,     0,   -12,     2,    15,    10,     0,    -6,     1,    -5,     3,    11,     6,     9,    -4,    -1,    -1,    -9,   -11,   -16,   -10,    -2,    -5,    -1,   -10,   -10,    -4,    -3,    -3,     3,    -1,     0,     2,    13,    -5,    -9,    14,     4,    -1,     5,     5,     5,    -1,     1,    -1,    -3,    -1,    -7,   -12,    -3,   -10,   -12,   -14,   -25,    -7,    -4,    -4,     7,    10,    -3,     8,    -3,   -17,   -22,   -13,    -9,     2,     4,     0,    11,    10,    -3,    -3,     2,    -2,     1,    -4,    -1,   -14,    -2,   -10,    -8,    19,     0,    -2,     1,     9,    10,     6,     0,   -27,   -20,   -29,   -17,    -9,     2,    -2,     6,    -3,    -6,     1,     0,     0,     5,     3,     7,   -10,    -6,   -16,    -8,     7,    -2,     0,     4,    12,    -1,   -13,    -4,   -19,    -6,   -21,   -39,   -47,   -19,   -21,   -21,   -11,    -8,     5,     5,     5,     0,    -3,     6,     2,    -8,   -16,   -16,    -7,    -3,    -5,     3,    17,     4,   -10,     7,     2,    12,    -1,    -5,   -16,   -11,   -24,   -22,    -9,     4,    -4,     0,    -3,     5,     8,     6,    -1,   -20,   -29,   -10,    -7,    -6,    -2,    -3,   -11,    19,     3,     3,     5,     2,     6,    -5,    -5,   -11,    -8,     5,    -1,     0,    -2,    -3,    -1,     0,    -3,    -6,   -10,   -13,   -21,    -9,    -8,    -4,    -2,     2,   -20,    15,    13,     1,    -1,     0,     8,     1,     5,     5,     4,     5,    -4,    -8,    -1,     0,    -4,    -4,    -1,    -9,   -15,   -19,   -18,    -5,    -4,    -1,    -5,     2,    -3,     7,    15,    -1,    -6,     4,    12,     0,     8,     3,     1,    -7,    -5,    -9,   -10,     3,    -2,   -13,    -6,    -6,   -10,   -21,   -16,    -6,     0,     1,    -1,    -4,    -1,     6,     5,     7,    -5,    -9,    -2,    -7,    -1,    -2,    -8,    -5,    -7,    -4,    -2,     6,   -11,    -2,   -12,   -14,   -20,   -19,   -16,    -7,    -2,    -1,    -2,     2,    11,    10,     2,    14,    -9,     3,    -6,    -2,    -4,     3,    -3,     0,     4,    -1,    15,    -1,     0,    13,    -7,   -16,   -27,   -21,    -9,   -14,    -1,     0,    -1,     0,    -2,     4,    -5,    -6,     2,    -5,    -5,     3,    -4,    -6,    -6,   -13,    -3,    -9,    -7,   -12,    -5,   -16,   -17,   -14,   -16,    -6,    -8,    -1,     1,     0,     0,     1,     1,   -10,    -4,    -2,    -7,   -13,    -8,    -2,     4,   -12,    -1,    -2,    -7,   -18,   -18,   -17,    -6,    -4,     0,    -6,   -15,   -10,     1,    -3,     1,     0,    -2,    -2,     0,    -7,    -3,     2,    -7,   -13,   -18,   -20,    -7,   -13,     5,    12,     8,     1,    -8,   -10,    -6,    -8,   -13,    -8,   -11,    -1,     2,    -1,     1,    -2,     1,     1,     1,     1,    -1,    -1,    -3,     0,     0,    -6,    -1,    -4,     1,    -3,    -7,    -1,    -8,    -7,     1,    -1,    -5,    -2,    -2,    -1,     0,     2,    -1,     0),
		     4 => (    1,    -1,     1,     0,    -1,     2,     2,    -2,    -1,    -1,    -2,     0,    -4,    -4,    -4,    -1,    -1,    -2,    -1,     2,     1,     0,     1,     0,    -2,    -1,    -2,    -1,     2,    -1,     1,    -2,    -1,     0,    -7,    -9,    -3,    -4,    -9,    -3,   -10,   -16,    -7,    -8,    -9,    -6,    -2,     1,    -6,    -3,    -5,    -7,     1,     1,     2,    -1,     1,     0,    -1,     2,    -9,    -2,    -9,   -11,   -16,    -7,    -8,   -17,   -11,   -11,    -7,    -6,   -15,   -12,   -12,    -3,   -15,   -13,   -12,   -10,    -3,    -9,     2,    -1,    -2,     1,    -1,    -7,   -18,    -9,   -13,    -8,    -8,   -11,    -6,   -11,   -12,   -11,   -10,   -11,   -18,   -22,   -11,    -2,     1,    -2,    -5,    -3,   -10,    -6,    -2,    -1,    -2,    -1,    -4,   -16,    -2,     3,    12,     3,    -5,   -16,   -10,    -5,    -4,   -14,   -24,   -19,   -11,   -18,   -10,    19,     9,     3,    12,    -7,    -8,    -4,    -8,    -2,    -2,    -1,    -8,    -6,    -1,     3,    11,    -4,    -3,    -5,    -5,    -5,    -3,   -21,   -24,     3,   -10,     3,    -8,     3,     1,     2,     2,   -14,    -6,    -4,    -4,    -2,     1,     0,    -1,    -2,    -6,    -5,    12,   -10,     4,     8,     2,    -8,   -16,   -35,   -32,   -18,    -5,     3,    12,     0,     0,     2,   -11,   -15,   -16,    -4,    -1,    -6,     1,   -10,    -2,     2,    -3,    -4,     6,    -1,     2,     3,     4,     4,   -15,   -28,   -38,   -15,    -6,    18,    12,    13,     5,    -2,   -10,   -14,   -14,    -1,    -4,   -14,    -9,   -22,     2,    -2,     5,     5,     7,    -2,     5,    12,    -2,    -4,     2,   -30,   -27,   -12,    17,    11,     7,    -4,   -10,     5,    -2,    -5,    -8,     2,   -13,   -19,    -2,   -14,     3,     2,    13,     6,   -16,    -3,     9,     1,     6,     8,    11,   -15,   -21,    -1,    24,     4,     2,     0,   -12,    -4,    -5,     1,   -15,     3,   -12,   -10,     2,    -7,     0,     6,     4,    -2,   -29,    -7,     4,    10,    -2,     5,    10,   -15,   -17,    11,    11,     2,     9,     7,    -8,   -15,    -9,   -18,   -19,     4,    -1,    -6,     0,   -11,     4,     2,     7,     2,   -10,    -2,     4,     3,     6,     7,     2,   -23,   -24,     2,     6,    -1,     3,    -5,   -14,   -14,    -7,   -13,    -6,     4,    -5,   -15,     2,    -7,     5,     7,     7,     7,     2,     2,   -10,    -6,     6,     0,     2,    -7,   -16,     7,     1,     1,     0,     2,   -10,     0,    10,    21,    21,    17,   -16,   -11,     0,    -5,   -10,     0,    11,     4,    -3,     0,    -3,     5,    10,     0,    -1,    -2,    -6,    -7,     4,    -1,     7,     1,     3,    11,    20,    10,     3,    -2,   -16,     0,    -2,    -1,   -10,     1,     6,    16,     2,    10,     5,    -2,    -1,    -3,    -5,    -3,   -11,     1,    -4,     3,     4,    10,     1,    14,    11,    -2,     6,    -6,    -9,    -1,     2,     2,     3,    -3,    13,    -1,    -1,    10,     0,     1,     0,     3,     2,     9,     6,     9,     7,     3,     4,    10,     0,    -3,     4,    -9,   -12,   -12,     5,    -2,    -2,    -2,   -14,     8,    13,    -7,    -8,    11,     1,    -4,     2,     1,    -2,     3,     9,     8,    -1,    -6,     6,     0,    -2,     4,    -9,   -13,    -2,    -4,    -6,     0,     0,    -2,    13,     9,    20,     0,   -12,     3,    -8,     2,   -11,    -8,    -4,    -6,     2,    -8,   -11,   -11,    -2,   -18,    -6,     3,    -5,    -8,     0,    -3,     2,     1,    -9,    -1,    10,    11,    14,   -10,   -11,   -13,    -7,    -3,    -8,   -11,    -7,    -5,    -6,   -18,   -13,    -6,   -12,   -13,    -5,     2,     2,    -3,    -5,    -7,     2,     0,    -1,     0,    -3,     5,    -1,   -16,    -3,   -17,    -9,    -3,    -2,    -1,   -10,    -1,     3,    -2,   -12,     4,    -9,    -3,    -5,    13,     4,     1,    -6,   -10,    -2,     0,     0,     0,    -3,   -10,   -23,   -15,   -14,    -3,   -11,   -13,    -8,    10,     4,    -1,     3,    -2,    -2,    -3,     7,     1,    -6,    -4,    -1,    -2,    -2,   -20,    -3,    -2,    -7,    -6,    -4,   -13,    -9,   -14,   -11,   -10,    -4,   -11,    -5,     2,     2,    -4,     6,   -11,     3,    -8,    -4,    -7,   -10,   -16,    -4,     4,     1,   -17,    -9,    -1,    -3,    -6,    -2,    -7,    -3,     0,     1,   -13,     3,   -17,   -12,     1,     2,    -6,    -2,    -6,    -1,    -5,    -3,   -11,    -9,   -14,     2,     7,    -1,     2,     4,    -1,    -2,    -2,    -4,    -7,     0,    -5,     8,     7,     2,   -21,    -2,    -7,    -7,    -6,    -5,    -7,     1,     1,    10,   -10,   -13,    -2,    -5,     4,    -6,     4,     1,    -1,    -2,     2,    -1,     2,   -17,    -5,    -7,    -5,    -1,    -4,   -10,    -4,    -9,    -6,    15,    -2,     9,     9,    12,   -11,    -1,     2,    -2,    -1,   -15,     1,    -4,    -1,     1,    -2,    -1,    -2,    -1,   -11,   -29,   -17,   -12,    -8,   -12,   -11,   -11,     2,     4,   -10,    -1,     5,     1,    -6,    -2,     7,    -8,     4,    -7,    -3,    -3,     2,    -2,    -1,     2,    -3,    -5,    -2,    -8,   -13,     3,    -3,   -15,   -25,   -22,   -17,    -8,   -13,   -22,    -5,   -14,   -18,   -22,   -21,   -17,    -4,    -6,    -1,     2,    -1,     2,     0,    -1,    -1,    -1,     1,    -8,    -7,    -9,   -10,    -8,   -17,    -9,    -7,   -19,    -6,    -8,   -11,    -8,   -12,   -14,   -13,   -10,    -3,    -1,     0,     0,     2),
		     5 => (    2,    -1,    -1,     1,     2,     0,     1,     1,    -1,     2,     2,     0,    -1,     1,     0,     2,    -1,    -2,     1,     2,    -2,    -1,     1,    -1,     1,     2,     1,     2,     2,     1,     2,    -2,     1,    -2,     0,     1,     2,     2,     2,    -2,    -5,    -5,    -5,    -5,    -3,    -5,    -2,    -1,    -3,    -1,    -1,     0,    -2,     2,    -2,     2,     2,    -2,     0,    -3,    -2,    -2,     1,     1,    -3,    -1,    -9,   -18,   -16,   -22,    -8,     8,     8,    10,    14,    11,    14,    11,    11,    12,    -5,    -3,     1,    -2,     2,     2,    -1,     4,     9,    -2,    -6,    -5,    -4,   -12,   -14,   -11,    -4,   -11,     9,    -4,   -17,   -13,    -1,    -3,     4,     7,    -5,    -2,     7,     6,     7,     3,     1,    -4,    -5,     1,   -13,   -13,   -16,   -19,   -26,    -8,   -20,   -13,   -13,     0,    13,     1,     5,    -1,     0,    -1,     3,     7,    10,    11,    14,    27,     7,    -2,     0,    -2,    -3,    -2,   -12,   -11,   -23,   -22,   -27,   -14,    -2,    -1,     5,     0,     2,    -3,     4,    10,     6,     2,    19,    16,     9,    16,    18,    25,    12,    -4,     1,     0,     5,    -4,   -12,   -21,   -21,   -13,    -6,   -12,    -3,     2,    12,     1,     0,     1,     5,     9,    19,     3,    16,     0,     1,    15,     5,    12,     8,     2,    -1,     2,    -2,    -7,   -10,   -14,    -6,    -1,    -4,     1,     0,    11,     8,     3,    -4,    -6,     2,     7,     8,     1,     9,     0,    -9,    -2,    -5,     5,     6,     4,    -2,    -3,    -7,    -6,    -8,    -5,   -13,    -6,   -10,   -14,     5,    14,     8,   -10,    -9,   -15,   -31,   -17,   -16,   -40,   -19,   -22,   -15,    -6,    -3,    -2,     4,     1,     0,    -4,   -15,   -17,   -16,    -2,   -15,   -17,   -14,    -8,    -7,    -4,    -5,    -9,   -17,   -38,   -48,   -55,   -60,   -58,   -40,   -31,   -28,   -16,   -10,    -8,     0,     3,     1,    -3,    -1,    -9,    -1,    -5,    -9,    -6,    -1,    -6,    -7,     2,    -7,     1,   -12,    -4,     1,   -12,   -34,   -36,   -35,   -29,   -27,   -18,   -10,     0,     2,     1,    -1,    -1,    -1,    -6,    -2,    -6,   -10,   -11,    -8,   -10,    -8,    -5,    -4,     0,    -6,    -5,     4,     1,     5,    -6,   -17,   -29,   -21,   -10,   -11,    -2,     3,    -5,     1,    -2,     0,    -6,    -1,    -5,    -5,    -9,    -5,    -8,    -4,     4,     4,     3,     3,     1,     2,    -5,    -5,     0,    -5,   -10,   -15,   -11,    -4,    -4,     0,    -7,    -1,     0,    -2,    -2,    -1,     4,    -7,     2,   -11,     4,     8,    15,     6,    -3,     6,     1,    -1,    -3,    -7,     2,     1,     6,    -6,    -4,    -8,     0,    -1,    -4,     4,    -2,    -1,     2,     8,    -8,   -14,   -12,    -3,    -4,     9,     1,     0,    -5,     2,   -10,     8,     1,     1,    -9,     0,     1,     0,     0,    -3,    -3,    -4,    -4,     0,    -7,    -5,    -3,     7,    -9,   -14,   -10,   -12,    -7,    -6,    -3,     5,    -6,   -11,    -3,    -9,     5,    -3,    -2,    -7,     2,    -1,     3,     2,    -2,    -2,    -1,     0,     2,    -6,     2,     0,   -12,   -13,   -20,   -20,   -33,   -26,   -16,     3,     2,    -9,     4,     3,    17,    -3,     5,     3,     4,     6,    -8,   -11,    -7,    -7,    -7,    -1,    -5,   -13,     3,    -6,    -8,    -9,   -20,    -9,   -25,   -35,   -12,   -14,   -19,   -14,     4,    -5,    -7,    14,     8,     9,     6,    -4,    -6,   -15,    -8,    -3,    -5,    -1,    -3,     1,     7,     0,    -7,   -11,    -3,     8,    -5,    -1,    -9,   -26,   -13,    -1,    -6,     3,     0,    10,    -5,    -1,     4,    -1,    -5,   -15,     2,   -13,   -10,     0,     0,    10,    -1,     2,    -9,    -2,    -3,     5,     9,     3,     8,     6,     3,     5,    -2,     5,    -2,     4,     3,     3,    -5,     0,    -8,   -13,     1,    -4,    -5,    -2,    -1,     7,     4,    25,    -1,     3,    -1,    13,     9,     1,     4,   -10,    10,     9,     4,     1,     0,    -5,     7,     5,    -6,     8,   -15,   -10,    -6,    -2,     1,     1,    -3,    -7,    -4,    16,    13,     0,    -3,     3,     1,     5,     8,     4,     6,    -2,     4,     5,    -6,    -9,     6,     9,    10,     9,     1,    -5,    -8,    -1,    -2,     2,     1,   -10,     2,    -7,    -4,    -7,    -4,    -5,    -4,    13,     2,     6,    -6,    -1,    -5,     1,    -3,     4,     2,    12,    -5,    -5,    -6,    -9,    -7,    -1,     1,     0,    -2,     5,     6,    -8,    -7,     3,     1,    14,     7,     2,   -11,    -5,    -4,    -1,    14,    -2,   -14,   -12,   -10,   -12,   -10,     1,     4,   -20,   -20,     3,     0,    -2,     0,    -9,    -1,    11,     9,    27,    13,    -2,     8,    17,     0,     5,     3,    10,    -8,   -13,    -7,   -10,   -12,    -2,     7,     9,    -2,     0,    -6,    -7,     2,    -2,     0,    -1,    11,    -5,    -1,     9,    13,     4,    11,     9,     8,     4,     2,    -7,    -3,    -6,   -13,     3,     6,     2,     3,     7,     1,    -1,     1,    -1,    -1,    -1,     2,     2,     0,    -5,    -6,    -3,    -1,     1,    -2,     6,     5,     4,    -4,    -5,    -3,    -2,    -3,    -3,    -2,     2,     1,     4,    -2,     1,     1,     1,     0,     0,    -1,     1,    -2,    -1,     0,    -2,     1,    -1,    -2,     2,    -1,     1,     2,    -3,     1,    -2,    -2,    -4,    -4,    -4,    -4,    -3,     2,     1,     0,     2,    -2),
		     6 => (   -2,    -1,     1,     1,     1,    -2,    -2,    -2,     1,     2,     1,     2,     6,     3,    -1,     1,     1,    -1,    -2,     0,     0,     1,    -2,    -1,     1,    -1,     2,    -1,     2,     2,    -2,    -2,     1,     1,     4,     5,     9,    13,    11,     5,    11,     8,    -4,     0,     5,    10,     1,     8,    10,     8,     7,    10,     2,     1,    -2,     2,     2,     1,     3,     7,    11,     6,     8,     8,     2,    -2,    -7,     9,    14,     6,     7,    18,    10,     4,     6,    -2,    -3,    -1,     2,    -1,     4,     4,    -1,    -2,     1,    -1,     0,    22,    12,    -3,    10,    15,    -3,     2,    -7,     4,     4,    10,     5,    -4,    -4,     0,    -8,    -1,     7,     0,    -1,    -3,    -3,     0,     2,    -2,     0,     1,    -8,    10,    -1,     6,     6,    -5,     1,     0,     5,     7,    -8,    -1,    -2,   -11,    -6,    -7,    -8,    13,    11,     5,    -6,   -13,    -7,    -7,    -2,     5,    -2,     1,     2,    -4,     0,   -15,   -11,    -5,    -8,     9,     0,    -7,     5,     8,    -4,    -5,   -12,     3,     4,     7,     3,     0,    -7,   -11,    -8,    -3,     3,     5,    -2,    -3,     3,   -11,   -10,   -19,   -15,    -3,    -8,     0,   -12,     9,    12,     2,    -2,    -4,    -4,   -10,     4,    -1,   -11,    -1,   -13,   -17,    -3,    -5,     7,    -2,    -1,    -3,     1,   -10,    -9,   -24,   -15,    -7,    -3,    -3,     3,    14,    10,     1,     6,    -8,   -10,    -9,   -24,   -19,   -19,   -11,   -16,   -20,   -12,    -8,     5,   -12,     1,    -1,     2,   -11,    -8,   -26,    -4,    -4,   -11,     7,     3,    -2,    11,     2,    -9,   -17,   -17,   -28,   -25,   -24,   -16,   -19,   -31,   -24,   -20,   -14,    -4,   -11,     2,    -2,    -5,    -7,    -6,   -28,    -1,     2,    -2,    -8,    -7,     1,    -5,   -11,   -11,   -21,   -20,   -29,   -29,   -25,   -15,   -27,   -26,   -18,    -5,    -5,    -6,    -4,    -2,     1,    -3,    -8,   -13,   -25,   -15,     1,     6,     0,    -7,    -1,     6,    -9,   -25,   -23,    -6,     7,    -1,   -12,    -9,    -7,   -12,    -5,    -4,     7,    -9,   -11,     2,     0,     2,   -15,   -11,    -4,   -11,     0,     8,    -6,    -2,     2,     5,   -20,   -18,    -5,     6,     8,     6,    -7,     0,   -17,    -8,   -12,   -11,    -2,   -15,    -8,     2,    -2,     3,    -8,   -10,   -11,    -6,    10,     6,    -2,    -7,     0,    -7,   -27,    -8,    -2,    10,     4,    -1,     7,     9,    -2,    -6,    -8,    11,    -4,    -9,    -8,     1,     0,    -6,    -5,   -17,   -15,     0,    12,     6,   -15,   -11,     0,    -5,   -11,    -9,     1,    -2,    -3,    -1,    10,    15,     7,    -3,     4,     3,    -4,    -9,     6,     0,     1,    -1,   -12,   -20,    -8,    10,     7,     3,    -4,     4,    12,    -3,    -3,     5,    -2,     5,    -8,     7,     6,     4,     8,    10,     3,    -3,     1,    -6,    -2,     1,     0,    -3,   -10,   -15,     0,    15,     9,    -3,     0,    -3,    16,     2,    -7,    10,    -4,     1,    -4,     6,     2,     2,     6,    12,     5,     0,     4,   -12,   -16,    -2,    -2,    -3,    -8,    -6,     9,    18,    -2,    -3,   -14,     8,    13,    -2,    -9,    13,    -3,    -3,     0,    -2,    -2,     5,    11,     7,     1,     3,     0,   -15,   -14,     2,     0,     0,    -5,    -1,    -6,     8,     4,    -8,    -8,    -1,     6,     3,    -3,     2,    -1,    -3,    -8,     4,    -5,    -8,    10,    11,     1,    13,    12,    -6,   -13,     1,     0,     2,    -9,     0,    -5,     3,     8,     0,   -11,     1,    -2,    10,     4,     7,   -10,    -4,    -9,    -3,     5,    -3,    12,     4,     9,     8,    16,    -8,   -13,    -2,     0,    -1,    -9,     7,   -14,   -10,     5,    -2,    -6,    -9,     2,     7,     7,    10,     8,     1,     1,    -7,     3,    -8,    -4,   -10,     9,     4,    11,    -4,    -1,     1,    -3,     0,    -9,     4,    -6,   -10,     0,   -14,    -6,    -4,     0,    -5,     1,    14,    15,     3,     1,    11,    -3,    -3,    -4,     4,     8,    11,    13,    -1,     1,    -1,     0,     0,    -1,     1,    -4,     2,    -1,   -12,   -15,    -2,   -10,   -16,   -12,     9,    10,    -3,     4,    -1,     2,     7,    -7,     8,    13,     5,     3,     5,     1,     2,     1,    -2,    -4,    -4,    -5,     7,   -16,   -29,   -29,    -2,    -7,    -9,    -8,   -10,    -6,   -16,   -10,     5,   -11,   -10,   -10,     4,    -5,   -24,   -15,     5,    -2,    -2,    -1,    -2,     0,    -8,     0,    -7,   -10,   -12,    -6,    14,     4,   -22,   -17,   -20,   -22,   -22,   -26,   -24,    -5,    -6,   -16,   -13,   -19,   -22,    -7,    -7,     0,     2,     1,    -1,    -1,    -2,    -3,    -4,    -1,    -4,    -4,    -8,     0,    -6,   -12,   -19,   -14,    -9,   -13,   -15,   -24,   -11,   -11,    -5,    -7,   -12,    -8,     1,    -1,     0,    -1,     2,    -2,    -1,     2,    -3,    -4,     1,    -5,    -2,     4,     6,     2,     0,    -1,     0,    -4,    -1,    -7,   -11,    -8,    -7,   -12,    -1,    -1,     0,     0,    -2,     1,    -1,     1,    -1,    -2,    -1,    -2,    -1,     0,     1,    -3,    -1,    -3,     0,     0,     1,     0,    -1,    -1,    -3,    -3,    -2,     1,     2,     1,    -1,     0,     0,    -1,     0,     2,    -2,     0,    -3,    -2,     1,     0,     1,    -1,    -1,     2,     0,     1,     2,    -1,    -1,     2,    -1,     0,    -3,     1,     0,    -1,     1,    -1),
		     7 => (    1,     1,    -2,    -1,     2,    -2,    -2,     2,     0,     2,     1,     1,    -1,    -1,     1,    -1,    -1,     1,    -1,     1,     1,     0,     2,     2,     0,    -2,    -1,     1,     0,     1,    -1,     0,     0,    -2,     1,     1,    -1,     2,    -3,    -6,    -2,    -5,    -6,    -6,   -11,   -11,    -7,    -2,    -1,     3,     4,    -2,     2,     0,    -2,     1,     0,    -2,     1,    -1,    -2,    -2,     1,    -4,    -6,    -2,   -12,   -21,   -10,    -6,    -4,    -3,    -5,    -3,     0,    -1,    -5,    -1,    -2,     4,     1,    -3,     1,    -1,     2,     0,     0,    -3,     0,    -8,   -12,   -10,   -12,    -2,    -2,    -8,   -14,   -18,    -9,    -8,    -8,    -4,     0,    -6,    -4,    -3,    -7,    -4,    -1,     0,     2,    -2,     2,    -1,    -2,    -1,    -5,    -5,    -5,   -15,   -20,   -10,   -21,    -6,     2,    -1,   -11,   -16,   -19,   -21,   -14,   -11,    -8,    -6,   -13,   -19,   -13,   -12,    -8,     0,     1,    -1,     0,   -16,    -4,    11,    16,     9,    15,     5,    -8,     3,     3,     4,     9,     5,     2,    -3,   -11,   -15,   -25,   -17,   -15,   -22,   -34,   -23,    -6,     2,    -2,     1,    -3,   -11,    -2,     8,     8,     8,     3,    -1,     8,     0,    12,     5,     5,    -6,    -9,    -6,   -11,     0,     0,    -5,   -13,   -13,   -26,   -13,   -14,    -5,    -1,     6,     0,     3,     3,     8,     4,    -1,    -1,    -8,     2,    -7,     6,    -3,    -8,   -14,    -7,    -9,   -13,   -12,    -2,   -11,     3,     4,    -4,   -15,   -16,    -6,    -7,    14,     7,     1,    13,    16,     0,     8,     2,     5,     2,    -9,    -6,    -4,    -6,     5,     4,     3,    -1,    -2,     1,     0,    -2,    -6,     0,   -22,   -20,    -7,     0,    10,     3,     7,    11,    15,     5,     3,    17,     5,    -9,   -11,    -8,    -1,    -2,     3,    -6,     0,     6,    -2,     5,     5,     6,    -5,    -7,    -1,    15,    21,     2,    -2,     1,    -5,     6,    -2,     8,    10,     9,    -1,    -1,     2,    -6,    -1,    -5,    -3,    -3,     6,    10,     4,     7,     5,     3,    -3,     0,    10,     6,    18,     0,    -6,     3,    10,    -1,    -4,    13,    19,    12,    10,     1,     0,     1,     2,     2,    -2,    -6,    12,    -6,    12,     6,    -4,    -7,    -9,    -5,   -15,    -4,    14,     0,     2,     2,    -7,   -11,   -20,    -1,    -1,     2,     0,    -8,    -6,    -6,   -14,    -9,    -2,    -6,   -10,     1,     0,    -1,    -2,    -6,    -4,    -3,     2,    10,    16,    -2,     4,    10,   -13,   -14,   -15,    -5,    -5,   -12,   -15,   -17,   -16,   -24,   -26,    -4,    -2,     0,    -4,    10,     4,     6,    -4,     3,    15,     6,     6,   -11,   -10,    -4,    -4,    -4,   -11,   -10,   -17,   -12,   -17,   -27,   -21,   -19,   -19,   -22,   -12,     2,     1,     5,    -1,     6,    10,    13,    -7,     2,    -2,    -7,   -18,   -13,    -3,     0,     0,    -6,    -1,   -18,    -8,    -7,   -23,   -12,    -9,    -1,    -2,     4,     0,     7,     8,    -5,     5,     3,    -4,    13,     2,     7,    -3,    -5,   -23,    -9,    -4,    -2,    -4,    -5,    -4,   -12,   -11,   -11,   -15,     1,     9,     9,     8,     9,     6,     6,    -8,    -7,    -1,    -2,     3,     0,     4,     7,    -8,   -26,   -25,   -11,    -7,    -1,    -2,    -1,    -8,    -8,   -10,   -14,   -18,     0,     2,   -10,    -1,     1,     5,     5,    -8,    -6,   -11,     4,     6,     2,    -4,     4,    -6,   -10,     2,    -2,    -5,     3,    -3,    12,    -6,   -12,   -20,   -22,   -14,    -8,   -23,   -15,    -3,    12,    13,   -12,   -12,    -9,    -4,    -2,   -10,    -8,   -11,    -6,   -10,    -9,    -5,     8,    -4,    -1,     4,     2,    -4,   -10,   -24,   -13,   -14,   -11,     4,    -7,    -7,    -1,    -3,    -8,    -6,    -2,   -12,    -7,    -5,    -6,   -11,    -9,   -11,   -19,    -2,   -10,     0,     2,    -3,     0,    -5,   -13,    -3,     2,     6,    -5,    -3,    -3,    -2,     3,     3,   -11,   -14,   -11,   -17,   -17,   -13,    -5,     1,     4,    -1,    -9,    -4,   -16,    -2,    -3,    -3,    -1,   -14,   -10,    10,    12,    -7,     4,     0,    -3,    -8,    -4,     4,   -24,   -16,   -22,   -24,   -14,   -15,   -12,    -2,    -3,   -11,    -9,    -3,    -4,    -3,    -6,    -4,    -4,   -22,     7,    11,    11,    13,    16,     5,     5,     0,    -6,    -9,   -16,   -15,   -16,   -13,   -18,   -13,   -14,     2,     4,   -24,   -14,    -2,    -5,     0,     0,     2,    -6,   -25,     6,    -1,     8,    21,     1,     0,    -3,     6,    -8,    -5,   -15,    -7,   -17,   -28,   -22,   -20,   -19,    -2,     0,   -11,    -8,    -1,   -12,     0,    -2,     0,     5,    -1,    10,    15,    11,     4,    13,     2,    -5,     4,    -4,     5,    -9,    -7,   -24,   -25,   -21,   -13,   -18,     1,    -5,   -19,    -3,    -7,    -2,     2,    -2,    -1,    -4,     9,   -10,     2,     0,     4,    -6,   -11,    -2,     6,    -3,   -13,   -18,   -13,   -16,    -9,    -6,    -9,   -22,    -2,    -3,   -14,     3,     0,    -3,    -2,     2,     1,    -1,   -11,   -13,   -14,    -4,     7,    12,     4,    -7,     0,     4,     8,    -9,    -3,    -1,    -5,     3,    -1,    -7,     7,    10,     4,    -4,     0,     2,    -2,     0,    -1,     0,     2,    10,    10,    -2,    -1,    -3,     0,     7,     5,    -5,    15,    10,     1,     4,     2,     2,    -2,     3,    12,     9,    10,    -1,     2,     0,     1),
		     8 => (   -1,     1,     0,     1,    -1,     2,    -2,     0,     2,    -1,    -1,     2,     0,     0,     0,    -2,    -2,    -2,    -1,    -1,    -2,    -2,    -1,    -2,     0,     0,    -1,     1,     1,    -1,    -1,     2,     1,     2,     2,    -2,     2,     2,     0,     1,     0,    -3,    -2,    -3,    -7,    -6,    -3,     2,    -1,     0,     1,     1,     0,     2,     2,    -1,     1,    -2,    -2,     2,    -2,     2,    -1,    -1,    -3,    -7,   -18,   -16,    -4,    -4,    -3,    -8,   -10,     8,    12,     4,    -8,    -8,    -7,    -7,    -3,    -4,     2,     0,    -1,    -2,    -6,    -5,    -4,    -7,    -4,   -14,    10,     8,    -4,   -11,   -10,    -8,    -7,     3,     2,     2,    16,     8,     0,    -5,    10,    14,     0,    -3,    -5,     2,     0,    -1,    -5,    -8,   -14,   -18,     0,     7,    -2,   -11,   -10,     6,    -3,    -1,     3,     4,     5,     1,    -2,     0,    -6,     0,     6,    -6,   -11,     8,    10,     0,    -1,    -1,    -4,    -8,    -8,   -13,     1,    -1,   -14,    -7,    -5,     0,    -2,     5,    -1,     4,    -5,   -14,   -17,    10,    -2,    10,     1,    -4,    -5,    -1,    -5,    -4,     1,     0,    -8,   -14,   -10,     2,    -2,    -6,   -11,    -5,     2,    -5,    -4,    -5,   -12,     0,    -7,    -7,    -7,     4,     1,    -4,    -4,   -10,    -9,    -7,    -1,    -1,     2,   -11,    -3,    -5,    -1,    -1,    -5,    -5,    -1,    -2,    -9,    -2,    -6,   -14,    -8,     4,    -3,   -10,    -7,     2,     1,    -2,   -10,    -8,    -8,    -1,     3,     7,    -5,    -8,    -2,    -2,    -6,    -1,    -9,    -4,     2,     5,   -12,    -9,    -6,    -2,    -5,    -5,    -8,   -11,    -6,     1,     2,     4,   -13,   -15,    -5,     1,    15,     7,    -1,    -3,    -8,     1,    -4,    -4,    -8,     3,    -1,    -5,   -12,    -1,    -4,    -8,   -11,   -11,    -6,    -6,   -12,     6,     2,   -13,   -14,   -12,   -10,    -1,     5,    -8,     2,    -4,    -7,     0,    -3,     2,    -7,    -7,    -2,     1,     6,    15,    -5,    -6,     4,     1,     1,     1,     4,     7,     1,    -5,   -10,   -15,    -7,    -9,     2,     3,     0,    -3,    -3,    -8,    -5,     6,     4,     0,     4,    10,     5,     2,    -6,   -11,    -4,    -3,     5,    -3,     1,    -9,   -10,    10,    -7,    -7,    -3,   -20,    -1,   -10,    -1,     1,    -7,     0,     7,    10,     6,    -2,     3,     9,     7,    -9,    -6,   -10,    -8,   -11,    -6,    -4,     0,   -11,    -1,     5,     6,     9,     3,   -17,   -18,   -14,     2,    -1,    -9,   -15,     2,     5,    -4,   -13,     7,    20,     8,     6,    -2,    -7,    -9,    -1,     1,   -16,    -5,     0,     5,    12,     9,     9,    -1,   -15,   -24,     3,     0,     1,     0,   -18,    -8,    -3,    -5,   -14,     3,     2,    -2,     0,     2,    -1,    -6,    -6,   -21,    -9,     7,    10,    10,     8,    -4,   -13,   -19,   -14,   -23,     0,    -2,     1,    -4,     5,     2,    -9,    -7,    -7,     1,    -1,     6,     8,    -1,    -1,    -8,   -17,    -6,    -4,    -7,     3,    -3,   -12,   -14,    -7,    -6,     0,   -11,    -9,     1,    -1,    -2,     9,    -2,    -8,    -9,    -8,   -20,   -13,    -4,     5,     6,    -7,    -5,    -4,    -1,    -2,    -1,    -8,    -2,     3,    -7,    -2,     1,    -2,   -13,    -7,     1,    -1,    -5,     7,    -6,    -9,   -11,    -6,   -17,   -31,   -12,     3,     9,    -2,    -1,     2,     2,    -5,   -13,   -12,     2,    -5,    -6,    -6,    -5,    -2,     2,    -4,    -3,     1,    -6,    -7,    -4,    -7,    -9,    -9,    -6,   -11,    -1,    -1,     5,     3,    -5,     6,     5,    -4,    -3,    -4,     1,    -7,    -4,    -8,    -3,    -1,    -2,    -6,     1,    -1,    -4,    -4,    -2,    -6,   -12,   -15,     4,     5,    -1,    -3,     6,     4,    -3,     9,    -7,    -2,     0,     1,    -9,    -7,    -6,    -5,     0,     0,    -8,    -9,     2,    -1,    -4,     0,    -5,    -4,   -15,   -16,    -4,     4,    -3,    -3,    -3,     5,    -7,     1,   -11,   -11,    -4,    -1,   -15,    -6,    -1,     1,     0,     0,    -6,     0,    -4,    -2,    -5,     0,    -6,    -8,   -12,    -2,    -9,    -8,    -5,     4,    13,     4,     5,     2,    -6,    -6,    -4,    -5,    -8,    -7,    -4,    -4,    -6,    -3,    -7,    -2,    -4,    -6,    -3,    -4,    -5,   -16,   -18,   -10,    -6,    -6,   -14,    -7,     8,     6,     6,   -10,    -1,     1,     0,     0,    -4,     0,     0,    -1,    -4,    -3,    -7,    -1,    -2,     0,    -6,    -2,    -2,    -8,   -15,   -20,    -7,    -1,    -7,    -1,    -7,    -3,   -10,    -4,     2,    -7,    -6,     1,     5,     5,     1,    -3,     0,    -1,    -8,     0,     2,    -1,    -1,    -2,    -3,    -6,    -6,   -10,    -7,    -7,   -18,    -6,    -8,    -8,    -4,     6,     5,    -5,     9,     5,     1,    -1,    -4,    -4,   -14,   -10,    -4,     2,    -1,     2,    -3,    -1,    -3,    -9,    -6,    -3,    -6,    -6,   -10,   -13,    -2,     4,    -3,     6,    -1,    -1,     5,     5,     2,   -10,    -3,    -4,     0,    -4,    -1,     1,     1,    -1,    -1,    -3,    -3,    -6,    -9,    -3,    -3,    -5,    -7,   -15,   -18,   -15,   -15,   -22,     0,    -2,    -2,   -19,   -17,   -10,    -7,     3,    -2,    -1,     2,    -2,     0,    -1,    -2,     1,    -4,    -1,    -3,    -2,     0,    -5,    -1,    -5,     2,    -5,     0,     0,     0,     1,     0,    -1,    -1,     1,    -2,    -1,     1,     2,    -1,     1),
		     9 => (   -1,    -1,     2,    -1,    -1,    -2,    -1,     2,     1,     0,    -2,     0,     0,     0,     2,     2,    -1,     0,    -2,     1,     0,    -2,     1,     1,     2,    -3,    -1,     0,     2,    -1,     2,     2,    -2,     1,    -3,    -1,     2,     0,    -1,    -1,    -7,    -4,    -1,    -1,    -2,    -2,    -5,     2,     0,    -3,    -2,    -3,     0,    -1,    -1,    -1,     0,     0,     2,    -1,     1,     2,     0,     0,    -2,    -3,    -3,     0,    -1,    -1,    -7,    -1,    -3,    -1,    -2,    -1,    -6,     3,    -3,    -3,    -2,     2,     0,    -1,     0,     0,     1,    -4,    -1,    -4,    -3,    -1,    -8,    -3,    -5,   -11,    -7,    -2,    -6,    -6,    -7,    -3,     6,    -4,    -6,    -8,    -7,     1,    -4,    -3,     0,    -1,     0,    -2,     0,    -4,    -4,     1,   -11,    -3,    -3,    -1,    -5,    -6,   -15,   -19,   -22,   -21,   -11,    -1,     8,   -11,   -16,   -11,    -8,    -7,    -6,   -14,   -10,     1,     0,     1,    -2,    -3,     1,    -2,    -4,    -6,   -14,    -8,   -12,    -4,    -4,     5,    -5,    -8,   -18,   -19,   -18,   -15,     2,    -8,   -10,   -12,    -7,    -7,   -16,     1,    -2,    -3,     0,    -4,     4,    -7,    -2,   -15,   -12,   -12,   -16,    -6,    -7,   -12,    -4,    -4,    -4,   -12,     1,    -8,     4,     7,     0,    -5,    -7,    -8,   -11,   -10,    -1,    -4,    -6,    -5,    -8,   -13,   -14,   -17,   -20,   -28,   -23,   -18,    -9,    -7,    -9,   -17,     5,     3,    -1,    -2,    21,     8,     8,     6,    -4,   -10,    -4,    -7,    -8,    -3,     2,     0,   -10,    -8,    -9,   -13,   -15,   -22,    -7,   -14,    -6,    -3,   -14,    -5,     2,     8,     8,     1,     1,    -1,    -1,     9,     3,    -6,    -9,    -5,    -2,    -5,    12,    -1,    -5,    -9,    -5,    -2,   -17,    -3,    -3,    -6,    -7,   -13,     3,    10,     2,     1,    -2,     7,    -8,     2,     4,     0,     7,     7,   -20,   -10,     0,    -3,    -8,    -7,    -1,    -6,   -11,   -14,    -5,    -1,    -2,     4,    -6,     4,    -3,    -9,   -10,    -8,   -18,   -16,    -8,    -3,    -6,    -2,    11,    24,    -8,   -15,     2,   -20,    -4,    -3,    -6,    -9,    -8,    -3,    12,     6,     8,    -3,     2,    -4,   -11,   -18,   -20,   -23,   -10,    -4,     6,    -2,     6,     3,    17,    22,    -2,   -13,     1,    -2,     2,   -12,     5,    -6,   -10,    -1,     5,     3,     9,    -5,   -14,   -10,   -17,   -12,    -5,   -18,     0,     0,    11,    -3,     7,     9,    -3,   -17,   -15,   -14,    -2,    -4,    -5,    -9,     6,    -8,    -1,     4,     2,     6,    13,     1,     1,     2,    -8,     7,    13,     1,     0,    13,     5,    14,     2,    -5,   -11,    -7,    -8,     1,     0,    -4,     1,    -8,     6,    -7,    -1,    -6,    13,    13,    12,     0,     5,     6,     5,     8,     1,     2,    -1,     6,    -4,   -14,    -6,   -18,   -16,    -3,     2,     0,    -1,     2,   -15,   -10,     7,    -7,   -10,    -8,     3,    -6,     2,     6,     6,    14,     0,     4,    -2,     1,     8,     3,   -12,   -14,   -19,   -15,   -12,    -3,    13,    -2,    -3,    -4,   -10,    -8,     5,    -5,    -2,    -1,    -7,    -3,     3,     5,    -5,     3,   -10,   -11,     0,     6,     3,    -1,   -17,    -6,    -5,   -18,    -9,    -1,    -2,    -1,     1,    -3,    -8,    -2,    -7,    -8,    -5,     7,    -7,   -12,    -9,    -6,    -4,    -2,    -6,    -3,     0,     9,     7,    -7,    -9,    -4,    -9,   -18,    -7,    10,    -1,    -4,     0,     2,    -8,    -3,   -17,   -12,     0,     6,    -8,   -13,    -3,     4,    -5,    -3,     5,    -6,    -2,    -4,     4,     1,    -8,    -6,    -1,    -7,    -4,    12,    -7,    -7,     0,    -2,    -9,    -6,   -18,   -15,    -7,    -6,   -11,   -16,   -10,   -13,    -1,    -7,    -1,    -9,   -10,    -6,    -3,     1,   -17,    -8,    -1,    -3,     4,    14,    -9,    -6,     2,     0,     6,    -5,   -13,    -8,   -22,   -17,     5,    -7,   -15,    -2,     8,     6,    -3,   -10,    -3,    -1,     1,    -4,    -9,    -8,    -6,    -2,     3,    12,    -2,    -2,    -1,    -2,    -2,    -6,   -13,    -6,   -16,   -11,     4,     5,     1,    -6,    -3,    -7,    -6,   -19,     1,    -4,    -4,     3,    -9,    -7,    -9,    -4,     3,    10,   -10,    -1,     2,     2,    -8,   -13,   -16,   -13,   -20,    -7,     4,     7,     7,     5,    -3,    -8,   -13,   -10,    -6,    -4,   -14,     0,     2,    -8,    -4,     1,     4,    -1,    -6,    -2,     0,     2,    -7,    -9,   -20,   -10,   -13,     2,    11,     8,     2,    -8,    -3,   -12,   -13,    -3,     1,    -2,    -3,    -3,     3,    -1,     2,    -8,    -3,     4,    -5,     2,     2,     2,    -4,    -7,    -9,     0,     1,     6,     3,     8,     3,    -3,     0,   -13,     2,    -9,    -8,     0,    -7,     5,     1,     0,     4,     0,    -1,    -1,    -3,     0,    -3,     2,     8,    -4,     3,    -2,    -4,    -1,     5,     3,     8,    -1,     7,     0,    -8,    -7,     2,    10,     6,     2,    -3,    -5,    -6,     5,     1,    -1,    -1,     1,     2,     3,     0,    13,     6,    -2,     8,     7,    -5,     1,     4,    12,     2,    10,     8,     4,    14,    17,     9,     7,    13,     2,    -5,     4,    -3,     1,     1,    -2,    -1,     1,     2,    -1,    -4,    -3,     4,    14,    12,     8,     8,    17,     9,     8,     6,     6,     3,     6,    10,    13,    -5,    -6,    -3,    -3,     2,    -1,    -2,    -1),
		    10 => (    1,     2,     1,    -2,     1,    -1,    -2,     0,     2,    -1,     1,    -1,    -2,     0,     0,     0,     1,    -1,    -2,    -1,     0,    -1,     0,     1,    -2,     0,     0,     1,     0,    -2,    -2,    -2,     1,     2,    -1,     1,     2,    -3,    -3,     2,     6,     1,    -4,     8,    10,    11,     0,     2,     2,     0,     0,    -1,    -1,     0,    -1,     1,     2,     2,    -3,     9,     8,    -2,    -2,     2,    -3,    -4,    -7,    -1,     0,    -5,    -3,   -12,    -2,   -14,   -12,   -12,   -10,    -4,   -12,    -7,    -6,    -2,    -2,     2,     2,     1,     1,     0,    -3,     0,    -3,    -1,     5,    -8,   -20,   -12,     1,     3,    -2,   -10,    -8,   -16,    -2,     0,     1,    -9,   -10,    -5,    -1,     2,   -17,     0,     2,     2,    -2,    -4,     3,   -13,    -8,   -10,    -7,   -13,   -14,   -11,   -20,   -21,    -4,     4,   -10,     3,    -5,     0,    -2,     1,     4,     3,    -9,   -14,   -15,    -2,    -2,    -2,    -6,    -2,     2,   -15,    -7,   -15,    -5,     0,   -17,    -7,   -13,    -8,    -1,    -2,    -6,    -1,    -6,    -2,   -17,    -8,     9,     1,   -14,    -9,   -12,    -9,     1,     1,   -10,    -1,    -3,    -1,    -6,    -6,     2,    -2,    -5,     1,    -5,     1,     1,    -6,    -4,     0,     2,     1,    -8,     6,    11,    -6,   -14,   -14,    -1,    -2,     0,   -12,    -7,    -4,    -3,     1,    -2,   -10,    -2,    -5,    -2,     2,    -2,    -5,    -4,     2,    -7,     2,     7,     3,   -14,    -1,    -5,    -6,   -20,   -14,   -10,     6,    21,   -17,     9,     4,    -3,    -4,    -3,   -12,    -6,    -6,     0,    -1,     3,   -20,     3,     8,     0,    11,     8,   -10,   -14,    -3,    -6,    -6,   -20,    -8,   -15,    -2,     2,    -4,    13,    -1,    -3,     3,    -8,     2,     4,    -5,     2,    -1,     0,     0,    -5,    -6,     8,     4,     7,    -3,     8,    -4,    -9,    -9,    -8,   -19,   -16,     0,    -1,     1,     8,     4,    -2,    -1,    -2,    -4,    -3,    -2,     3,    -1,     0,    -4,     2,   -17,    -6,     6,    -1,     0,    -4,    -8,     1,    -2,   -12,   -11,   -13,    -1,    -2,    25,    -8,    -9,   -10,     2,     4,    -8,   -16,   -14,    -2,     1,    -3,     4,   -11,   -18,   -14,    -3,     5,     7,    -1,   -15,   -16,   -11,   -15,   -15,    -9,     1,     0,     3,    -4,   -11,     9,    11,     3,    -6,   -23,    -2,     4,     2,     8,    -1,   -14,   -19,    -8,     2,     8,    11,     3,   -12,   -14,    -6,   -12,   -15,    -6,    -2,    -2,     6,     7,    -9,    18,     9,     6,     1,    -8,     7,     4,    -2,     1,   -10,   -24,   -33,   -12,     1,     3,    12,    16,   -10,    -6,     7,     2,    -1,   -10,    -4,     2,     1,    -2,   -12,     1,    11,    -8,     2,     6,     6,     3,    14,    11,    -3,   -17,   -13,   -11,    -8,     6,    16,    14,   -11,     0,    10,    -1,    -6,    -5,    -3,     2,    -2,    -9,   -15,   -10,    -6,    -6,    -2,     5,     2,     6,    12,    24,    -9,   -25,   -13,    -5,    -1,    13,    -3,     6,   -13,    -1,     6,    -3,    -4,   -20,    -4,     2,     1,    -7,    -9,    -7,    -3,   -10,   -10,     7,    -2,    -4,     6,     7,   -18,   -26,    -2,     4,     5,     6,     5,   -10,   -17,   -12,    -4,    -8,   -11,   -17,    16,     1,    -4,    -8,   -11,    -2,    -7,   -14,    -4,     3,    -3,     1,     0,     4,   -15,   -14,    -2,     5,     4,    -4,     4,    -2,   -17,    -7,    -8,    -8,   -10,   -10,    25,    -1,    -3,    -9,    -9,    -9,   -18,   -11,    -6,     1,    -3,     4,     2,   -10,   -12,    -8,     1,    13,     4,     2,    -6,    -8,   -10,     0,    -8,    -4,    -7,   -12,    -6,     1,     7,     0,    -7,   -10,   -10,   -15,    -6,     9,     2,    -1,     2,    -2,     2,    -5,    -4,   -12,    -6,     8,    -4,    -4,     1,    -8,    -9,    -1,   -13,    -8,    -3,    -2,     9,    -4,    -8,    -2,   -10,   -18,    -8,     4,     2,     7,     7,     9,     5,    -2,   -16,   -12,    -2,    -8,     1,    -5,     3,    -9,    -3,   -11,     1,     6,     2,     2,     1,    -5,   -11,   -12,    -6,   -11,    -7,     1,     3,    13,     1,    12,     5,    -8,    -7,    -7,    -7,     2,     6,     0,    -5,   -10,    -2,     0,     3,    31,     7,     2,    -2,   -10,   -17,   -14,    -7,   -12,    -9,    -5,     8,    -1,    -1,     1,   -13,     3,     6,     6,    -8,   -14,    -3,   -13,   -11,    -7,    -5,    -1,     5,    17,     7,    -2,     1,    -1,   -11,   -13,   -21,    -9,    -7,    -8,     9,    17,     6,     3,    -3,    -1,    -8,     1,    -5,     0,    -3,   -13,   -10,    -3,    -3,     0,     0,   -14,     0,    -1,    -1,    -4,     0,     7,     5,   -13,   -17,   -19,   -14,   -12,    -7,    -2,    -9,   -12,    -7,    -9,    -4,     6,   -16,   -10,    -9,    -6,    -2,     2,     3,     1,     1,     2,    -1,    -3,     0,   -10,    -8,    -9,   -14,    -4,    -7,   -18,   -21,   -35,   -34,   -35,   -27,   -16,   -13,   -13,   -13,   -16,   -13,    -7,    -6,     1,    -1,    -1,     1,     2,    -2,     1,     2,    -6,    -9,   -22,    -7,    -9,   -17,   -11,   -13,    -9,    -9,    -4,   -12,   -12,   -13,   -17,   -14,   -13,   -10,    -5,    -6,     0,     1,     1,     1,    -1,    -2,    -2,     2,    -1,     2,    -2,    -4,    -5,     0,    -1,    -1,     0,    -3,    -3,    -3,    -2,     0,    -2,    -1,     1,    -3,    -1,    -3,     1,    -2,    -2,     0),
		    11 => (    0,     1,    -2,    -2,     2,    -2,     2,     1,     0,     1,     2,    -2,    -1,    -2,     2,    -2,     1,     2,    -1,     0,     0,    -2,     1,    -2,     2,    -1,     2,    -2,     0,    -1,    -2,     2,     0,    -2,     0,     1,     2,     0,     0,    -3,    -1,    -4,     0,    -3,    -5,    -4,     0,    -2,     1,    -2,    -1,     2,    -2,     2,    -1,    -2,    -2,    -2,    -2,    -2,    -2,     0,     2,     1,    -4,    -2,     3,     2,     1,    -2,    -3,    -8,   -18,   -22,   -18,     5,     6,    -8,    -3,    -6,    -2,    -2,     1,     1,     1,    -2,     7,     1,    -1,    -2,    -2,     8,     8,    10,     8,     2,     2,     0,     2,   -12,   -19,   -14,    -2,    -6,    -6,   -10,     3,     8,    -7,     0,     0,     2,    -1,     2,     6,     5,     2,     5,     7,     6,    -2,     1,    -7,    -6,    -5,    -7,    -7,   -15,   -11,    -5,     2,     4,    10,     0,     0,    -4,   -12,    -9,   -13,   -11,    -1,    -1,     1,    11,     8,     8,    -2,     0,   -13,    -7,   -11,   -12,    -5,    -4,   -22,   -24,   -16,     2,     5,     3,    -1,    10,     8,     3,     2,    -8,    -9,    -1,    -1,     0,    -2,    10,    17,    -3,    -6,    -1,   -15,     9,     7,    -1,   -22,   -25,   -32,   -26,   -12,    -8,     0,    -3,    -3,     2,     0,     2,    -7,   -10,    -7,    -5,     1,    -4,    -6,     0,    -7,    -9,    -6,    -8,   -17,     0,    11,     1,   -14,   -20,   -22,   -17,    -6,    -3,     6,     0,     1,    -2,    -2,     3,   -14,   -21,   -13,    -4,     0,    -9,    -7,    -2,    -4,    -5,    -5,   -10,   -10,    -4,     1,   -14,   -11,   -12,   -22,   -11,     0,     5,     3,    -1,     5,    -3,    -1,    -1,   -14,   -17,   -13,    -4,    -1,     1,    -7,    -3,    -4,    -6,    -4,    -5,    -5,    -1,   -18,   -20,   -22,   -35,   -31,     0,     8,     2,     4,    -2,    -3,    -3,     1,    -1,    -3,   -10,    -4,    -7,    -2,     1,    -3,    -1,     0,     0,   -11,   -12,   -16,   -10,   -18,   -18,   -24,   -29,   -14,    -1,    13,     2,    -4,    -2,     0,     4,     3,    -1,     2,    -5,    -6,    -5,    -2,     1,     3,     2,    -3,     2,    -5,   -13,   -15,   -12,   -15,   -10,   -14,   -11,    -7,    16,     6,     6,    16,    -3,     0,     2,    -9,   -13,    -9,     1,    -7,     1,    -1,     1,    -7,     4,     0,     5,     2,   -11,     1,   -18,   -11,   -12,    -4,    -8,     4,    12,     1,     6,     2,     4,   -12,    -1,   -10,    -2,    -7,     1,    -4,     0,    -2,     1,    -5,     0,     1,    -6,    -3,    -6,    -5,   -10,    -4,    -2,    -8,     2,    12,     8,     2,     8,     5,    -5,   -27,   -12,   -12,    -4,    -5,    -3,     0,     1,    -1,    -1,    -1,     0,     3,    -4,    -3,     0,    -2,     7,     9,    -3,    -1,     8,     3,     4,     7,   -11,   -15,   -32,   -35,    -4,     5,     0,    -3,    -6,    -4,    -1,     0,    -2,     6,    12,    -1,   -13,    -1,     2,    17,     7,     6,     1,    -3,     2,     2,     6,     2,   -10,   -29,   -36,   -21,    -3,     3,     1,   -23,   -17,   -11,     0,     2,     0,     2,    -4,     4,    -3,    -7,     1,     7,     7,   -10,    -1,    -4,    -1,    -9,     5,     6,    -2,   -20,   -19,    -3,     5,     6,    13,    19,    -7,   -12,    -3,     0,     0,    -1,    -6,     0,   -15,    -7,     4,     0,     0,    -3,     8,     7,    -1,     2,   -10,     2,    -1,     3,     8,    10,    17,    21,    20,    15,    -1,   -21,    -8,     0,     0,    -2,    -1,    -9,   -24,   -15,     2,     1,    -1,    -3,     7,    -3,    -2,     1,    -3,    -7,    -1,     4,     6,     6,    -1,    12,    10,     0,     4,    -1,     6,    -1,     2,     2,    -9,   -15,    -4,     1,     4,     3,    -2,    -5,    -2,    -2,    -9,   -19,   -14,    -9,   -14,   -11,    -7,    -6,    -4,     7,    10,     9,    10,    -1,     3,    -1,    -1,     0,    -7,     3,     8,     7,     1,     3,     0,    -5,     6,    -7,   -14,   -14,   -10,     5,    -7,   -15,    -9,   -10,    -3,     8,     8,    14,     0,     2,     4,     5,     6,     1,     0,    -2,     0,    -1,     2,     2,    -4,    -4,    -2,    -5,    -3,    -4,     3,     7,     6,    -8,    -7,   -10,    -5,     2,    14,    12,     5,     2,     2,     8,     6,     1,     1,     3,    13,     4,     0,     3,     8,    -4,    -7,   -11,    -1,    -9,     8,    10,     0,    -8,   -11,   -10,   -10,     1,     2,     3,     0,     3,     1,     0,     0,    -3,     6,     1,     1,     1,     1,    11,     6,    -4,    -9,     2,     4,     5,     9,     3,    -6,    -7,    -9,    -4,    -1,    -2,    -2,     7,    13,    15,     1,     0,     1,     2,     4,   -12,    -8,   -12,   -15,    -3,     9,    -2,    -7,     9,    14,     2,     1,    -1,     0,     0,    -4,     0,     2,     2,     2,    -8,     2,     0,     1,     0,    -1,     2,    -5,   -10,   -10,    -3,   -21,    -5,     4,    -4,     3,    11,     3,   -15,    -9,    -8,   -14,    -8,    -5,    -3,    -7,    -6,    -5,    -5,    -2,     0,    -1,    -1,    -2,    -1,    -1,    -9,    -7,    -8,   -11,   -14,   -12,    -8,    -4,    -7,    -8,    -6,    -7,    -9,   -10,    -4,     0,    -1,    -2,    -1,    -1,     1,     0,    -2,    -2,     1,     0,    -2,     1,    -1,    -1,     0,     1,     1,    -2,    -8,    -4,    -2,    -1,    -5,    -3,     2,     1,    -2,     0,     0,     0,     2,    -1,    -1,    -1,    -2,     2),
		    12 => (    2,    -2,     2,    -2,     0,    -1,    -1,     2,     1,     1,    -2,     2,     1,    -2,     4,     2,    -2,    -1,     1,    -1,     1,     1,    -2,    -2,     1,     1,     1,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,    -4,    -8,    -3,    -3,    -4,    -4,    -7,    -2,     2,     2,    -1,    -3,    -8,    -5,    -4,    -1,     2,     0,     1,    -2,    -1,     2,    -1,    -3,    -7,    -5,     2,    -1,    -3,     1,     2,     3,     8,     3,    -4,    -3,    -7,    -9,    -5,     3,     3,     1,     2,    -7,    -2,    -4,     2,     2,     2,     0,     2,    -3,   -14,     1,    -7,    -4,    -7,    -1,     8,    14,    10,     8,     2,     1,     1,     0,     0,    -4,     0,     1,     3,    -7,   -13,    -6,    -6,    -2,     1,     0,    -1,    -1,    -6,     2,     4,     9,    13,     1,     0,     4,    11,    10,    12,     0,    -2,     0,    -6,    -1,    -8,    -5,    -7,    -8,    -8,   -13,   -11,   -11,    -2,     2,     2,    -9,    -1,     1,     5,     9,    17,     8,     4,     4,     1,     3,     3,    -5,    -4,    -6,    -4,    -5,    -3,     1,     2,    -3,    -7,   -12,    -5,    -6,    -2,    -2,    -2,     0,     0,    -1,     1,    12,    10,     6,     6,     2,     1,    -3,     0,    -4,    -5,    -4,    -4,    -1,    -7,    -1,     3,     2,    -7,     0,    11,    -6,     1,     2,    -2,    -1,    -1,    -3,     2,     1,     3,     0,    -6,    -5,     0,    -4,    -5,    -3,     2,     3,    -8,    -7,    -9,     1,     5,    -3,    -8,     4,    13,   -17,    -7,    -7,     5,    -3,     1,    -2,     0,    -3,     2,    -8,   -10,    -5,    -6,    -2,     1,    -1,     1,     2,    -3,    -6,    -3,    -2,    -1,    -3,     3,     2,    -1,   -16,    -8,     1,    -7,     8,     0,    -4,    -3,    -5,    -4,    -7,    -9,    -5,    -6,    -1,    -2,     9,     2,    -6,    -2,    -5,    -4,    -1,     3,     3,    -1,    -4,    -9,     0,    -6,     2,    -1,     2,    -2,    -8,    -3,    -6,   -10,   -15,   -13,   -15,    -5,    -2,    -4,    -4,     0,    -9,    -3,   -10,    -3,    -8,     3,     5,    -5,   -10,    -4,     5,    -9,    -1,    -5,    -3,    -8,    -6,    -5,     0,   -14,   -15,   -15,   -14,    -5,    -1,     2,     4,    -4,   -10,    -6,     3,    -1,    -4,    -4,    -3,    -4,    -7,    -3,     0,    -4,    -1,    -3,    -9,   -10,    -4,    -2,    -6,    -8,    -3,    -4,    -4,     2,     7,     0,    -1,    -2,    -5,    -3,    -5,     1,    -9,   -10,    -4,    -8,   -11,     1,     4,     2,     2,    -3,    -5,    -6,    -7,   -10,    -4,    -9,    -6,    -3,     0,    -2,     0,    -1,    -2,    -3,    -7,    -6,     3,     0,    -4,    -4,    -7,    -9,    -2,     3,     8,     0,     0,    -6,    -4,    -3,    -8,   -11,    -2,    -7,    -5,    -6,    -5,    -9,    -8,    -5,    -5,    -7,    -9,    -9,     1,    -2,    -2,   -11,    -8,    -7,    -2,     6,    11,     6,     0,    -7,    -5,     1,    -6,     1,    -6,    -4,     0,    -6,    -3,    -5,    -7,    -1,    -2,    -8,   -14,   -10,    -1,     0,     1,    -4,    -7,    -9,     4,    10,    13,    10,     1,    -4,    -2,     7,     6,     0,    -4,    -5,    -3,    -2,     2,     1,     3,     3,     2,    -5,    -8,    -7,    -8,    -6,    -4,    -3,    -6,    -8,     1,     8,    16,    10,    -2,    -2,     2,     8,     7,    -2,    -1,    -9,    -4,    -3,    -4,    -4,     7,     1,    -4,    -5,    -9,    -9,    -6,    -9,   -11,    -6,    -7,   -12,     0,    13,    10,    12,     2,     0,    -3,     2,     8,     0,    -8,    -3,     0,     2,    -1,    -7,     0,    -2,     0,    -2,   -11,    -4,    -9,    -7,    -4,    -4,     1,     0,     8,     7,     8,     9,     0,    -1,     0,     3,     2,    -4,    -1,    -3,    -2,    -4,     2,     3,     0,     1,    -6,    -5,    -1,    -3,     5,   -12,    -5,     3,     6,     9,     9,    10,    17,    18,     1,    -3,     2,    -1,     4,     4,    -3,    -3,    -5,    -1,     1,     6,     0,    -3,    -5,    -6,    -3,    -5,     5,    -8,    -2,     5,     7,    10,    11,     6,     5,    -2,     1,     1,     4,     5,    -3,     2,    -1,    -6,    -7,    -6,    -5,    -2,    -5,    -4,    -6,    -4,    -1,     2,    -3,    -5,     3,     6,    11,    10,     5,    -1,     2,    -4,     0,     1,     1,     3,     5,    -4,    -2,    -4,    -2,    -4,    -7,    -4,    -3,    -3,     3,    -5,     4,    -4,    -6,     0,     1,     4,    10,     9,     3,     7,    -8,    -4,     0,     1,     1,     3,     2,     0,    -2,     0,     4,    -5,    -3,     5,     1,     2,     3,     3,     0,    -7,    -9,    -7,     1,     4,    10,    13,     0,     6,    -4,     2,    -1,     2,    -5,    -3,    -5,    -6,    -6,    -1,    -3,    -2,    -7,     0,     5,     0,     6,     0,    -7,    -5,    -5,     0,    -6,    -3,    -7,     5,     3,     2,     1,     0,    -2,     1,    -9,    -2,    -1,    -2,     0,    -2,    -6,    -8,    -9,    -3,    -7,   -14,    -5,    -6,   -10,    -2,    -6,     0,    -7,    -6,    -7,    -5,    -3,    -1,     0,     2,     0,     2,     0,     1,    -4,    -8,    -5,    -6,    -7,   -11,   -10,    -5,    -4,    -7,   -13,   -10,   -20,   -21,   -18,   -15,    -8,    -6,   -10,    -7,     1,    -1,     2,    -2,     1,     1,     1,    -1,     0,     2,    -3,    -4,    -6,    -3,    -6,    -7,    -4,   -11,    -7,    -6,    -7,    -6,    -9,    -3,    -5,    -4,    -6,     2,     0,    -1,    -2,     2),
		    13 => (   -1,    -2,     2,    -1,    -2,     1,    -2,    -2,     2,     1,     2,    -2,    -2,    -3,    -1,     0,     2,     2,    -1,     1,     2,     1,    -1,    -2,     1,    -1,    -1,     1,     1,     1,    -2,     2,     0,    -1,    -2,    -1,     2,     0,    -1,     1,     0,    -1,    -4,    -2,    -5,    -1,     2,    -1,    -2,     0,    -1,     1,    -1,    -2,     2,     1,     1,     1,     0,    -1,     2,    -1,     1,     0,    -6,   -11,     9,     6,    10,    -3,    -4,    -5,    -3,     1,    -1,    -1,    -5,    -3,    -8,    -4,     0,     0,     1,     2,     0,     1,    -1,     1,     1,    -4,     2,    -3,    -6,   -10,   -12,    -8,   -10,   -25,   -35,   -27,   -22,    -3,     3,    -1,    -9,    -8,    -6,   -11,    -1,    -1,     0,    -2,     2,     7,     0,     4,    -9,   -11,    -7,    -5,    11,    -7,     6,    11,    -9,    -6,     0,    -3,    -9,     8,     2,    -9,    -4,     7,    -5,    -5,    -9,    -4,    -3,     0,     2,    -1,    10,     0,    13,    15,     8,     7,    -6,   -10,     0,     0,    -1,    -4,     2,     0,    -5,    -4,    -3,    -2,   -14,   -13,    -6,   -11,    -4,   -11,    -5,    -2,    -1,     0,     2,     4,    11,    12,     4,     0,    -5,     0,    -1,     8,     0,     7,     4,     2,    -1,     6,     1,   -24,    -1,    -8,   -17,    -9,    -4,    -4,    -1,    -2,    -2,     2,     4,    -6,    15,    -6,    14,     4,     2,     7,     1,     5,     1,     5,     5,   -11,    -6,     0,     2,    -6,    -4,     0,   -16,   -11,    -7,    -6,    -8,    -2,    -1,    -2,     4,    -6,    14,     3,     2,     4,     0,    17,     9,     5,    -4,    -1,    -6,     0,    -1,     4,     7,    -5,   -10,     1,    -9,   -24,   -15,    -4,   -10,     2,     2,    -7,     9,     4,    10,     1,    16,    18,     8,     8,    -1,   -15,   -11,    -2,     2,     6,     0,     1,     1,     5,     2,    -4,   -17,   -18,   -19,    -7,    -5,     0,     2,    -9,    10,    15,    13,     8,     9,     5,   -16,   -23,   -31,   -15,   -12,     3,     4,    10,    -2,    15,    -1,     2,     2,    -5,   -13,     0,   -10,    -7,    -6,     1,     2,    -5,     1,    15,     5,    -8,   -15,   -24,   -39,   -20,    -4,    -5,     6,    13,     1,    -1,    -8,    -6,     3,    -1,     4,    -1,   -17,   -13,    -7,    -6,    -2,     0,    -1,    -1,    12,    14,    -9,   -19,   -32,   -19,   -19,     2,    11,     7,    10,     8,     2,    -7,   -12,    -9,   -10,   -20,   -12,   -25,   -13,   -19,    -8,     0,     0,    -3,    -2,     1,    -3,    -4,    -3,   -12,   -19,   -15,    -8,     1,    10,     3,     5,     3,     3,    -9,    -4,    -7,   -11,   -11,   -15,   -16,    -7,    -4,    -4,    -8,    -6,    -4,    -2,     5,     1,     6,     0,    -9,   -11,    -7,    12,    -1,     3,    -1,     2,    -1,     7,    -4,    -4,    -5,   -14,     3,    -9,    -9,   -10,     4,    -1,   -19,    -9,    -5,    -4,     4,     4,    10,    -6,    -8,    -5,    -3,    -2,     6,    10,    18,     0,     2,     3,     5,    -1,   -10,   -11,     0,     1,     9,   -11,    12,    -1,    -9,    -4,    -6,     3,     2,     5,     9,   -11,   -15,    -9,    -6,     4,    13,     0,     1,    10,     9,     7,    -3,     1,    -2,     0,    -7,     2,    14,     6,     7,    -2,   -14,   -14,    -6,     1,     3,     5,    10,   -12,   -22,   -21,   -18,    -8,    -5,   -13,    -2,     2,     6,     1,     1,     6,     1,    -2,     2,    -5,    11,    12,     1,    -7,   -21,   -10,    -4,    -4,    -1,     9,    17,    -4,   -12,   -17,   -23,   -36,   -48,   -40,   -42,   -40,   -30,   -20,   -26,    -7,    16,     2,     5,     5,     4,    18,    10,    -7,   -17,    -9,    -7,     0,    -3,   -15,     9,     8,     9,    -8,    -9,   -15,   -21,   -32,   -35,   -32,   -27,   -22,   -25,   -13,    -6,     2,    11,    10,     8,    12,    13,    -2,   -11,   -14,    -8,     1,     2,   -10,    -6,    -2,     9,     3,    -3,    -1,   -11,   -11,   -10,    -8,    -2,    -3,   -13,   -15,    -2,     0,     8,     7,    -3,     2,    25,    -2,   -11,     1,     1,    -1,     1,     7,     7,     6,    -1,     7,     5,    -1,    -3,     1,    -1,     5,     6,    -5,    -2,    -6,    -1,     5,     3,    12,    -6,    -7,    -2,    -9,   -10,    -3,     1,     2,    -2,    10,    10,    13,     8,     4,     6,    11,     4,    -1,    -5,    -1,     6,    -8,     1,    -1,    -8,     3,     2,     5,     4,    -1,     5,   -17,   -12,     0,    -2,    -1,     1,    11,    14,    13,    -1,     1,     5,     4,     3,    -2,     6,    -5,     5,    -5,    -3,    -5,    -5,   -13,     0,   -10,    -4,   -10,    -1,   -11,    -2,     2,     2,     2,     2,     3,    -2,    15,    10,     4,    14,    10,     0,    11,     8,     4,    -2,     3,    -5,    -6,     2,    -3,    -9,   -16,     1,     7,     2,   -10,     1,     0,     0,     2,     1,    -2,    -9,     3,    12,     3,     6,     9,     5,    -2,    -6,    -8,   -11,   -14,    -9,    -3,   -15,   -16,   -16,   -11,    -9,    -5,   -28,   -12,    -2,    -2,     0,     2,     0,     2,    -6,     1,     1,    -8,    -4,   -11,   -13,   -15,   -15,   -13,     5,    -5,   -10,    11,    -1,     3,    -2,    -2,     1,    -8,    -1,    -1,    -2,     1,     0,     2,    -2,    -1,    -1,    -3,     2,    -2,     2,    -1,   -12,    -9,    -7,     1,    -8,    -5,    -6,    -3,    -1,    -4,    -9,   -10,    -2,    -4,    -2,    -1,    -2,    -2,     1),
		    14 => (    0,    -2,     2,    -2,     1,     2,     1,    -2,     0,    -1,     0,     0,    -7,    -4,     0,    -1,     1,    -2,    -1,    -2,     2,     0,    -1,     2,     2,     1,     2,     2,     1,    -1,     2,     2,     1,     0,     0,    -5,    -2,    -3,    -8,    -7,    -9,    -6,    -2,   -21,   -17,   -13,    -4,    -3,    -8,    -4,    -2,    -2,    -1,    -1,     0,     2,     2,    -2,    -1,    -7,   -21,     0,    -2,    -7,   -12,    -9,   -17,   -17,   -17,     0,     4,     4,   -16,   -11,    -6,    -5,   -16,    -8,     1,    -1,    -2,   -11,     0,    -2,    -1,     0,     0,    -7,   -21,   -16,    -7,    -3,    -4,    -6,   -15,   -16,   -11,     1,     6,     1,   -12,   -15,     0,     8,    11,     9,    -4,   -11,   -17,    -9,     1,     0,     2,    -1,    -3,   -14,    -6,    -8,    -4,     3,     6,     9,    -1,   -16,   -17,     1,     2,    -3,    -4,    -5,     6,    -2,     9,     2,    -1,    -8,   -16,   -10,   -12,    -2,     0,     2,    -6,    -2,    -5,     0,     6,     4,    10,     5,    -2,   -14,   -14,    -9,    -1,    -6,   -11,     2,     3,     7,    -1,    -2,     0,    -1,    -5,     6,   -13,    -3,    -1,     0,   -10,    -4,     7,     7,     2,     3,     0,    -6,     1,    -5,     6,     5,    12,    24,    24,    18,    11,    10,     2,    11,    -6,    -2,    -3,    -7,     1,    -5,    -1,   -18,    -5,     3,     4,     5,    11,    11,     1,     4,     5,    -1,     6,     7,     6,    16,    18,    14,     2,    -3,     0,     0,     1,     1,    -5,     3,    -2,   -18,    -8,   -21,    -2,     1,     1,     2,    13,     8,    11,    -2,   -10,    -2,    -5,    -1,    -4,     2,     1,    -4,     0,     0,    -2,     2,    -2,    -1,     3,     7,    -1,   -16,    -1,    -9,   -11,     1,     0,     3,    -1,    -1,    -2,   -16,   -16,    -3,    -9,   -14,   -17,    -8,    -6,    -7,    -1,    -7,     1,     7,     2,     2,    -6,    -3,    -6,   -12,     1,    -8,     2,     0,    -5,    -4,    -8,    -6,    -9,    -9,    -6,    -6,    -8,   -20,   -23,   -15,   -12,    -8,     2,    -4,    -9,     9,    -3,   -16,   -19,   -12,    -7,    -4,    -1,    -7,    -6,     0,    -9,     0,    -8,    -4,    -9,    -9,    -8,   -10,     0,    -8,   -18,    -2,    -7,     3,     3,     5,    -4,     5,    -8,   -23,   -22,   -15,   -10,   -15,    -1,     1,     2,     4,    -5,     3,     6,    -1,     5,     5,     6,     2,     9,     7,   -11,     5,     4,    -1,    -1,     4,     6,    18,     4,    -5,   -13,    -8,   -18,   -19,    -1,    -3,    -8,    -1,    10,    -2,     0,    -2,     6,     4,     1,     8,     5,    -3,     3,    14,     7,     8,     9,    10,     7,     4,    -4,    -4,   -14,    -6,   -13,    -1,    -2,    -4,   -21,    -4,     9,    -3,    -2,    -1,    -2,     0,    -7,    -3,    -9,    -4,     2,    13,     4,     9,    13,     9,    10,     3,     1,    -6,     1,    -8,    12,     2,     1,     0,    10,     3,     7,   -13,    -6,     0,    -3,    -9,   -20,   -12,    -7,     6,    11,    19,    17,    15,    15,    -2,     1,     3,     4,    -4,   -10,   -11,    13,   -10,     1,     0,     2,     6,     7,    -9,   -10,    -5,    -7,   -12,   -16,    -2,     3,    14,    21,    17,    20,     5,    13,    -5,     1,    -2,    -4,    -6,    -5,     2,     1,    -4,     2,    -1,     5,    -4,    15,   -12,    -5,    -6,    -1,   -11,    -3,     6,    15,    14,    13,    14,    20,     6,    10,    -8,    -4,    -2,     2,     1,    -8,     1,     9,   -11,   -13,    -2,    -1,    -2,    12,    -8,    -5,    -7,   -22,    -5,     3,     5,    11,     2,    13,    12,    14,     5,    -1,   -10,     2,     1,    -2,    14,   -12,   -15,    -4,    -2,     0,    -3,    -8,    10,    -1,    -2,     1,     1,    -2,     5,     6,    17,     0,    -8,     7,     7,    -1,    -7,     8,     3,    -4,     2,    -1,    -1,    -9,    -7,    -5,    -2,     2,     1,    -4,    -8,   -14,   -12,    -9,     1,    10,     8,    10,    10,     9,     9,    -2,     4,    14,     1,    10,     5,     8,     3,     2,    -1,   -12,   -18,   -10,     0,    -2,    -3,   -13,    -6,   -16,    -2,   -18,    -1,     5,     3,     1,    -6,   -13,   -12,    13,     9,     5,     4,    -2,     5,     4,    -4,     6,     3,    -4,   -27,   -16,     1,    -3,    -4,    -3,   -11,   -33,   -15,    -3,    -2,     2,   -16,     1,    -5,    -7,    -4,    -3,     7,    -1,   -10,    -5,     4,    -3,     5,     0,     6,    -8,   -14,    -6,    -4,     1,     0,     0,   -18,   -28,   -25,     7,    -1,   -11,   -11,    -5,    -8,    -9,    -4,     4,    -4,    -5,    -5,     3,     9,     2,    -5,    -9,    -1,    -6,    -2,    -3,    -1,     2,     0,    -3,    -4,   -20,     3,    -1,    -7,   -13,   -11,   -12,    -7,    -6,     2,    -2,    -7,     1,    -6,     0,    13,    -8,   -11,    -3,     3,   -13,     7,    -9,     1,     0,     2,    -1,    -1,    13,     9,   -12,   -14,   -11,    -1,   -12,     3,    -1,     7,     3,     3,    -2,    -9,    -6,    -3,   -12,   -15,    -5,     6,    -3,   -10,   -10,    -2,    -2,     1,     2,   -10,    14,     1,    -8,   -19,   -11,   -10,   -13,    -8,   -22,   -17,   -19,   -20,   -14,   -19,   -15,    -7,   -21,   -32,   -34,     1,    -1,    -1,    -2,     0,     1,     1,    -1,     1,    -2,    -4,    -5,    -9,   -10,    -9,   -17,   -14,   -10,   -11,   -20,    -2,   -11,   -14,    -9,   -12,   -14,   -11,   -13,    -1,    -2,    -1,     1,     1),
		    15 => (   -1,    -2,     0,     2,    -2,    -1,     1,    -2,     2,     2,    -1,     0,     1,     0,    -1,    -1,     2,     2,    -1,    -1,    -2,    -1,     2,     0,     1,    -2,     0,    -1,    -2,     0,    -1,     0,     2,     2,    -2,     1,     2,     0,    -2,    -3,    -5,    -6,    -5,    -4,    -5,   -10,    -5,    -4,    -4,    -2,     1,     1,     0,    -2,     0,    -2,    -2,    -2,    -2,    -3,    -1,     2,    -3,    -7,    -6,   -14,    -6,    -2,    -6,   -11,   -13,   -17,    -7,    -4,     1,     0,    -3,    -8,    -2,     1,    -4,    -3,    -2,    -1,     1,    -1,    -5,     5,     2,    -5,     0,   -11,   -11,   -11,   -11,    -6,    -5,   -11,   -12,   -18,   -21,   -12,    -5,    -2,    -2,     4,     3,    -2,    -5,    -6,     1,    -2,    -2,     1,    -3,     3,    -3,    -2,    -1,     4,    -5,     3,   -11,    -9,   -14,   -15,    -3,     4,   -11,    -5,    -6,    -4,   -10,    -2,    -6,     4,     5,    -6,   -11,   -11,     1,    -2,    -3,     0,    -2,     3,     6,     5,   -10,    -9,     2,    -2,    -7,   -13,     2,     4,    -3,    -8,    -7,    -6,     2,    -3,   -11,   -16,   -12,    -3,    -5,    -8,     1,    -3,    -1,    -6,    -5,     6,     5,    -2,    -7,    -8,    -6,     2,    -5,    -1,     9,    -7,   -10,   -14,   -11,    -1,    -2,    -5,    -1,    -2,    -7,    -1,    -1,     8,     2,    -3,    -3,    -9,    -2,     2,     2,    -6,    -8,   -13,     2,     1,    -5,    -9,     3,    -8,   -13,   -13,   -25,   -23,   -20,    -8,    -1,    -3,     4,     3,     3,     6,    -1,   -11,   -10,   -11,    -8,     9,     0,    -3,   -16,    -5,     6,    -8,    -3,     1,   -10,   -20,   -11,    -9,   -20,   -19,   -10,    -8,    -8,    -2,     1,    -8,   -19,     0,     0,    -2,    -4,   -10,    -6,     8,    -8,   -15,    -5,    -1,     4,     0,     1,   -17,    -4,   -15,     4,     4,     5,    -5,    -7,    -1,    -4,     2,    12,     4,    -4,    -3,    -2,    -4,    -1,    -2,    -9,    -4,    -1,   -12,    -2,    -1,     5,     1,    -4,     8,    -3,     3,    12,    12,    13,    13,    11,     6,     7,    22,    14,    18,     4,    -4,     1,    -2,    -3,    -3,    -5,    -6,     6,    -6,    -1,     2,     5,    11,     1,    -3,    -3,    -3,    10,     1,     7,     9,    15,    18,    20,    22,     6,    10,     1,     0,    -2,    -1,    -1,    -8,   -13,    -5,    -1,    -4,    -1,    11,    10,     2,     3,     0,     6,     1,    -4,    -2,     0,     3,    18,     9,    15,    11,     2,    10,    20,    -3,    -1,    -1,    -2,    -4,   -16,    -3,    -9,    -7,     4,     3,     9,     2,     2,    -2,    -6,   -17,    -4,    -2,   -25,   -15,   -10,   -13,    -2,    -5,    -2,     1,    18,    -6,     0,    -1,    -5,   -12,     8,     6,    -2,    -1,    11,     4,     5,    12,     5,     7,   -16,   -17,   -14,   -13,    -8,   -18,    -6,    -9,    -4,    -9,   -11,   -12,    -6,     1,     3,     2,    -4,    -7,    17,    -1,     3,    -2,    -3,     7,    -2,     3,    12,    -1,   -12,    -9,   -16,   -16,    -5,   -11,    -8,    -5,    -7,   -12,    -1,   -18,    -4,    -5,    -3,    -4,    -4,    -1,   -15,   -10,   -16,    -6,   -12,    -7,    -4,    -4,     1,     0,    -4,    -2,    -1,    -1,    -2,   -10,   -13,    -3,   -13,    -3,    -6,   -16,    -8,    -6,    -2,    -3,    -4,    -6,    -9,   -13,   -14,   -21,   -18,    -3,   -15,     0,    -4,   -12,     1,    -1,    -5,    -1,    -1,    -5,    -1,    -4,   -16,     8,   -11,   -19,   -10,   -17,    -2,     0,    -4,     2,    -1,    -2,     0,    -4,   -13,    -7,    -6,     5,     4,    -7,   -11,   -14,     8,     4,     1,    -8,    -2,    -7,    -8,     5,    -7,    -4,   -11,    -9,    -1,    -2,     5,   -11,    -2,   -11,     7,     6,    -8,    -5,    -1,     2,    -4,     0,     5,     2,    10,     2,     6,     1,    -4,   -10,     3,     9,    -4,   -12,   -11,   -10,    -1,    -6,     4,   -10,    -8,    -6,     6,    10,    -2,     4,     9,    -6,    -2,     3,    -7,     1,     8,     7,    -3,    -3,    -8,     3,     8,     2,    -3,    -1,   -15,     2,     0,    -2,    -2,    -1,    -8,     4,    10,    11,     2,     0,     3,    -7,   -11,     4,    -9,     4,     3,    -1,     8,     1,     7,     5,    -1,    -1,   -12,    -2,   -11,    -2,     0,     2,    -2,     6,    -1,    -3,     4,    -3,     5,     1,     6,     5,    11,     4,     6,     6,     1,     4,     0,     4,     7,     2,    -4,    -2,   -10,    -1,    -4,    -1,     0,     1,     5,    -4,    -9,   -12,    -4,    -2,     9,     4,     4,     2,     7,    13,     8,    -5,    -2,     2,    -8,     4,     6,    -4,    -8,     1,    -1,     1,    -2,     0,    -2,    -2,    -5,    -1,    -1,   -11,   -11,   -10,     9,    10,     7,     3,     2,    -3,     8,     3,     3,     8,    -4,     3,     1,   -11,    -5,     3,    -1,   -11,    -3,     2,     0,    -2,    -2,     2,    -6,   -15,    -8,   -18,   -11,   -17,   -11,    -8,   -11,   -14,   -10,    -6,   -12,   -17,   -11,    -8,    -4,    -3,    -4,    -2,    -1,    -1,     2,    -2,     0,     2,    -2,    -3,    -2,   -11,   -14,   -13,     0,    -6,     3,    -4,   -10,   -18,   -17,   -17,   -14,    -8,   -11,    -2,    -3,     2,     0,    -6,     0,     2,     1,    -2,     2,    -1,    -1,    -2,    -4,     0,    -2,    -3,     0,     1,     1,    -1,    -3,    -3,   -15,    -7,    -5,    -1,    -1,    -6,    -7,   -10,   -10,    -3,    -2,    -1,     0,    -2),
		    16 => (    1,    -2,     2,     0,     2,    -1,    -1,     0,     3,     0,     0,    -1,     4,     1,    -2,     0,    -1,    -1,     2,     2,     0,     0,     0,    -2,    -1,    -1,     2,    -2,     0,     1,     1,    -2,     1,    -2,     1,     7,     2,     2,     2,     3,     9,     4,    -7,     1,     4,     4,     2,     1,    11,     2,     3,     2,     2,     1,     0,     2,    -1,    -1,     4,     1,     3,     3,     5,     6,     5,    -3,    -4,    -1,    -9,    -7,     4,     3,    15,    17,     2,    -9,   -12,     6,    10,     7,     3,    -3,     0,     0,    -2,     0,    -3,     0,     4,     7,    -2,    -1,     0,    -5,    -4,    -2,   -11,    -3,     7,     9,    16,     7,    -3,     3,    14,     7,    -6,    -2,     1,     0,    -1,    -2,     2,     1,    -7,    -7,    12,    11,    -2,    -3,    -6,    -4,    -4,   -10,   -11,    -5,   -10,     1,    -2,     1,    -7,    -3,     1,   -10,     1,    -9,    -8,    -4,     6,     6,     2,    -1,    -5,    -1,    14,    12,     1,    -1,    -3,    -1,   -13,   -21,    -7,   -13,    -3,    -4,     6,     6,    -4,    -3,   -16,   -13,    -1,    -9,    -2,     0,     5,     2,     1,     0,     1,    -7,     8,     7,    -1,     0,    -3,    -6,   -18,   -20,   -12,    -2,     3,    11,     1,   -11,     6,     5,    -2,   -16,    -3,    -3,     1,    -1,    -2,     3,     2,    -1,     0,   -12,     6,     8,    -1,    -6,    -5,    -8,   -15,   -19,   -11,     1,     2,   -15,    -9,   -15,    -9,     1,     1,     6,     7,     1,    -2,     3,     1,    -4,    -1,     1,    -2,   -12,     7,     8,     2,    -1,    -8,    -9,   -14,   -21,    -5,     2,     2,   -10,    -5,    -9,   -14,   -10,    -4,    11,     4,    -4,    -3,    -1,    -8,   -12,     1,     0,    -1,    -6,    12,     9,     1,     3,    -4,   -10,   -11,    -3,     4,     5,    -2,     2,   -10,    -7,   -12,   -10,   -10,    -9,    -9,     1,    -2,     1,     0,    -3,     2,    -2,    -4,    -7,    11,    12,    -3,    -4,    -7,    -3,    -2,    -8,     5,     0,    -1,   -16,   -10,   -11,   -21,   -15,   -12,   -14,    -7,     1,     2,     1,    -4,    -2,    -1,     2,     0,    -9,    14,    13,    -2,    -4,    -7,   -11,    -9,     3,    -1,    -5,    -8,   -11,    -7,   -14,   -19,   -15,   -10,   -16,   -12,     3,     4,     1,    -3,    -6,     1,     0,    -2,    -7,     8,    11,    -4,    -8,    -8,    -4,    -1,    11,     3,    -6,    -5,     0,   -11,   -17,   -12,    -7,    -5,   -14,   -12,     7,     6,     0,    -7,    -5,     1,     1,     2,    -6,     9,     8,    -1,    -5,    -4,    -6,    -1,     5,    -1,    -1,     3,     4,    11,     3,    -6,    -6,    -3,   -10,    -9,     4,    -7,    -9,    -7,     0,     2,     2,    -2,    -2,     0,     7,     5,     1,    -2,   -13,     0,    -1,    -1,    -4,    -7,    -2,     9,    -7,   -11,     0,     6,    -8,    -9,    -2,    -4,    -4,    -5,    -3,     2,     0,    -3,    -7,    -2,     2,     3,     0,    -5,    -9,    -1,     1,    -1,   -17,    -3,    -3,     3,    11,     0,    12,     9,    -7,    -2,    -4,    -7,    -7,    -3,    -9,    -1,     2,    -2,    -8,    -3,     3,    -1,     5,     4,   -10,    -1,    13,    11,   -10,    -3,   -12,    -2,     3,    -7,     6,    -1,   -10,    -5,    -8,    -4,    -2,    -5,    -4,     1,     2,     1,    -9,    -5,    -3,     2,     3,     4,   -10,     7,    16,     4,   -18,   -16,    -6,     2,    -7,    -1,     5,    -1,    -9,    -7,    -4,    -7,   -13,    -2,    -7,     2,     0,     0,     2,    -6,     0,     0,     0,   -11,    -9,     0,     2,     7,     1,   -13,   -10,     0,     5,     4,     4,   -13,    -8,   -12,   -10,   -12,   -13,    -2,    -7,     1,    -1,     1,     0,    -3,    -6,    -7,    -8,    -8,   -12,    -1,    13,     7,     8,     0,    -4,    -8,     6,     3,     3,    -8,    -5,   -10,    -9,    -9,    -7,    -7,    -3,     1,    -2,    -2,    -2,     0,    -4,    -6,   -10,   -11,   -16,   -14,    -1,     4,     9,    -2,     1,    -3,     9,    -1,     5,     3,    -5,    -4,    -5,    -4,    -4,    -1,     0,    -1,     0,     1,    -1,     2,    -2,    -3,    -7,    -9,   -14,   -13,   -13,     0,     6,     1,    -2,    -5,    -2,     0,    -1,   -11,    -6,    -4,    -3,    -5,    -7,     0,     1,     2,     0,     0,    -3,     1,    -2,     2,     0,    -7,   -16,     2,    -5,     0,     2,     8,     8,    -5,   -12,   -13,     4,    -3,    -4,     1,    -3,   -10,    -3,     2,     1,     1,    -2,    -1,    -3,     1,    -1,     0,    -3,    -3,   -10,   -12,    -7,     2,    -3,     1,    -3,    -4,    -5,    -1,     1,    -5,    -4,     1,    -1,    -1,    -3,     2,     1,     2,     1,     0,    -3,    -3,    -4,    -3,     0,    -6,    -3,    -7,     2,     3,     4,     0,    11,    19,     8,   -13,   -19,    -5,    -1,     0,    -1,    -2,    -3,     0,     1,     1,    -2,     0,    -2,     2,    -3,    -2,    -2,     0,    -4,    -2,     1,     5,     4,    -2,    -1,    -3,    -1,    -2,    -3,    -6,    -1,    -3,    -4,     1,     2,     1,     0,     0,     1,     1,     1,    -1,    -1,     2,     1,     1,     0,    -2,    -3,    -1,     1,     2,    -3,     0,     0,     1,    -2,    -1,    -4,     1,     0,     2,     2,    -2,     1,    -1,    -1,     2,     2,     0,     0,    -2,    -1,     1,    -2,    -1,     1,     0,     1,     1,    -3,    -2,     0,     2,    -1,     1,     1,     1,    -2,     2,     0,     0,     0),
		    17 => (   -1,     1,    -2,     1,     0,    -1,    -2,    -2,     2,     1,    -2,     2,     1,     2,     2,    -2,     0,    -2,     2,    -1,    -2,     1,    -1,     2,    -1,     0,     1,     1,    -1,     0,     2,     0,     2,     2,     1,    -1,    -1,     1,    -2,   -10,    -9,    -6,    -2,    -8,    -8,    -6,     1,     1,     2,     1,     0,    -2,     2,     1,     1,     0,    -1,     1,     1,    -5,    -4,     1,    -2,     0,    -4,    -3,    -2,    -8,    -4,    -4,     0,    -6,    -6,    -1,    -1,     2,    -1,     1,    -2,     0,     2,     1,     2,    -1,     1,     0,     1,    -9,    -2,    -3,    -3,    -7,    -9,    -7,    -5,    -4,    -5,    -7,    -4,    -7,    -2,    -2,    -4,    -3,    -3,    -4,   -12,    -5,    -1,    -3,     2,    -2,     1,    -1,    -2,    -1,   -12,    -5,    -2,   -16,   -15,    -8,   -16,   -25,   -22,   -20,   -15,    -8,    -5,    -1,     1,    -2,   -10,   -12,    -7,   -13,    -3,    -5,    -3,     1,     2,     3,    -1,    -2,   -12,    -6,    -4,     4,     3,    -2,   -10,    -6,     2,     1,   -14,   -17,   -18,   -34,   -39,   -36,   -35,   -20,    -2,   -12,    -8,    -6,    -3,    -1,    -2,     2,    12,    13,    -1,    -2,     0,    -6,    -6,   -11,   -16,     6,     9,     5,    -6,   -20,   -15,     0,    -2,    -2,    -5,    12,     7,     3,    -9,   -10,   -16,    -5,    -2,    23,    21,    14,     2,    -2,     0,    10,    -3,     0,     2,    -6,     5,    -2,    -7,   -10,   -10,    -3,    -1,    -4,    -8,     1,    -3,     6,     5,    -1,   -12,    -6,   -15,    25,     8,     2,    -5,    -8,    -6,    -2,   -11,    -1,    10,     1,     4,    -9,    -7,    -5,    -7,     5,     6,     1,    -3,    -9,    -4,    10,    16,     4,    -9,    -8,     1,    14,   -11,    -1,     4,     1,     6,    -2,    -6,     2,     2,     5,     3,     1,    11,    -1,    -7,     4,     8,     7,     1,     2,     2,     6,    17,    -2,   -16,     0,     2,    11,     8,     2,     4,     2,    10,     4,     5,    -1,     1,     9,     9,    13,    -1,   -10,    -8,     3,     0,     7,    10,     9,    -7,    -5,    -7,    -6,   -13,     4,    -1,     2,     9,    12,     4,    14,     3,    -6,   -10,    10,     4,    17,    19,    -1,   -16,   -10,    -6,    -2,    14,     7,    10,    -3,    -9,     0,    -4,   -11,    -6,     2,     3,     3,     5,     8,     1,     7,     3,    10,     7,     5,    11,     6,    12,   -31,   -33,    -5,     5,     5,     7,     0,     4,    -4,   -10,   -10,    -6,    -8,    -1,     7,     0,     4,    11,    -3,    -2,    12,     8,    11,     9,    -1,     1,     1,    -7,   -42,   -28,   -15,     7,    -1,     8,    -7,     0,     5,    -9,   -17,    -1,   -13,    -4,    -2,    -3,     8,    22,     8,    -6,    13,     4,    -3,    -2,     9,    13,     3,   -20,   -55,   -25,    -9,     5,    -2,    11,     6,    -2,    -2,    -2,    -2,     1,    -8,    -6,    -1,    -2,     0,     6,     8,   -20,     5,     7,     7,    -9,    -5,    14,    -7,   -48,   -34,   -18,    -8,     7,     6,     4,    10,     0,    -4,     1,    -8,   -11,   -11,    -1,    -4,    -3,    -3,     3,     3,   -10,    -7,     2,    14,    -2,    -1,    15,   -20,   -47,    -6,     1,    -3,    -3,     2,     9,     8,   -10,    -1,     6,    -6,    -6,   -10,    -1,    -9,    -2,     1,     7,    -4,     2,    -7,     2,    -1,    -8,   -16,   -23,   -32,   -25,    -2,     3,    -2,    -3,    -5,     8,    -7,     2,    -1,     8,   -24,   -31,    -5,     0,   -11,     6,    -2,    13,   -20,    -8,    -2,     5,     1,   -12,   -24,   -40,   -11,    -3,     6,    11,    -2,     4,     6,     6,    -7,     8,    -6,    -9,   -30,   -28,     3,     0,    -4,    -2,     7,     5,   -16,    -3,     3,     4,   -25,   -25,   -29,   -31,   -10,    -1,     0,     3,     0,    -3,    -6,     5,     0,    -5,   -12,   -19,   -22,   -14,    10,     0,    -2,     0,     9,    -1,   -10,    -6,    -5,   -10,   -24,   -24,   -32,    -7,    12,     8,    -6,     0,    -8,    -5,     2,    -7,    -2,    -8,   -19,   -16,   -23,    -9,     0,    -1,    -1,    -1,     0,    -4,   -12,   -23,    -6,   -21,   -20,   -18,    -7,    16,     5,    -5,    -8,    -5,   -14,    -8,    -1,     7,     2,    -1,    -4,    -1,    -3,    31,     2,    -2,     1,     0,     2,    -2,    -6,   -15,     2,     1,     0,     2,     5,     1,     3,    -6,     0,     1,     0,    -3,     1,     3,     6,     2,    -5,     0,    -4,    -2,     0,    -6,    -1,     1,     1,    -2,   -15,    -8,     9,    11,     7,     8,    -1,     4,   -16,     1,     5,     0,     0,    -6,    -5,     5,   -10,    -5,    -2,   -21,   -14,    -2,    -5,    -2,    -2,    -2,     0,     4,     4,    -1,    10,    -4,   -12,     7,    -1,     2,     4,     3,     0,     7,    -4,    -7,    -5,   -15,   -10,    -5,     3,   -17,   -17,    -4,   -14,     2,     1,     2,     0,    -2,    -1,   -18,   -22,    -8,    -6,     0,    -2,     4,     3,     5,     1,     8,     0,     5,     7,   -10,    -3,    -4,     4,    -1,   -11,     5,    -3,    -2,     1,     1,     1,     2,    -1,   -19,   -18,   -15,   -16,    -7,   -10,    -9,   -12,     2,    10,    10,     1,     7,    -3,     0,     5,    -4,    -5,    -3,     0,    -5,     2,     0,     1,     2,     2,     1,    -1,     6,     6,     2,     5,    10,     3,     5,     3,    -3,    -2,     3,    -5,    -6,    12,    11,    -9,     5,    18,     4,     9,    -1,     2,     0,     0),
		    18 => (    2,    -2,     0,     0,     2,     0,     0,    -2,     0,    -1,    -2,    -1,    -1,     2,    -1,     1,     1,     1,    -1,    -2,     1,     2,    -2,    -2,     0,     1,    -2,     1,     2,    -2,    -1,    -1,    -2,     2,    -2,    -1,     2,    -2,     1,     1,    -2,    -4,    -6,   -11,   -17,    -8,    -3,    -4,    -3,    -5,    -5,     0,     2,     2,    -1,     0,     2,    -1,    -3,     0,     0,    -1,    -7,    -4,    -5,   -15,   -18,   -10,    -3,     1,    -3,   -12,    -8,    -3,     4,    -6,   -19,   -16,   -18,    -5,    -4,    -3,     2,     1,    -1,     1,    -7,    -8,     0,    -6,    -9,   -20,     4,     2,    -2,    -9,   -10,   -14,   -21,    -1,     3,     2,     7,     4,    18,    15,     7,     6,    -7,    -2,    -5,     0,     0,     2,    -1,   -12,   -11,   -19,     0,     0,    -8,   -13,     2,    -6,   -17,   -14,     7,     1,     3,    -2,    -2,     6,    13,    15,     8,     5,     0,    18,     8,    -3,    -2,     1,    -9,   -13,   -19,    -6,    -1,     1,     5,    -2,    -1,     0,    -7,    -7,    -6,     2,     0,    -8,   -10,    -4,    13,     7,     3,    16,    17,     7,    -7,    -1,     1,     1,    -7,   -12,    -3,   -10,     3,     5,     5,    -1,    -4,    -7,     4,     0,     3,     0,   -12,   -12,    -4,     7,     1,    -6,   -12,     4,    -1,    20,     1,   -10,    -1,   -14,    -8,    -2,     0,   -12,     5,    13,    -1,    -7,    -5,    -3,     1,     0,     2,     5,   -12,    -3,     8,     3,    -6,     1,     6,     6,     4,    -2,    -2,   -11,    -4,    -4,    -7,     4,    13,    -5,    10,    10,    -9,     5,    -3,     2,     2,    11,    -5,   -16,    -7,    -5,    -6,   -13,     1,    12,     7,    -1,     2,     8,     7,     4,    -1,     2,    -2,     8,     4,   -12,    -5,    -3,    -6,    -4,     4,    10,    -3,    -4,   -12,   -17,    -1,    -2,    -9,     5,     5,     4,     2,    10,     2,     3,   -12,   -27,     1,    -3,    -4,    -8,    -1,   -12,    -8,   -14,     3,     7,    10,     2,    -2,   -10,   -10,   -10,     2,    10,    -4,    -5,    -3,    -4,     0,     7,     0,   -19,   -10,   -21,    -1,    -2,    -7,   -10,   -10,    -7,    -4,     1,    -6,     7,     0,    12,    10,    -2,    -4,    -7,     0,    -6,    -4,   -17,    -9,   -20,    -9,     9,    18,     2,    16,   -12,     0,     1,   -12,    13,    -7,    12,     1,     3,   -12,    -5,     0,    -8,     5,     9,    -2,    -7,    -8,     0,     3,     8,   -12,    -3,    11,    21,    20,     6,     5,   -22,     0,    -1,   -11,    11,    -3,    -7,   -21,    -8,    -9,   -10,    -2,    -2,     2,     6,     1,    -2,   -14,     3,    -1,     5,     7,    17,    25,    21,    11,    -6,    -7,     3,    -4,     0,     0,   -18,     0,   -17,    -8,    -8,   -14,   -18,     0,    -8,     0,    11,     3,     2,   -12,     9,   -11,     5,     0,    11,     2,    17,    11,    -6,   -15,     0,     0,     1,    -3,     7,    -2,     4,     1,    -5,     0,   -16,    -4,     2,     6,     3,    -1,    -5,     7,   -21,    -7,     3,    -8,   -16,    -4,    13,    13,     0,   -18,   -12,    -1,    -2,    -5,     9,   -13,    12,    -3,     3,   -10,   -12,    -6,    -1,    10,     2,    -1,     3,   -10,    -5,    -4,   -14,   -18,   -13,    -9,     6,     2,     5,   -13,   -10,     0,    -2,    -6,     5,   -19,    -3,    -2,     8,    -6,    -9,     1,     8,     9,    -6,    10,     9,    -3,    -3,   -18,   -15,    -8,   -13,    -8,     0,    -2,     2,    -3,    -7,    -4,    -2,    -2,    -7,   -13,    -6,    -4,    -8,   -10,    10,     7,    14,    -7,   -22,    -4,    11,     0,    -3,    -5,     6,    -4,   -22,    -6,     1,   -14,     2,    -1,    -7,     1,    -2,    -5,    -5,   -15,    -6,    -6,   -13,    11,     4,    12,    11,   -10,   -21,    -9,     4,     2,     8,   -10,    -2,    -7,   -13,    -1,    -9,    -9,     0,    -9,    -3,     0,     2,    -3,    -7,   -22,    -2,   -11,     7,     5,     5,    10,    13,     2,    -6,    -2,     2,     0,    -5,     0,     1,    -7,    -7,    -7,    -9,     0,     3,   -10,     1,    -2,    -7,    -6,    -1,   -19,   -23,     2,     4,     4,     4,     1,    -1,     4,   -10,    -8,     5,   -11,    -6,     3,    -6,   -22,   -12,    -2,    -8,    -4,     6,   -12,     0,    -3,    -2,    -3,    -9,   -13,   -28,   -13,     3,    -3,     1,     0,     6,    -3,     6,    -7,    -2,   -20,     0,     2,   -19,   -29,   -13,    -8,    -8,     1,     6,   -17,     0,     0,     1,    -7,   -12,   -16,   -19,    -7,     1,    11,    -7,   -12,     1,     6,     3,     4,    -9,    -3,    12,   -13,   -29,   -26,   -12,   -13,    -4,     6,     5,   -17,     1,    -1,    -1,    -2,    -1,   -17,   -23,   -13,    -1,     6,     1,    -2,     3,    10,    10,     5,    -2,     5,   -10,   -14,   -17,    -8,    -6,    -8,    -3,    -6,   -14,   -13,     0,     0,    -1,    -8,    -5,    -8,   -12,    -5,    -2,   -10,   -10,    10,   -12,   -14,    -6,    -3,     7,    -5,     0,     4,     8,     8,    -3,    -9,    -4,   -11,    -6,    -6,    -1,    -1,     0,     2,    -2,    -3,    -9,   -13,    -1,     1,    -7,   -18,   -13,   -10,   -14,   -20,   -19,    -8,    -4,    -1,    -4,    -7,    -8,    -7,    -2,    -1,     1,     2,     1,    -1,     0,    -2,     2,    -4,    -2,    -1,    -6,    -8,    -4,    -4,    -4,    -1,    -5,    -4,     1,    -2,    -2,     0,    -1,    -2,    -2,    -2,     1,     0,    -2,     2,     0),
		    19 => (   -1,     1,    -1,    -1,     0,     1,     0,    -2,     1,     2,    -1,    -1,    -1,    -1,     2,     0,     2,     2,     0,     0,     1,     1,     0,    -1,    -2,     0,    -2,     2,     1,     2,    -2,    -1,     2,     0,     2,    -2,    -3,    -2,     0,     3,    -3,    -3,     0,    -6,    -5,    -8,    -3,    -2,     1,    -3,     0,     0,     2,     2,    -2,     0,    -2,     2,     2,    -1,     0,    -1,    -1,    -1,     0,    -3,    -2,    -2,     1,    -1,    -6,    -3,     0,    -2,    -5,    -1,    -4,     1,    -1,    -2,    -2,    -2,    -1,     2,     0,     1,    -2,     0,    -3,   -11,    -1,    -1,    -8,    -1,    -1,     0,    -1,     0,    -7,   -16,    -8,     3,    17,     6,   -10,    -5,    -6,     0,    -1,    -3,    -2,     2,    -2,    -1,    -2,    -3,     0,    -6,    -6,     0,    -3,     1,     2,    -2,    -8,   -11,   -15,   -23,   -26,   -26,   -16,   -19,   -23,   -12,   -11,   -14,    -9,   -13,    -7,    -1,     1,     1,    -5,    -1,    -2,    -1,    -3,    -1,   -11,    -1,    -4,    -9,   -22,   -25,   -32,   -32,   -25,   -22,    -7,    -6,     1,    -3,   -10,   -18,   -13,   -10,   -12,     1,    -1,    -4,    -8,    -8,     5,    -1,    -6,    -7,    -8,   -17,   -13,   -30,   -33,   -18,    -1,    -4,    -1,    10,     8,    -8,    -3,    -5,   -11,   -16,    -9,    -8,   -10,   -11,     1,    -7,    -9,    -4,    -5,    -4,    -7,   -10,    -4,   -24,   -33,   -20,    -6,     5,     5,    14,    13,    -6,     7,    -1,    10,    -7,    -5,     4,   -14,   -10,    -8,    -6,   -10,    -7,    -8,     2,    -2,     0,    16,    -7,    -1,   -11,   -13,    -7,     4,     6,    -5,    -9,    -1,     2,     4,     8,   -14,     1,    12,     9,   -16,   -16,    -9,    -3,    -1,    -8,     8,     7,     9,     2,    -3,    -7,   -19,    -6,     3,     6,     7,     0,   -13,     0,   -14,   -24,    -8,     0,    -8,    -7,    19,    -7,    -8,   -17,    -3,    -7,     1,   -11,   -19,     9,    10,     3,    -9,   -16,    -7,     5,     5,    10,     3,     2,     1,    -1,   -11,   -13,     0,     0,    -4,     1,     0,    -9,    -3,   -14,   -11,    -6,     0,    -5,    -8,     2,    -2,    -2,    -5,    -1,    -6,    -5,    -2,     9,     1,     6,     0,    -1,     3,    -6,     9,     1,    -4,     2,     3,    -6,    -4,    -6,   -12,    -6,     0,     0,     4,     1,     3,    -8,   -10,    -1,    -2,    -6,     4,     2,     3,     0,    21,    14,     9,    -2,     2,   -14,   -25,    -5,   -14,    -4,   -10,   -16,   -13,   -14,     2,    -5,    -5,    -4,    -3,    -6,     1,   -10,     1,    -5,    11,    15,     8,     6,     6,     7,    -4,     1,    -3,   -31,   -29,   -10,   -14,    -4,     1,    -7,    -7,     1,    -3,    -2,    -8,    -4,    -3,    -2,    -3,     2,    -8,    -7,     1,     2,     0,     2,     9,     3,    -1,    -2,     0,   -26,   -18,   -13,    -8,    -5,     2,     0,    -1,    -2,    -1,    -1,   -10,    -3,    -4,   -10,    -1,    -1,     2,    -6,     5,     2,     4,     4,     8,     5,    12,     5,     7,   -35,   -23,    -7,   -11,     5,     5,    -4,    14,     2,     1,    -2,    -7,    -1,    -2,   -21,   -15,    -6,     1,     1,    19,     9,     8,    -9,    -6,    -1,     1,     2,   -29,   -40,   -12,    10,     3,     1,    16,   -10,    -3,     1,     2,    -3,    -5,    -3,    -3,   -18,   -18,   -10,   -12,    -6,     9,     4,   -12,     0,     9,    -1,    -6,    -8,   -18,   -19,     7,    14,   -11,    -7,    13,    -5,   -11,     0,     7,    -1,    -6,    -4,    -7,    -8,    -5,   -24,   -26,   -10,    -2,    -5,   -15,     3,     5,     5,   -13,    -9,   -15,   -16,    12,    12,     1,    -3,     0,     1,   -13,    -7,     0,    -7,    -8,    -4,   -11,   -15,   -12,   -18,   -32,   -25,   -19,   -18,    -2,     2,    -3,    -2,   -13,    -6,   -17,    -4,     6,    16,     2,    -5,    -3,     0,    -5,    -7,    -1,     0,    -6,    -6,   -11,    -2,    -7,   -21,   -15,    -8,   -12,     0,     0,    -7,    -1,   -15,   -11,   -10,   -13,     9,     3,    -3,    -2,    -4,     9,     5,    -2,    -1,    -2,     0,    -8,    -8,   -10,    -5,     3,    -4,     1,    -2,    -2,    -7,     1,    -3,    -4,     0,    -5,   -15,    -8,    11,    11,    -1,     0,    11,   -17,    10,    -7,    -2,     0,     2,    -6,   -11,    -1,     4,    -8,     1,     5,     1,    -6,     2,    -9,   -13,    -7,    -6,    -7,   -20,    -8,     8,    15,     0,    -4,    10,    15,    -1,     1,    -1,    -1,    -1,    -4,    -3,   -11,     2,    -4,    11,     2,     3,     2,   -11,    -4,    -8,   -10,   -14,    -8,   -13,   -10,     6,    18,     3,    -1,    -4,    11,    -7,     1,     1,     0,     0,    -2,    -8,    -5,     4,     1,     8,    -1,     2,    -3,    -9,    -1,    -6,    -8,   -11,    -6,    -5,   -16,    -9,     6,    -2,     0,     1,   -10,    -6,    -9,    -2,    -2,     0,     7,    -3,    12,    -3,     1,     9,     1,   -12,    -7,     7,    -4,     4,    -9,    -7,    21,     7,    -9,    -5,     4,     4,    -3,     3,   -13,   -11,    -8,     0,    -2,    -1,     1,    14,    15,     2,    -2,    10,    -2,     6,    -5,     8,    15,     6,    14,     3,    27,    24,     1,   -16,     1,     6,    -4,    -4,     1,    -2,     0,    -2,    -2,     2,    -1,    -1,    -1,    -1,     1,     1,     1,     1,     8,    17,    14,    15,    18,    11,     6,    -3,    -5,    -3,    -5,    -4,     1,    -3,     1,     0,     1,     2),
		    20 => (    0,    -2,    -1,     0,    -2,    -2,     2,     2,     0,     2,     0,    -2,    -2,    -3,    -2,    -3,    -1,     1,     1,     2,    -2,    -1,    -2,    -1,    -1,     0,     2,    -2,    -2,    -3,    -1,     1,     2,     2,     0,    -4,    -8,   -10,   -11,     3,     2,     1,    -1,     9,     5,     5,    -3,    -1,    -1,    -1,    -2,    -1,    -2,     1,    -2,    -1,     0,     2,    -1,     3,     7,    -2,    -3,    -1,    -5,   -10,    -7,    -1,     1,    -4,   -11,    -9,     1,    -1,     2,    -2,    -1,    -3,   -11,    -9,    -3,    -4,     0,     2,     0,     1,    -2,     4,     1,    -9,    -5,    -2,   -10,   -19,    -7,    -7,    -6,   -15,   -11,    -5,    -5,     1,    -5,    -3,   -13,   -13,   -10,   -16,    -6,    -7,   -11,     1,     1,     0,    -4,    -7,    -6,   -17,    -6,    -4,    -6,    -4,     0,     0,   -10,    -8,    -7,    -3,     6,     8,     6,     6,    -4,    -9,    -8,   -10,     1,   -19,    -8,     2,     1,    -1,    -5,    -2,     3,    -8,    -4,   -10,    -9,     0,     2,     2,    -3,    -6,     1,     4,    12,    10,    12,     6,    -3,    -2,   -15,   -11,    -1,   -17,    -8,     0,     0,    -1,    -6,     0,    -1,     0,    -1,    -4,   -10,    -9,    -3,    -3,    -7,     1,    -3,     6,     8,     8,    10,     5,    10,     5,     0,    -2,    -5,   -11,    -3,     6,    -2,    -8,   -11,    -8,    -6,    -3,     0,     1,   -12,    -6,    -3,    -2,    -3,     1,     4,     1,     2,     6,     1,     4,     6,    -3,     4,     1,     0,     4,   -10,     2,     5,   -15,     2,    -7,    -9,    -5,   -10,    -6,   -10,    -8,    -6,    -1,     0,    -1,    -4,    -7,    -4,     1,     5,    -2,     1,     6,     2,     1,    -2,    -7,    -9,    -2,    -3,    -3,     3,    -1,    -9,    -8,   -15,    -4,   -10,    -7,    -9,    -1,    -3,    -5,   -13,   -10,    -6,    -9,   -12,   -12,    -7,    -7,    -6,    -5,    -2,   -13,   -14,     0,    -2,     2,     7,    -1,   -10,   -13,    -6,     0,    -9,   -10,   -12,   -14,   -16,   -16,    -8,   -11,    -7,    -5,   -11,   -10,   -18,   -20,    -6,    -4,    -7,    -6,   -11,    -2,    -1,    12,   -12,     1,    -9,    -3,     5,    -5,   -16,   -12,   -12,   -13,   -12,    -8,    -8,    -4,    -7,    -5,    -5,    -3,    -7,   -10,    -2,    -5,    -3,    -5,    -4,    -2,    -1,     2,   -15,     4,    -5,    -1,    -1,    -6,    -5,    -1,    -4,    -1,     1,     2,     2,    -2,    -1,    -3,     3,     1,     1,    -1,     2,    -3,    -4,    -7,    -6,    -3,     0,     4,    -1,     3,    -1,    -2,     1,    -3,    -8,    -1,    -6,    -3,    -2,     1,     0,    -8,    -4,     0,     8,     1,    -8,     1,     2,     3,    -1,    -1,   -10,    -7,     1,    -1,    -3,   -10,     1,     0,    -2,     2,     2,    -1,   -13,    -9,    -6,    -5,   -15,   -12,    -9,    -1,    -1,    -9,    -4,    -2,    -1,    -8,    -3,     7,   -11,    -1,     1,     1,    -3,   -13,     4,     4,    -9,     3,     3,   -10,   -14,   -16,   -10,   -23,   -23,   -11,    -8,     0,    -2,    -2,     5,     1,    -6,   -10,    -2,     2,   -14,    -5,     2,     0,    -8,    -3,    11,     0,    -8,    -9,    -2,   -14,   -18,   -13,   -18,   -22,   -14,     0,     0,     6,     2,     0,     6,    -4,    -7,    -1,     5,     4,   -19,     3,    -1,    -1,    -8,    -2,     2,     0,     3,     1,    -1,    -1,   -11,   -11,    -6,    -7,    -4,     6,     3,     7,    -1,     4,    -2,    -5,    -4,     6,     4,     2,   -17,     3,    -3,    -2,    -6,    -2,     5,    -3,     2,     3,     3,     3,    -3,    -9,   -11,    -8,     0,     9,     7,     5,    -1,    -5,    -5,    -4,     1,     4,     1,    -1,   -10,    -7,     1,     1,     0,     0,     2,     2,    -2,     7,     4,     4,    -3,    -3,     0,   -10,     0,     6,     1,   -10,   -15,   -10,    -1,     9,     5,     2,     9,   -16,    -7,    -6,    -2,     4,     4,     2,     1,     2,    -4,    -3,    -2,    -4,    -1,    -4,    -5,    -9,    -1,     0,    -6,   -13,    -5,    -1,    -1,    -2,    -1,     5,     4,    -5,    -2,    -2,     2,     1,    -3,     0,    -2,    -1,    -3,    -2,     1,     0,    -4,   -12,    -8,   -14,    -7,     1,    -5,    -6,     1,     2,     1,    -9,    -2,     5,     5,     0,     4,     1,     0,    -2,    -9,     0,     5,     1,    -1,    -2,    -2,    -1,   -10,    -3,    -5,    -3,    -1,   -10,    -2,    -9,     0,     0,    -5,     0,     4,     2,     1,    -2,     0,     1,    -2,     0,    -9,    -8,    -7,    -4,    -3,    -2,   -11,    -8,    -3,     2,     1,     1,    -6,    -4,    -3,     2,     4,     3,    -3,     4,     5,     2,   -13,    -9,    -6,     1,    -2,     1,    -1,    -6,    -7,     3,   -11,    -4,    -4,    -9,   -19,   -14,   -10,    -9,   -11,    -8,    -6,     3,    -2,    -1,    -4,    -4,    -3,    -5,    -5,    -1,    -1,     1,    -1,     1,     0,    -8,   -13,    -7,    -8,    -7,    -7,    -5,    -8,   -14,   -15,   -18,   -16,   -11,   -13,    -5,    -3,   -15,   -10,    -9,   -10,    -6,     1,    -1,     2,    -1,     0,    -1,    -2,     1,   -10,   -12,   -15,    -7,    -5,    -9,    -9,    -2,    -4,    -9,    -8,   -12,   -10,   -15,   -15,   -17,   -13,   -12,   -10,    -4,     2,     0,     0,     1,     0,    -1,     1,     0,     0,     1,    -5,    -8,    -7,    -6,    -1,     1,    -1,    -6,     2,    -3,    -4,    -6,    -4,    -6,    -2,    -4,    -6,    -4,    -2,    -1,     3,    -2),
		    21 => (    2,    -1,    -2,     1,    -1,    -2,     1,    -2,    -2,    -2,    -2,     2,     2,     2,     0,     1,     0,    -2,     2,    -1,     2,    -1,    -1,     0,     2,     0,    -1,    -2,     1,     2,     1,     2,    -2,     1,     2,     0,     2,    -1,    -2,     2,     0,    -6,    11,    12,    -2,    -9,    -3,    -5,     1,    -1,    -1,     2,     2,     1,    -1,    -2,     1,     0,     1,    -2,    -2,     1,    -1,    -1,    -2,   -12,   -11,    -8,   -20,    -5,   -11,   -11,    -2,   -11,    -5,    -3,    -3,   -14,   -18,   -10,    -8,    -4,     1,    -1,     0,    -2,    17,    11,    -1,   -10,    -2,    11,     9,    11,     3,   -15,   -10,    15,    -2,   -14,   -11,    -4,    -5,    -9,    -3,   -24,   -16,   -10,    -9,    -3,     2,     2,    -2,    -2,    15,    15,     2,    -5,    -1,    15,    15,    13,     9,    -4,    -1,     5,    -2,     0,   -12,   -12,    -4,     1,    -6,   -16,    -8,    -9,    -8,   -18,   -19,   -14,    -1,     0,    14,     2,     4,     7,     7,    14,     5,    12,    19,    20,    10,    10,     1,    -6,    -7,    -4,    -7,     3,    -5,   -12,    -9,     7,     1,   -30,   -14,   -12,     0,     0,    -7,     1,     6,     3,    10,    18,     5,     6,    22,     9,     4,     8,     2,     0,    -3,     0,    -1,     0,    -2,   -11,    -6,     8,     0,   -13,   -17,    -8,    -1,   -12,   -17,   -14,   -21,     8,    13,    21,    -7,    -8,     9,     3,     9,    -4,     9,     0,     4,     3,   -10,    -8,     7,    -6,     8,     7,    -4,   -11,   -27,   -17,    -3,   -12,   -16,   -23,   -22,    -2,    14,    15,    -8,   -18,     9,    -9,     3,    12,     8,     6,     2,     8,    11,     4,    -4,    -2,     6,    -2,   -13,   -11,   -29,   -11,     2,    -5,   -16,   -22,   -16,    -7,     0,    11,    -4,    -5,   -10,   -13,    -5,    14,     3,     3,    -1,    10,    14,    -3,     2,     5,     1,    -8,   -11,   -12,   -11,   -17,     1,    -8,   -14,   -21,   -17,   -10,   -10,     0,     7,    -8,   -12,   -14,    -3,     9,     0,    -1,    14,    16,     5,    -3,    -1,    -7,   -10,   -14,   -16,   -10,   -18,     2,     0,    -1,    -5,   -13,     1,    -4,    -6,    13,     5,     1,    -7,   -10,    -2,     3,     0,     2,    18,    27,     7,    -1,    11,   -13,   -17,   -13,   -17,   -14,   -18,    15,     1,     2,   -22,    -9,    -1,     2,    11,    12,     2,    -6,    -6,     0,     5,     0,     5,    12,    11,    16,    10,    -3,     2,   -15,   -16,    -4,   -17,    -5,     2,    14,     1,    -2,   -11,     0,    -7,     6,    11,     5,    -7,   -11,    -5,    -7,    -2,    -5,     1,    -4,     1,    19,    -9,     2,     0,   -12,   -12,   -24,   -19,     5,    11,     1,     0,    -2,     2,     4,    -9,     2,    -8,   -10,     0,    -7,   -10,     3,    -2,    -2,     9,    -1,    -5,    -2,   -21,    -7,     3,    -4,    -5,   -10,   -17,     6,    20,     0,     1,    -2,     2,    -6,   -16,   -11,    -5,     0,    -5,    -2,     3,    -8,     0,     2,     6,     1,    -6,   -12,   -20,   -15,    -4,     3,   -16,   -16,   -23,    -9,    -1,    -5,     0,    -1,     3,   -15,   -14,     3,     1,   -10,   -10,     6,     0,    -5,     0,     8,     7,   -12,   -20,   -20,    -6,    -8,     0,    -1,    -4,    -1,     8,     1,    -7,    -5,     0,    -2,    -3,   -22,   -11,     6,    -2,    -8,    -7,   -12,   -10,     7,     9,     6,     9,   -19,   -16,   -21,   -14,    -1,     3,     7,    13,    14,    11,     0,   -10,   -13,    -2,    -2,    -6,   -22,   -15,   -14,   -24,   -15,   -13,    -8,    -5,     0,    -2,     3,     1,    -6,   -12,   -11,    12,    13,    15,    13,     2,    -1,     5,     9,    -7,     5,     2,     0,     3,   -26,   -19,    -7,    -4,    -3,    -1,     2,     7,     7,    -6,    -8,     6,    -4,    -5,     1,     2,     9,    24,    12,     2,    10,    14,    12,    -5,     2,    -2,    -1,   -12,   -21,    -4,    -1,     7,    -3,     5,    11,    16,     5,    -1,    -6,    -4,     2,     0,     7,    16,    14,    23,     8,     1,    -1,     6,     4,    -1,     0,     5,     4,   -17,    -1,    -4,     4,    -1,     2,    -2,     5,    11,    -5,   -12,    -8,    -5,     8,     5,    -3,    19,    17,    21,    18,    -2,    -5,     7,     5,    -7,     1,     2,     2,   -15,   -12,    -5,     5,    -2,    -3,    10,     3,     5,    -4,    -9,     0,    -9,    11,    -3,     5,    31,    20,    13,    18,     4,     0,     7,    10,    -2,     0,    -2,     2,    -5,    -1,   -12,    -3,     2,     1,   -13,    -3,    -6,    -1,    13,     4,     7,    20,     8,    12,    14,     9,    13,     4,    -1,   -11,   -15,    -9,     9,    -2,    -1,    -2,     0,    -3,   -13,   -11,   -12,    -2,   -16,   -18,     4,    -9,     1,     2,     2,     9,     6,    16,     5,     6,     2,    10,     5,   -12,   -10,     5,     2,     1,     1,     0,    -1,    -7,   -12,   -22,   -25,   -26,   -15,   -38,   -36,   -29,    -3,    -1,    -7,     1,   -14,   -27,   -25,   -31,   -26,   -20,    -8,    -8,    -9,    -7,    -6,     2,     1,     0,    -1,    -6,   -17,   -31,   -29,   -20,   -38,   -38,   -21,   -14,   -19,   -24,    -2,    -2,     5,   -15,   -12,    -4,    -7,   -14,    -1,    -2,     2,     2,    -1,    -1,     2,     2,     0,    -2,    -4,    -4,    -4,     0,    -1,    -3,   -17,   -10,    -3,    -5,    -8,    -4,    -2,    -1,     3,    -2,    -3,     1,    -1,     0,     0,     1,     2,    -2),
		    22 => (    0,    -1,    -1,     0,     0,     0,     0,    -2,     1,     1,     0,     1,    -4,    -6,     4,     4,    -1,    -1,     0,    -2,    -2,     0,     0,     0,     1,     0,     0,    -2,    -2,     0,     1,     2,     1,    -1,    -6,    -6,   -14,   -11,    -6,    -9,    -6,   -13,    -4,     0,     0,    -3,    -6,   -24,   -14,    -8,    -8,    -5,     2,     0,     0,     2,     0,    -1,    -2,    -4,    -8,    -3,    -2,    -8,     5,    11,    13,    12,    10,     7,    -7,    -5,    -3,    -7,   -13,   -15,   -14,    -9,    -6,    -2,     2,    11,     2,     0,     1,     1,    -5,   -14,   -13,    11,     9,    -7,    -1,    20,     8,    14,    14,     5,     2,    -5,     0,    -2,   -13,   -10,    -5,     9,     0,   -13,     1,     3,    -2,     1,    -1,    -1,     0,    -5,    11,    -4,     5,    10,     6,    16,    10,     9,     9,     8,    -1,     3,     5,     8,     4,    -2,    -1,   -10,    -5,    -8,    -6,    -7,    -5,    -6,    -1,     1,     4,     3,     9,     7,    -2,     5,     6,     3,    -1,    -1,     0,     2,     3,     4,    14,     5,    11,    -6,    -4,    -2,     3,    -7,    -7,    -7,    -5,    -5,     0,     0,     3,     1,     0,     4,    -4,     2,    10,     3,     2,    -2,     5,     0,    11,    19,    12,     1,     3,     2,   -12,    -8,    -6,   -14,   -23,    -1,    -3,    -4,    -2,     0,     3,    -7,     1,    -3,     9,     8,     7,     8,     0,     3,     0,     5,     2,   -10,     0,    -2,    -3,    -4,    -9,   -12,    -7,   -23,    -9,     2,    -6,    -1,    -8,     6,    -9,   -11,    -2,    -6,    -3,     1,    -4,     0,    11,     3,    -9,    -4,    -3,    -3,    -3,     2,     6,     6,     2,     0,   -15,   -14,    -9,    -8,    -3,    -6,     1,     0,    -2,   -13,   -12,   -16,   -14,   -11,   -17,   -17,    -1,    -2,    -1,    -8,   -11,   -11,     0,    -4,    -2,    -7,     1,    -5,    -5,   -16,   -18,   -13,     2,    -3,     0,     0,    -1,   -17,   -10,    -4,     2,    -7,   -15,   -18,   -12,   -17,   -11,   -22,   -16,   -16,    -6,     4,     5,     7,     3,    -8,   -23,    -8,    -3,    -4,    -2,    -6,    -2,    -7,    -7,   -14,   -10,   -17,   -17,   -31,   -27,   -28,   -27,   -26,   -23,   -16,   -16,   -22,   -11,    -1,    -8,     7,    -2,    -6,    -5,     6,     6,     0,   -16,    -5,     0,   -11,   -12,   -11,   -22,   -20,   -20,   -31,   -24,   -15,   -13,   -20,    -6,     0,    -4,    -8,    -4,    -5,    -3,     6,    -4,    -2,    -5,    -8,   -20,     4,   -12,    -3,    -1,   -10,    -4,    -8,   -15,   -17,    -9,    -1,    -5,   -10,    -9,     7,    19,    14,     9,    -6,    -3,     1,     9,    -3,    -2,   -12,    -6,     0,     9,     8,     8,     3,    -2,   -11,   -10,    12,    -2,    -5,     4,     6,     7,    12,    17,    19,    21,     4,    11,     5,     6,     1,     6,    -3,     0,    -7,     0,     2,    11,     2,    11,    12,     1,    -5,     0,    10,     9,    16,    10,     1,     6,    14,    13,    10,    -2,    -1,     5,     7,     1,    -3,     3,    -3,    -9,     4,    -2,    -4,    -3,    11,    10,    18,    -2,     2,     9,     2,    14,     5,     9,     6,     1,     4,    -2,     6,     0,    -3,     3,     3,     5,    10,     7,     7,    11,    13,     6,     2,    -4,    19,    16,     4,     2,     0,     7,    -5,     4,     6,    11,     0,    11,     0,     8,    -4,     0,   -12,     3,     8,    -4,     9,     7,     3,    -1,    -8,     4,    -4,   -19,    12,    -3,     9,    -1,     0,    -5,   -16,    -7,    12,     8,    10,    17,     7,     1,   -10,   -12,     0,     3,     4,     7,    -3,    -7,     2,     7,    -8,    10,     1,     6,     0,    -4,    22,    -1,    -7,    -2,   -20,    -5,   -17,     2,     3,     5,     0,    -1,   -15,   -12,   -12,     2,    15,     4,     4,     3,    -8,     0,    -3,     4,    -7,    -1,    -6,    13,    19,    -1,   -10,     9,    -1,     3,     2,   -14,     1,    15,    -2,   -10,    -3,    -6,    -3,    -6,    -7,    -7,    -8,     7,    -5,     1,    -7,    -4,   -10,    11,   -11,    11,     0,     2,     3,     6,    10,     6,    -2,    -1,    -1,     3,    -1,     8,     0,    -6,    -4,    -5,   -18,   -19,   -10,    -8,     1,    -8,     6,     0,     3,   -12,   -10,   -25,    -1,     2,     2,     6,    18,     8,     2,     2,   -10,    -7,     1,    -5,    -1,   -15,    -8,   -22,   -33,    -6,   -14,     2,     1,   -12,   -10,     5,     2,    -3,   -16,   -26,     0,     2,    -1,     3,     4,    -4,    -3,   -13,   -10,    -6,    -4,     0,    -6,    -8,   -23,   -15,   -20,   -16,   -16,    -9,   -27,   -17,   -12,     2,   -11,    -9,   -14,   -25,     1,    -1,    -1,   -13,    -6,   -16,   -10,   -30,   -14,   -17,   -22,   -24,   -16,   -27,   -31,   -28,   -27,   -19,   -10,   -32,   -32,   -20,    -8,    -4,   -18,     3,     4,     0,    -2,     2,     2,     0,    -2,    -1,    -5,    -6,   -12,   -20,   -24,   -14,   -10,   -15,   -17,   -16,   -17,   -23,   -25,   -18,   -22,   -17,    -8,    -6,     0,     6,    10,    11,    -1,     1,     0,     1,    -1,    -2,    -4,    -4,    -2,    -3,    -5,     0,    -2,     1,    -3,    -3,    -6,    -9,   -11,    -8,    -3,    -4,     2,    -8,    -1,    -4,     2,    -2,    -2,    -2,    -1,     2,    -1,    -2,     2,    -1,    -2,     0,     1,    -2,    -3,    -1,     0,    -3,     0,     0,    -1,    -2,     1,    -3,    -5,    -3,     0,     2,     0,     2,     1),
		    23 => (    0,    -1,    -1,    -1,     2,    -2,     0,     0,    -1,     1,     1,     1,    -1,    -3,     1,    -1,     0,     0,    -2,    -2,     0,    -1,    -1,     2,    -2,     2,     0,     1,     1,    -2,     0,     1,    -1,     0,    -1,     1,    -1,    -1,    -6,    -6,    -7,    -4,    -6,    -6,    -6,   -10,    -9,    -3,    -3,    -3,    -2,    -2,     2,     2,     0,     0,     1,    -1,     1,     2,    -2,    -3,     0,    -3,   -13,   -10,     1,     0,    -8,    -6,    -8,   -13,   -20,   -14,   -10,   -11,    -7,    -3,    -5,   -10,    -1,     1,    -1,    -1,     2,     1,    -3,     4,    -4,     9,    14,    20,     9,     5,    -8,    -2,    -1,     2,    -7,     3,     7,    -4,   -24,   -15,    -5,   -16,   -10,   -17,    -5,    -5,     2,     0,    -2,     4,     1,     3,    11,    11,     2,     7,    15,    11,     1,    -3,     2,     3,     3,    -1,     0,     1,   -14,   -20,   -27,   -11,   -13,   -24,   -14,    -3,    -3,     0,     2,     1,     8,     1,     3,    10,     7,     1,     2,     0,     6,     7,     2,    10,     2,     3,     4,    -8,    -9,    -6,   -23,   -21,   -26,   -22,   -11,   -10,    -5,    -2,     2,     3,     4,     7,     3,    13,    13,     3,     9,    12,    13,    -3,    -1,     6,     1,     4,     3,     2,     6,    -3,    -7,   -22,   -23,   -21,    -6,    -6,   -12,    -2,     0,     1,     0,    10,    16,    16,     5,     3,    -3,    -2,     0,    -3,    -7,     6,     2,     0,     9,     5,    -3,    -3,   -18,   -23,   -24,   -26,   -13,    -2,   -11,    -6,    -4,    -2,     3,     6,     1,    13,    12,     9,    -1,   -18,    -7,   -31,   -20,    -6,    -5,     5,     7,     1,     1,    11,   -15,   -17,   -24,   -26,   -18,    -6,   -13,     0,     2,    -4,    -3,    -5,    -4,    -4,    -5,   -24,   -38,   -34,   -21,   -21,    -6,    -3,     8,     9,     5,     3,     0,   -16,   -33,   -23,   -21,   -12,   -10,    -6,   -12,     1,    -1,    -7,     3,     1,   -14,   -25,   -42,   -45,   -27,   -10,     9,     1,     2,     8,    12,    -1,    -1,     5,   -15,   -26,   -33,   -26,    -6,     1,   -10,    -5,    -7,    -4,     2,    -3,    -2,    -4,   -26,   -28,   -25,   -19,    12,     8,    11,    18,    10,    12,     6,     0,   -15,   -16,   -11,   -19,   -17,   -16,   -11,     1,   -13,    -3,    -7,    -2,     2,    -4,    -6,    -9,    -8,    -2,    -4,    12,    11,    18,     8,     3,     0,     2,    -2,     4,   -12,   -16,    -7,   -11,    -9,   -10,    -5,    -7,   -12,    -1,    -6,    -2,     2,    -2,    -4,    -8,     0,     4,    11,    27,    18,     7,     0,    -8,     0,    -2,    12,     2,    -1,   -14,    -6,    -3,    -1,    -1,    -8,    -2,   -13,   -12,    -9,    -6,     0,     1,     1,   -10,     2,    -5,    -5,     0,     5,    -2,    -3,    -7,    -8,     1,     0,    -8,    -3,    -5,    -5,     5,     1,    12,     2,     6,    -1,   -25,    -2,    -7,    -3,     6,     0,    -6,    -1,    -1,    -5,   -19,    -8,   -14,    -8,   -14,    -6,    -1,     0,   -16,     0,     7,    -2,    -3,    -1,    13,     3,     6,    10,   -14,    -2,    -3,     0,     1,     1,    -8,    -7,    -7,   -14,   -25,    -6,   -15,   -16,   -25,   -36,   -21,    -7,   -11,    -2,     6,     1,     6,     2,    12,    14,     9,     7,   -26,   -22,    -5,    -2,     4,     7,     5,    -8,    -6,    -4,     2,    12,     2,    -5,   -25,   -31,   -23,   -24,   -12,    -1,     4,   -10,   -12,    -2,     4,     6,   -10,    -5,   -27,    -5,    -7,    -3,     5,    -3,    12,     7,     8,    19,    -8,    19,     3,    -4,    -2,    -5,   -11,    -8,    -6,     8,    -7,    -6,    -1,     1,     1,    -1,   -12,   -10,   -14,    -8,    -6,    -2,    -1,   -13,     3,     6,     5,    -5,    -5,     7,    -4,    -5,     7,    13,    10,    -4,    -2,   -11,    -4,    -3,     1,    -5,   -10,     1,    -4,     3,    -8,   -13,    -6,     1,    -1,   -11,     4,    -7,     3,     6,    -3,     4,     6,     0,    -8,    -7,    -7,     1,    -6,     1,    -1,     2,    -9,     1,   -14,   -11,    -4,     5,    -4,   -11,    -3,    -3,     0,     4,     1,     0,     1,     3,     4,     4,     7,     1,     5,     9,     1,    -9,    -9,     2,    -7,    -2,     1,    -4,   -10,    -3,    -3,    -8,    -3,    -7,     0,     0,     0,     0,     8,    15,     4,    11,     3,     0,     4,     4,     2,    -1,     0,    -1,     0,   -10,    -4,    -4,     1,    -4,    -2,     4,     5,     4,   -10,    -1,    -2,    -1,     1,     5,    20,    20,     4,     3,    10,     3,     2,     2,     0,    -7,     7,    -3,     1,    -3,    -5,     5,     0,     3,     1,    -7,     2,     8,     1,    -2,     1,     0,    -1,    -5,     4,    -2,    -2,   -15,     7,    -6,    -6,    -5,     5,     0,    -1,    -1,    -6,    -6,    -5,    -2,    -7,    -7,   -12,   -13,   -11,    -7,    -3,     1,    -1,    -2,    -1,     2,    -4,    -3,    -5,     8,    12,    11,    -3,    -5,   -10,   -23,   -10,   -12,    -7,     5,     1,    -1,    10,    -3,   -13,   -19,   -12,     1,    -3,    -2,    -2,     0,    -2,     2,    -5,    -6,    -7,    -5,    -1,    -7,   -10,    -6,    -8,   -14,   -15,   -18,     0,     4,    -4,    -3,     2,    -6,    -9,   -13,     0,     0,    -1,     1,    -1,     1,     1,    -2,     2,    -1,    -2,    -2,    -1,     0,    -3,    -5,   -14,    -9,   -17,     0,    -4,    -1,     1,    -1,     2,    -4,    -2,    -5,    -2,     2,    -2,     2,     0),
		    24 => (    0,    -1,    -2,     1,     2,    -1,     2,    -1,    -2,     0,    -2,    -1,    -7,    -7,    -3,    -4,    -1,     2,     1,     1,     1,    -2,     1,     2,     1,    -2,     0,     0,     1,    -1,     1,     2,     1,    -1,    -7,    -8,    -4,   -11,   -14,    -6,   -21,    -3,     7,    -7,   -14,    -8,   -11,    -4,    -8,    -2,    -4,    -9,    -1,     0,    -1,    -1,    -2,     0,    -3,   -23,   -25,    -5,    -8,   -17,   -18,   -12,   -16,   -22,   -22,    -8,    -3,   -16,   -14,   -13,    -8,   -17,    -8,    -3,    -2,     0,     0,    -3,     1,     0,     2,    -1,    -2,   -19,   -19,     0,    -9,   -18,   -15,   -22,    -2,   -12,   -25,   -15,     0,     0,     9,     6,     7,     0,    -6,    -1,     7,     6,    10,    -6,     1,    -1,    -2,     2,    -1,    -5,     4,   -15,    -2,    -6,    -5,    -1,    -3,     3,    -6,     6,   -10,    -2,     4,    -2,    -8,   -12,     9,     8,    19,    22,    12,     2,   -10,    -3,    -2,     0,    -4,     6,    -8,    -2,    -7,   -11,    -9,    -6,     1,     6,     3,    -5,    -8,    -8,   -17,   -19,    -9,    -4,     6,    -1,    -1,     3,     2,    -1,     1,     2,    -2,    -2,     1,    -4,    -5,     5,    -9,   -13,    -4,     6,     4,    -8,   -10,    -3,    -7,    -6,   -37,   -45,   -19,    -1,    12,     3,     8,     3,   -11,    -4,     1,   -10,    -1,    -2,    -2,    -7,    -3,    -5,    -7,    -6,     3,     2,     1,    -1,     2,     3,    -3,   -23,   -42,   -37,   -11,     7,     6,    11,    20,    14,    -8,   -14,    11,    -8,    -4,    -7,     7,    -5,   -11,   -10,    -7,    -4,    -4,   -12,    -2,    -7,    -4,     7,    -8,   -21,   -37,   -29,    -5,     5,     1,     2,    11,    10,    -6,    -2,     6,   -11,    -1,    -4,     7,    -7,    -7,    -5,    -4,    -7,     1,     2,    -3,    -7,     4,     3,   -14,   -32,   -39,   -23,    -4,    16,     8,    -1,    10,     6,     1,    -1,    -9,    -3,     1,     0,     6,     9,    -5,    -6,   -10,    -5,     3,     0,    -2,     5,     5,    -2,   -27,   -36,   -24,   -13,    13,    13,     3,    -2,     0,     3,     2,    -3,    -3,    -7,    -1,    -5,    -4,     3,    -6,    -6,    -3,    -6,    -1,    -5,     5,     4,    -2,    -5,   -11,   -22,   -15,    -3,     3,    14,    -5,    -1,     0,     3,    -3,    -7,    -7,   -12,     0,     1,     6,    -7,    -6,   -10,    -5,     2,     2,    -3,     0,    -1,     5,    -7,   -24,   -13,   -15,    -3,    13,     7,     1,    -7,    -1,     3,    -9,   -11,    -7,   -13,    -2,    -4,    -4,    -8,    -4,     0,    -2,    -2,     5,    -2,    -1,    -6,     0,   -10,   -12,   -11,   -10,     0,    -6,    -5,    -2,     5,     5,    -2,   -19,    -3,    -8,     0,     0,     0,   -10,    15,     3,    20,    -3,     4,   -11,     5,     1,     0,    -8,   -12,    -7,    -9,    -6,     0,   -10,     3,    -1,    -4,    -2,    -6,    -7,   -14,    -1,    -1,     0,     2,    26,    13,     4,     7,    -7,    -2,    -2,    13,    10,     1,    -8,    -4,   -11,   -11,   -10,     5,    -2,    -1,    -2,   -11,     6,    -4,   -24,   -14,   -10,    -3,     2,     2,     8,     1,   -20,    -3,     9,    11,    19,    12,    23,    -1,    -6,     0,    -8,    -2,     1,    -1,     0,     0,     3,     0,     8,   -15,   -14,   -15,    -6,    -7,    -2,    -1,    -2,   -13,   -13,    -6,     4,    13,    18,    10,    14,     7,    -8,    -1,     2,     0,    -2,     2,    16,    10,     5,    10,     6,    -1,   -17,   -11,     6,    -7,    -3,     1,    -1,   -25,     3,     2,    -2,     3,     3,     1,     1,     2,     9,    -2,     4,     8,     5,     8,    10,     8,     4,     6,     4,    -9,   -18,   -11,     0,    -1,     0,     0,    -2,   -16,    -4,     8,    10,     2,    -2,     2,    -4,    -6,   -10,    -3,     1,     7,     1,     0,     4,    11,    -1,   -11,    -6,    -9,    -2,   -18,    -6,    -1,    -1,    -2,     1,   -18,   -15,    -4,   -10,    -7,   -10,   -17,   -18,   -16,    -4,    -7,     4,    -2,    -7,    -3,   -10,    11,     4,    -6,     2,     2,     3,   -14,    -7,     0,     0,     0,    -4,   -15,    -5,    -7,    -7,    -4,   -15,   -28,   -27,   -10,    -8,    -4,     0,    -6,    -1,    -2,    -1,     6,    -2,    -6,     8,     7,    -2,   -16,    -8,    -2,    -2,     0,    -2,   -13,   -15,    -9,   -12,   -17,   -22,   -20,   -21,    10,    -1,    -7,    -9,    -3,    -1,    -7,    -5,     2,    -9,     7,     9,    11,    -7,     2,    -4,    -2,    -1,    -2,    -1,    -4,   -11,    -6,   -12,   -15,    -6,    -6,     0,     8,     4,    -3,    -2,    -9,     4,    -3,    -2,    -3,   -14,     8,     1,     3,   -10,    -6,    -3,    -1,     1,     1,    -1,    -3,    -6,     2,    -2,   -11,    -3,     0,    -1,    -3,    -2,     0,    -8,    -1,     7,     5,   -12,    -6,   -16,    -1,    10,     7,   -12,    -8,    -3,     1,    -2,     1,    -6,     2,    -3,    -2,    -4,     0,     1,    -3,     1,    -7,     0,     2,   -17,    -1,    -6,   -11,     3,    -3,   -13,   -15,    -4,     3,    -7,    -1,    -2,    -1,     2,    -1,     1,    -2,    -1,    -3,    -3,     0,    -2,     5,     6,     4,     7,     3,   -26,   -18,    -7,    -9,   -13,    -3,   -16,   -19,   -17,    -7,    -4,    -1,     1,     2,     2,     2,    -2,    -2,    -1,     1,    -5,    -7,    -8,    -3,    -7,    -6,    -3,     1,     0,    -2,   -10,   -13,    -3,    -7,    -5,   -11,    -9,     0,     0,    -2,    -2,     0),
		    25 => (   -2,     2,     1,    -2,     1,     0,     1,     2,     0,    -2,    -1,     1,     0,    -3,    -2,     0,     0,     2,    -1,     1,     2,    -2,    -2,    -1,     2,    -2,    -1,     1,     1,    -2,     2,     2,    -1,     2,    -1,     0,     0,     2,    -3,    -5,    -2,    -4,    -2,    -5,    -6,    -9,    -7,    -4,     0,     0,     0,    -1,     2,     1,     2,     1,    -2,     1,     0,    -2,     1,     0,     1,     0,    -4,     0,    -6,    -6,    -5,    -3,    -8,    -1,    -6,    11,     8,    -9,     3,    -1,    -3,    -2,    -3,    -7,    -1,     1,     0,    -2,    -2,     3,     5,    -8,    -4,    -5,    -3,    -3,    -4,    -7,   -10,   -16,    -5,     3,     2,     7,     9,    -6,     4,     9,     3,    -9,    -7,    -3,     8,     1,     1,    -1,    -4,     5,    -3,     1,    -2,    -2,    -3,    -2,    -7,   -23,   -16,   -18,    -1,     8,    -7,     5,     8,     0,    -5,    -1,    -6,     5,     5,     4,     1,   -14,     0,     1,    -6,     1,    -2,    -1,    -3,    -3,    -3,    -8,   -18,   -21,   -10,    -8,    -7,    -3,     1,    -3,    -5,    -1,     0,    -9,    -4,    10,     4,    15,    -3,    -8,     0,     2,     2,    -2,    -4,    -7,     1,    -6,    -4,    -8,   -10,   -29,    -4,    -5,    10,     1,    -1,    -8,     0,     9,     4,    -3,    11,    10,    12,    12,    -1,    -1,    -1,    -1,     1,    -5,    -4,    -3,     3,     0,    -6,   -22,    -4,   -21,    -9,    -3,    -2,     3,     5,     2,    -6,     0,    -3,     5,    10,    11,     8,    18,     3,     2,    -2,    -8,    -9,    -4,    -2,    -2,     5,    -6,    -8,    -6,    -2,     1,    11,    -2,    -3,    -2,    -6,    -6,     3,     2,    -6,     5,    11,    17,    15,    16,     0,     8,    -2,     0,   -10,    -6,    -1,     4,    -6,    -6,     0,    -2,     6,    -4,     5,    -8,     0,    -2,    -6,     2,    -3,    -5,    -2,    -1,    11,    16,    27,    16,     0,    12,     0,    -4,    -2,     0,    -4,    -1,     0,     0,    -4,   -14,     7,    -5,     4,     5,    12,     0,    -5,    -7,     6,     6,     8,    -8,     3,     4,    16,    11,     9,    10,    -2,     1,    -3,    -2,    -1,    -1,     3,    -1,    -1,    -3,     7,    -1,    -1,    -2,    -7,    -7,   -18,   -15,   -13,     3,   -17,    -8,    -2,     2,    -3,     4,    13,     4,     2,     1,     1,    -2,    -5,    -1,     3,     2,     7,     0,     3,    -3,     2,     8,    -5,   -17,   -32,   -35,   -32,   -35,   -32,   -32,   -21,   -10,   -11,     0,     8,   -13,    -2,    -3,     1,     0,    -6,    -2,     7,     6,    -3,     2,     5,    -7,     3,     2,     2,   -14,   -20,   -25,   -34,   -27,   -29,   -29,   -29,   -17,     1,     0,    12,    -7,     4,     1,    -4,     0,    -3,    -5,    -2,     1,    -2,    -5,     6,    -7,    -1,     0,    -4,    -5,   -12,   -26,   -32,   -26,   -22,   -19,   -15,   -13,     2,     2,     0,    -7,     1,    -4,    -6,     0,    -5,   -14,   -12,   -13,    -1,    -3,    -3,    -2,     9,    -5,     2,     4,    -2,     0,   -14,   -21,   -25,   -18,   -14,    -8,    -4,     0,    -2,    -3,     2,    -4,    -6,     7,    -5,   -11,   -19,   -21,    -8,    -9,    -5,    -3,    -1,     1,     5,     0,     4,     2,   -11,   -18,   -26,   -17,   -13,   -12,    -3,    -4,    -7,    -3,     2,    -1,   -13,    16,     5,   -11,   -19,   -20,    -9,   -14,   -16,    -3,     6,    -1,     2,    -2,     6,    11,   -12,   -15,   -21,   -13,    -9,   -14,   -11,    -4,    -8,    -8,     0,    -3,     1,    18,    13,     7,     0,    -2,   -13,   -16,   -13,   -12,    -7,     3,    -3,    -4,    -6,    -6,   -11,    -7,   -21,   -10,    -7,    -9,    -3,    -3,    -9,    -3,     0,    -1,     3,     2,    12,     9,    12,    15,    -2,   -11,     1,    -9,   -10,     6,    -9,     0,    -1,    10,   -11,    -8,   -10,    -5,    -6,    -8,    -3,   -13,    -6,    -6,    -2,    -2,     1,     2,    -4,     9,     9,    17,     8,     1,    -2,     2,     3,     7,     1,     3,    10,    -1,    -4,   -13,    -8,    -5,    -3,     0,    -1,     0,    -4,    -1,     1,    -1,    -1,    -3,    -8,    -7,    -9,     8,     9,     4,    -1,     5,     5,     2,    10,     5,     3,    -4,    -2,    -7,    -8,    -2,    -3,    -3,     0,     1,    -3,     0,     0,     2,    -6,     8,    -1,    -9,     1,     4,     1,     0,     1,    12,     7,    -1,     1,     2,    -8,     1,    -1,    -7,    -9,     0,     1,    -2,     1,    -5,    -1,    -2,    -1,    -1,     7,     5,     7,    -3,     0,    15,    13,    12,     5,    13,     8,     3,     5,     0,    -1,     9,     1,    -1,    -4,     0,    -1,    -1,     2,    -3,   -10,     0,    -1,     0,    -5,    -2,     0,    -8,     3,    10,     2,    16,    11,    10,     9,     5,     1,    -6,    -7,     5,    -5,     2,    -1,    -2,     0,    -1,    -1,   -14,    -5,     2,    -1,     1,     1,     0,   -11,   -10,    -2,    -9,    -6,     8,    -2,    -5,    -5,    -1,   -14,   -12,    -8,    -5,     9,     4,     0,    -4,    -2,    -2,     1,     0,     0,     0,    -2,    -1,     0,    -1,    -5,    -5,   -18,   -18,    -7,    -3,     5,     9,    11,     5,   -14,   -18,    -5,     0,    -5,     0,     1,     2,     2,    -6,     2,    -1,     0,     0,     1,     2,     1,     0,    -4,     0,    -4,     0,    -2,    -1,    -1,     2,     2,    -1,    -3,     0,     1,     1,    -1,    -2,     1,    -2,    -9,     0,     0,    -2,    -2,     0),
		    26 => (    1,    -1,     2,    -1,    -2,    -2,     1,     2,    -1,    -1,     1,    -2,    10,     7,    -1,     1,    -1,    -1,     1,     1,     0,    -1,     1,     0,     1,    -1,     2,    -1,    -2,     2,    -1,     1,    -2,    -1,     7,    10,    11,     7,    22,    19,     3,     9,    -9,     2,    -4,     1,     7,     9,    26,     9,     5,    10,     2,     0,     1,    -2,    -2,     0,     4,     6,    13,    18,     8,    12,    24,    19,    10,    11,   -18,   -12,     0,    -1,    -1,    12,     7,    -1,     8,     8,    15,     8,     2,   -10,    -2,     1,     2,     1,   -21,    -4,    -1,    18,    15,     5,     2,     2,    -3,   -13,   -18,    -3,     8,     5,    -3,     8,     8,     6,    -1,    -6,     2,    18,     9,   -14,   -11,     1,     0,     1,   -19,     0,     0,    14,    -1,    -4,    10,    13,    -5,   -10,   -30,    -8,     1,    -9,     4,    -3,   -10,     1,    -5,     8,     9,    17,    -2,   -20,    11,    17,     2,    -1,   -16,   -12,     6,    -7,   -18,    10,     7,     3,   -12,   -26,   -10,    -6,     1,     0,   -15,    -3,   -15,    -9,    -1,     0,     3,    11,     2,   -10,    23,    15,     0,    -2,     6,    -4,     3,    -6,   -12,     6,    -5,   -18,   -11,   -13,     2,   -14,   -13,    -1,    -6,    -4,    -2,     3,    -4,    -8,    10,     0,     5,    -8,     7,     9,     0,     1,     1,    -8,     4,    -3,    -6,    -3,    -8,   -13,   -13,    -2,    -3,    -6,    -5,    -7,    -2,    -4,   -11,    -3,    -5,    -2,     0,     2,     2,    -1,     4,     7,    -2,     2,   -10,    -8,     6,    -8,   -12,   -12,    -8,   -16,    -2,    -5,    -8,    -6,   -11,   -11,    -8,   -10,   -21,     0,   -18,    -1,    -5,    -4,     6,   -25,    -5,   -17,     2,     0,   -12,     4,     3,   -19,    -5,   -14,   -12,     1,    -2,     2,    -9,    -7,    -3,   -17,   -26,   -23,   -25,   -14,   -15,   -14,   -37,   -13,     3,    -1,    -6,   -18,    -2,    -1,   -15,   -12,    -7,   -14,   -20,   -21,   -12,     5,    -8,    -3,     2,    -1,    -9,   -11,   -19,   -14,    -9,    -7,    -7,    -7,   -12,     9,    11,    17,   -10,   -22,     1,    -1,     1,    -9,    -6,    -7,   -11,    -1,    -2,     3,     7,     5,     3,    12,     4,    -4,    -2,    -6,   -14,   -17,     4,   -10,    -8,     3,     3,    -5,   -12,    -6,     1,     0,    -2,   -10,    -8,   -15,     0,     6,    12,    16,    15,     5,     1,     3,    -2,    -3,     4,    -3,   -11,   -24,   -18,    -5,     8,    17,    12,    -2,   -20,    -4,     2,     0,    -5,    -8,    -8,    -1,    15,     7,     3,    11,    15,     4,     2,    -6,    -4,     0,    -1,     1,    -9,    -7,   -12,    -7,     5,    18,    11,     6,    -6,     2,     0,     2,    -2,   -16,   -13,    11,     5,     6,    12,    17,     5,    10,    -1,    -9,    -2,    -1,     4,    -4,    -4,    -3,    -4,     7,    13,    11,     4,     5,   -16,   -11,     1,     1,    -6,   -18,   -16,    13,    14,    15,    22,    20,    13,     9,    10,     3,    -5,    -9,    -3,     0,    -2,     4,     2,    -4,    13,    11,   -13,    -7,   -21,   -11,     1,    -1,     0,   -15,    -2,     9,     8,    17,    26,    24,    17,    16,    16,     1,     3,    -2,     6,    -3,    -5,    12,     7,     3,    10,    13,    -8,   -13,   -19,   -11,    -2,    -2,    -1,   -14,   -15,     6,     6,    11,     9,     9,    19,     7,    16,    20,     2,    -1,    -3,    -6,    -3,     5,     5,    10,    -1,    -3,    -5,   -15,   -23,   -18,     2,    -1,    -2,    -1,    -9,    -6,    -2,     9,    -5,     6,     5,     0,    14,    20,     6,   -12,     1,     0,    -7,   -11,    -1,    -3,    -5,    -9,   -24,   -17,   -12,   -12,     1,    -1,   -12,     1,     0,   -17,   -12,    -4,   -10,     0,    -3,     7,     6,     3,     0,    -4,    -5,     7,    -7,    -5,    -5,    -1,    -2,    -2,   -11,     3,    -9,   -15,     2,    -3,    -1,   -17,     4,   -13,   -11,   -10,    -8,     2,    -3,    -1,    -3,   -10,     8,    -2,   -11,    -7,    -1,    -5,    -3,    -5,    11,     0,     9,    17,    -3,     0,    -2,     0,    -6,    -8,    -8,    -6,   -11,    -4,    -2,     3,     2,   -10,    13,    13,     1,    -8,    -2,     0,     2,     8,    -2,    -1,    10,    12,    11,     5,    -2,    -5,     1,    -2,     0,    -6,    -8,   -22,   -22,   -14,     6,    -8,     1,    -6,    11,    13,     4,     6,    10,     2,     2,     5,    -4,     8,    -4,     0,    -7,   -18,    -2,    -3,     2,     0,     2,    -2,   -10,   -17,   -21,   -16,    -9,    -5,    -6,     1,    -7,     2,    -2,     4,    -7,     0,    10,    14,     1,   -12,   -19,   -15,   -14,   -14,   -21,     1,     2,     1,    -1,     0,    -6,    -5,    -3,   -14,   -14,   -21,   -23,   -16,    -6,   -10,     2,     7,     9,    10,     3,   -25,   -10,   -24,   -15,   -11,    -7,    -9,     1,     0,     2,    -1,     0,    -2,     0,    -4,    -4,   -13,    -6,    -8,   -11,    -1,    12,     0,   -10,    -4,   -11,   -10,    -4,    -9,   -18,    -6,    -7,    -6,    -5,    -1,     0,    -1,     2,     0,     1,    -2,     0,    -4,    -6,    -3,    -1,    -3,    -8,    -6,    -1,    -2,     0,    -3,    -1,     1,    -1,    -2,    -3,    -4,    -3,    -2,    -3,     1,     0,     2,    -2,     0,    -2,     2,    -2,    -2,     2,     1,    -1,    -1,     0,     1,     2,    -1,    -2,    -1,     0,    -3,     0,    -3,     0,    -4,    -1,    -1,    -1,    -2,     0,     0),
		    27 => (    2,     1,     2,     0,     2,     2,    -1,     2,     1,    -1,    -2,     2,    -1,    -2,    -1,    -1,     1,    -2,    -2,     0,    -2,     2,     0,     0,     0,     1,    -2,     0,    -2,     1,     0,    -2,    -2,    -2,    -1,     2,     2,    -1,     0,   -11,    -8,   -10,    -1,    -2,    -4,    -2,     1,    -1,    -1,    -2,    -3,    -2,     0,    -1,    -2,    -2,    -2,     1,     2,    -3,    -4,     0,     0,    -3,    -3,    -2,    -3,    -6,   -11,    -7,    -2,    -2,    -1,     2,    -1,    -3,     0,    -1,    -4,     0,     1,    -2,     0,     2,     2,    -2,     0,    -5,    -5,    -4,    -4,    -6,   -10,    -9,    -7,   -13,    -9,    -5,    -2,    -3,    -7,    -6,    -1,    -6,     0,    -8,    -6,    -4,    -2,     1,     2,     1,    -2,     2,     0,    -1,   -13,     0,    -3,   -13,   -11,   -16,   -22,   -20,   -18,   -22,   -16,   -17,   -13,    -6,    -5,    -3,     0,    -9,   -14,   -11,    -9,    -6,    -4,     1,    -1,     2,     1,    -8,     2,     3,    -3,   -13,    10,     8,   -11,    -9,   -14,   -13,   -11,   -15,   -19,   -40,   -49,   -32,   -22,    -8,    -1,   -22,   -17,   -16,    -8,     0,    -1,     1,     2,    22,    17,    13,    -6,   -13,    14,    -2,    -8,    -1,     7,     8,     1,   -15,    -3,     2,     9,    -2,     6,    19,    -1,   -28,   -21,   -19,   -14,    -1,    -1,    16,     0,    17,    16,    -5,     0,     1,     2,     7,    12,    10,     7,     0,    -2,    -3,     4,     4,     1,    12,     8,    11,    16,    18,    -1,    -8,   -16,    -8,   -12,    19,     4,    12,     6,   -10,    -9,     3,     7,     2,     1,     5,     3,     4,    -1,     4,     5,    -2,     4,     5,     3,     8,     6,     3,     6,   -11,   -21,    -5,    -1,    12,    -6,     2,     7,     5,     0,     9,     9,    12,    12,     8,    12,     0,    -3,    -1,    -4,     2,    -1,    10,     4,    18,     4,     0,    -2,    -4,   -20,     0,     0,     7,    -1,    -8,    13,    10,     2,     5,     6,     6,     2,    14,     2,    -4,   -17,    -9,     1,    14,    -2,     7,    10,     5,     4,    -5,   -10,   -12,   -13,     3,     1,    -6,    15,    -3,    12,     4,     4,    10,     1,     2,    16,    21,    -3,   -25,   -38,    -6,     4,     7,    -2,    -2,     9,    -4,    -2,    -4,     3,   -18,    -4,     1,     0,     8,     2,     1,     1,    10,    -8,     6,     2,     0,    10,    -3,   -23,   -57,   -38,    -4,     5,    -1,     4,   -17,    -1,     3,    -2,   -21,    -1,    -7,    -5,     3,    -1,    10,     1,    -2,    -9,    -3,     3,     7,    10,     8,     6,    -1,   -35,   -61,   -22,    -7,     2,     0,   -12,   -16,     1,     2,   -16,   -20,    -7,    -5,    -6,    -4,     0,     2,     9,     2,    -2,    -6,    11,     6,     4,     5,    13,   -19,   -51,   -52,    -1,    -2,     3,    -3,   -14,    -2,     0,    -8,    -8,     1,     8,    -5,    -3,    -1,     0,    -2,     8,    -2,    -8,     2,     0,    10,     0,    -3,     0,   -33,   -56,   -13,    -7,   -11,    -2,    -5,    -3,    -2,     4,    -4,    -2,     3,     9,    -1,     0,    -2,     3,     1,     7,    -7,    -9,     0,    -6,     0,    -2,   -13,   -16,   -33,   -19,    -6,    -9,    -6,    -9,    -4,    -7,    -4,     2,    -2,    -5,   -16,   -18,    -8,    -1,    -5,     1,     0,     0,    -6,    -9,    -6,   -22,   -12,    -9,    -9,    -6,    -5,   -17,   -14,    -8,    -5,     1,     1,     9,     3,    -1,     3,     0,   -16,   -21,   -10,     0,   -11,     3,    -2,    13,   -14,   -16,    -3,    -9,   -10,   -11,    -2,    -3,   -13,   -15,    -9,    -2,   -10,     1,     5,     5,     4,    -1,   -14,    -7,   -11,   -24,   -19,     0,    -7,     2,     6,     1,   -16,     2,     8,    -3,   -19,     9,    10,    -6,     0,    -6,    -4,     3,    -4,    -3,    -8,    -8,    -2,    -1,   -11,     3,   -11,   -12,    -6,    -2,    -2,     0,    12,    -3,    -4,    -7,   -18,   -14,    -4,    -1,     2,     2,    -4,    12,    -5,    -2,    -2,   -12,    -8,   -10,    -1,   -10,   -25,   -19,   -19,   -15,    -1,    -6,     2,    -1,     2,    -1,    -9,   -17,   -14,   -13,   -20,    -5,    -8,     2,    11,     4,    -1,     1,    -4,    -4,   -11,    -4,     1,    -2,     5,     4,    -9,     1,    -1,    -7,     0,     1,     1,    -3,    -8,   -11,     4,   -13,    -9,    -3,     1,    -1,    -5,    -5,     3,    -3,     2,    -7,    -5,     4,     4,    -9,    -4,    -6,    -9,    -4,     1,   -20,     1,     0,     1,    -4,   -10,     3,    12,     5,     2,    -8,     5,     9,    -6,   -14,     2,    -7,     1,     1,     1,    -6,    -2,   -11,     1,   -13,    -8,    -4,    -2,   -11,    -1,     0,    -1,     6,    13,    28,    17,    -2,    -5,     1,    -7,    10,    -5,    -4,   -15,   -19,     3,    -4,    -3,    -6,    -2,    -9,     2,    -7,    -4,    -1,    -5,    -1,     1,     2,     2,   -13,    10,     2,   -15,   -11,    -2,     4,     0,   -13,    -6,    10,    -2,     9,     4,     0,     2,     1,    -4,     3,    17,     9,    -9,    -3,     1,     1,     0,     0,     0,    -3,    -8,   -13,   -18,    -7,    10,    14,    -3,   -14,   -11,    -9,     4,     0,     8,     4,    -6,     0,    12,     8,    -2,    -1,    -3,    -4,    -3,    -1,    -2,     0,    -2,     1,     0,    11,    12,     4,     1,     7,     7,     5,     1,     2,    12,    12,    -3,     0,    12,     3,    10,     7,     3,     2,    15,    -2,    -1,    -2,     1),
		    28 => (    0,    -2,    -1,     0,     0,     2,    -2,    -1,     0,    -1,     2,    -2,    -2,    -2,     0,    -2,     2,     1,    -2,     0,    -1,     2,     0,     0,     0,     0,     0,     1,     1,    -2,     1,     2,     0,     2,     1,     0,     2,    -2,    -2,    -9,    -9,   -10,   -10,   -19,   -15,   -19,    -3,    -4,    -1,     4,     1,     1,     1,     0,     1,    -3,     2,     0,     0,    -2,    -3,    -1,    -5,     0,    -7,   -17,   -28,   -25,   -13,   -10,    -4,   -23,   -23,   -20,    -9,   -16,    -9,   -11,   -14,   -11,    -4,    -4,     2,     0,     2,    -2,    -9,    -6,    -4,   -17,   -28,   -34,   -41,   -44,   -28,   -25,    -6,    13,    -7,    -1,    -7,   -14,   -28,   -27,    -7,     4,    10,    12,     8,     0,    -6,    -1,    -1,   -10,    -6,   -17,   -21,   -33,   -16,   -15,    -5,    -6,    -1,   -11,   -11,     6,     5,     0,    -3,    -7,   -10,     5,     9,   -10,    -8,    -8,     7,   -10,    12,    -2,     1,    -1,   -15,   -13,   -11,   -28,     0,    -2,     3,    -1,    -9,    -2,    -4,     0,     7,    -7,    -3,    -2,   -15,    -3,    -3,    11,     7,    -4,    18,    15,   -13,     3,    -1,     0,    -5,   -23,    -8,   -11,     8,     1,     0,    -2,    -2,     4,     4,    -7,    -7,    -3,     3,    -2,     7,    -6,     5,     8,     9,    13,     5,   -10,   -11,     1,    -2,    -8,    -5,   -20,     1,     5,    -2,     8,     2,    -2,     6,    -1,    -4,    -7,   -12,     1,     1,     0,     2,     0,   -11,     9,    16,     5,    -5,    -8,   -16,     2,    -8,   -11,   -17,    -1,    -2,    -5,     5,     5,    -2,     9,    -2,    -9,    -6,     3,    -6,   -17,   -11,     3,     8,     1,     0,    -2,    11,     7,    12,   -10,     8,     8,    -2,    -8,   -19,    -2,   -15,    -3,    -3,    -6,     8,    -2,    -5,    -5,    -7,    -4,   -11,   -15,    -6,     5,   -13,    10,    -5,    -6,    -3,    10,    14,    -1,     6,    -8,    -2,    -3,   -26,   -23,     5,    -3,    -4,     7,    -1,     8,    -6,    -2,    -3,    -8,    17,     3,    -5,    -7,    -4,     3,     2,     0,     2,    21,    11,   -12,     4,    -3,     0,    -2,   -16,    16,     5,     4,    -3,    -2,     5,    -1,     2,    -1,     4,     9,    16,    18,     2,    -1,    -4,    -3,     5,     5,    -2,     6,    25,    25,    13,   -10,     1,    -1,   -11,    19,    11,     8,    -6,     1,    -1,   -11,   -11,    11,    17,    18,    10,    11,     6,    14,    -5,    15,     4,     0,   -16,    -3,     6,    17,     8,   -11,    -1,     0,    -7,    22,     1,     2,    -4,     5,    -7,     1,     3,    16,    11,    17,    15,    13,     9,     8,     9,    13,    -4,   -17,     2,    -8,   -15,    -2,    -6,     1,    -2,    -2,    -3,    16,     5,     3,     5,    -8,   -12,    -2,    20,    12,     9,    17,     8,     1,     8,     7,     7,     5,   -15,   -20,   -11,    -8,   -13,    16,   -16,     0,    -1,    -1,    -6,     0,   -22,   -15,    -5,     5,     2,    13,    14,    10,     9,    16,    11,     5,    10,     7,    -2,    -8,   -11,   -16,     3,     4,   -18,    18,   -36,   -12,    -3,    -2,    -3,    -3,    -5,    -4,     4,     2,     5,     7,    20,     6,    18,    -2,     4,     3,    17,   -11,    -7,     1,   -14,    -7,    -3,    16,   -20,     8,   -30,   -13,    -1,    -2,    -3,   -13,    13,     5,    20,    -3,    -8,     9,    14,    19,    17,    19,    14,     0,    18,     1,   -12,    -5,    -9,    -6,     4,    25,     8,   -15,    -7,   -18,    -2,    -3,    -6,   -16,    15,    -2,    -5,     3,    -3,     2,     9,    12,    25,    30,    13,    11,    -3,    -8,    -6,   -14,    -4,    -8,    -5,     6,    -4,   -17,    -9,    -7,    -2,    -2,   -19,    -8,    -8,    -1,     6,    -4,     7,     3,     3,   -10,     2,    14,     4,    -8,   -18,   -10,     0,    -4,     3,    -4,     6,    -8,    -3,   -21,   -28,    -7,     0,     0,    -7,    -1,    -2,     2,     7,     3,   -14,    -4,    -6,   -11,    -8,    -8,    -4,    -7,    -5,   -11,     0,    -4,     6,    -7,     9,   -11,    -9,   -16,   -17,     1,    -8,    -2,   -12,     3,    -5,     2,    -1,    -7,   -12,     0,   -14,   -20,   -16,   -11,    -9,   -12,   -13,    10,    11,    -6,     1,    -3,    -2,   -11,   -26,   -16,   -28,    -5,    -5,    -4,    -6,    -1,     4,   -12,    -4,     1,     2,    -2,    -6,   -13,    -8,   -15,   -11,    -3,   -10,   -14,    -4,    -6,    -2,    11,   -10,   -14,   -20,     4,   -12,    -1,    -1,    -1,    -9,     4,     1,     0,   -15,    -1,     3,     7,   -10,    -8,    -9,    -2,   -12,    -2,    -1,     1,     0,     9,    15,    -9,     4,     9,    -9,     4,   -17,    -1,     2,     2,    -8,    -6,   -28,   -21,   -18,   -25,   -15,    -1,     0,    -4,    -1,    -3,   -11,    -7,   -13,   -18,    -9,    12,    -5,   -16,    -6,     3,    -6,    -9,    -4,    -2,     1,    -1,    -8,    -6,    -6,    -2,    12,     9,    -4,    -2,    17,     2,   -16,    -8,    -1,     6,     9,     0,     5,   -11,    -6,   -11,   -16,   -11,   -17,   -11,    -7,    -1,     0,     1,     1,    -7,    -7,   -15,   -20,   -20,   -24,   -35,   -28,   -14,   -12,   -12,   -13,   -34,   -18,   -11,   -15,   -27,   -21,   -12,    -8,    -8,     0,    -2,     0,    -2,    -1,     1,     1,    -1,     0,    -2,    -2,    -9,   -15,   -17,   -10,    -2,    -5,   -13,   -15,   -18,   -11,   -12,    -7,    -9,     1,    -2,    -1,     0,     0,     0,     2,    -1),
		    29 => (    2,     0,     1,    -2,     0,     0,    -2,     2,     0,     2,    -3,     0,     2,     2,    -2,     2,     0,    -1,    -1,    -2,    -1,    -2,    -1,     2,     0,     0,    -1,    -2,     0,     0,     2,     0,    -2,     1,     0,     1,     1,    -2,     0,    -4,    -6,    -4,     1,    -3,    -8,   -11,    -9,    -5,     2,    -4,    -1,    -1,     2,    -2,     1,    -2,     0,     2,    -1,    -3,    -4,     0,    -1,    -5,    -2,    -4,    -4,    -8,    -1,    -1,   -15,   -11,    -9,    -3,    -3,    -2,   -18,    -7,   -12,    -7,    -3,    -2,     0,     2,    -1,     1,     1,    -3,    -6,   -16,   -15,   -13,   -17,   -17,   -30,   -30,   -20,   -23,   -44,   -17,   -22,   -32,   -24,   -16,   -25,   -27,   -18,   -10,    -7,    -3,    -1,     1,     2,    -1,    -7,    -7,    -8,   -26,   -36,   -13,   -16,   -20,    -9,    -6,    -4,    -3,    -7,     3,    -4,   -15,    -5,   -37,   -32,    -9,   -14,    -7,    -5,   -18,   -12,    -2,     1,    -2,    -1,    -3,    -2,   -10,   -12,   -12,    -6,     2,     3,    10,     2,     7,     5,    -3,     3,     6,    12,    12,     4,   -16,   -17,   -15,    -5,   -12,    -9,     1,    -2,     2,    -2,   -10,    -9,   -17,    -6,   -12,     0,    11,     5,    -6,   -11,     2,     3,     6,     4,    -1,    15,    10,    11,    -4,    -5,     7,     2,    -4,    -9,   -15,    -1,    -2,   -12,    -8,   -12,   -14,   -17,   -15,     0,     4,     2,    -6,     0,    -9,    -1,    -6,    -4,    -1,     0,     4,    -5,   -10,   -12,    -3,     2,     7,   -10,    -5,    -8,    -9,    -5,    -4,    -4,   -13,     3,    -3,     5,    12,     8,    -3,    -3,    -2,    -6,    -3,    -2,    -4,     2,    -6,   -17,   -14,   -15,    -9,     5,    -2,   -12,    -4,    -2,    -9,     5,    14,    14,     6,     7,     0,     6,    13,    -2,    -2,    -4,    -7,    -7,    -8,     4,    10,     9,    -5,    -2,    -5,   -13,   -20,   -12,   -17,   -27,   -10,     1,   -12,   -11,     8,    30,    16,    18,    11,     2,     3,    -4,    -5,     4,    -5,    -5,     4,    22,    18,     2,    -6,    -7,    -5,    -9,    -7,    -8,     4,    -8,    -5,     2,   -24,    -2,     1,    16,    17,    16,     2,    -8,    -2,    -2,     3,    -3,     7,    11,     6,    25,    17,     1,   -12,    -7,    -2,     6,     5,     2,    13,    -3,    -7,     2,    -6,     3,    -5,    12,    10,    14,    -4,    -1,    -3,    -4,    -1,    -1,     5,    25,    18,    10,     2,     4,    -4,     5,    -2,     3,     5,    -7,    -8,   -10,    -6,    -1,    -7,    -4,    -7,     9,    14,    -2,     0,    -6,    -7,    -3,     2,     1,    19,    23,    25,    11,     3,     5,    -6,     0,     4,     6,     3,    -1,    -4,    -8,    -4,     1,    -8,   -10,    -7,     2,     2,     9,     1,     2,     3,    -3,     2,     9,    22,    26,    18,    17,     5,     7,     7,     6,     0,    -6,   -10,    -8,    -8,     1,     1,     2,     2,   -17,    -7,    -3,    -4,     6,    -2,    -9,    -4,    -4,    -1,     7,    24,    24,    14,    15,     5,    14,     8,    12,     5,    -8,   -16,   -17,    -7,    -2,    -4,     1,    -4,   -16,   -14,    -4,    -8,    10,     4,     7,    -7,     8,     6,    11,    11,    21,    15,     1,     7,    14,    13,    18,     1,    -5,    -9,   -21,   -15,    -4,    -6,    -1,     0,   -15,    -3,    -6,   -14,    10,    13,    -3,     4,     2,    17,    12,     8,    19,     7,     3,     8,    11,     8,    13,    -1,    -3,    -9,   -20,    -8,   -12,    -5,     7,    -1,   -16,    -7,   -15,   -16,    12,    15,    14,     9,     7,     3,    -1,     3,     3,     5,     1,    20,     8,    13,     9,    -6,    -1,   -13,   -24,   -11,   -12,   -12,     0,     0,   -21,    -5,   -18,   -16,     7,    15,    10,    12,     6,     3,    -3,     1,    -9,     2,    17,    12,     7,     1,     1,     1,     5,    -2,    -6,    -4,    -6,    -5,     1,    -2,   -19,    -8,   -18,   -11,    -9,     3,    11,     3,    -5,     1,     5,    -5,    -9,    -3,     7,     4,     0,     0,    -2,    -6,    -5,     0,    -2,     6,    -7,     1,     0,     1,   -18,    -8,   -15,    -1,    -6,     2,   -10,    -4,    -7,     2,     4,    -8,    -9,     7,     1,     0,   -10,    -7,    -4,    -5,    -9,    -4,     4,     0,   -16,     0,    -1,     0,   -12,    10,   -10,   -15,    -5,    -7,    -7,    -3,    -3,     1,     2,   -13,    -4,     2,   -12,   -13,   -15,    -7,    -7,   -14,   -10,    -8,     3,   -11,    -4,    -1,     0,     1,    -8,     3,    -6,    -9,    -2,   -12,   -14,   -13,   -12,    -1,     4,    -2,     1,    -8,   -14,   -11,   -11,    -9,     9,   -10,   -11,   -14,     2,    -3,    -9,    -1,    -2,     2,   -11,   -15,    -4,     3,   -12,   -12,    -5,    -6,    -5,    -5,     2,     0,    -7,   -17,   -14,    -9,   -11,   -11,    -6,    -6,     0,    -6,     0,    -2,    -1,    -1,    -1,     1,     8,    -5,    -3,    -4,   -13,   -20,   -11,     0,    -8,    -7,     0,    -5,    -5,   -17,     2,    -5,    -3,   -11,    -6,    -6,     0,     9,    -4,     0,    -3,     1,    -2,    -1,    -1,    14,    -7,   -14,   -10,   -12,    -9,    -8,    -9,     0,     2,    -1,     0,    -4,    11,     7,     6,   -14,    -1,     2,    -2,     2,     2,     2,     2,    -2,     2,    -1,    -1,    -2,    -1,    -4,     7,     8,     4,     5,     3,     1,     0,    10,     4,    -3,    -2,    -9,     0,     0,    -4,    -9,    -3,    -8,     0,     0,     0,    -1),
		    30 => (    2,    -2,    -1,     0,    -2,    -1,     2,     1,     0,     0,     0,    -2,     1,    -1,    -4,     0,     0,    -1,    -2,    -1,    -2,    -1,    -2,     1,     1,     2,    -2,     2,    -2,    -2,     0,     0,     2,     0,    -1,   -11,   -10,   -16,   -10,     8,     3,     2,    -7,    10,    14,    10,    -6,    -3,    -2,    -3,    -3,    -2,     0,     1,    -1,     1,     0,     0,     1,    14,    13,     0,    -2,    -2,   -10,   -12,   -19,   -24,   -14,   -21,   -18,   -31,   -26,   -28,   -18,   -15,   -14,   -12,   -17,   -10,    -6,    -5,     0,    -1,     1,     1,     0,     9,    -5,    -9,    -9,   -14,   -13,    -5,   -16,     3,     8,    11,    -6,   -21,    -7,    -5,   -18,   -25,    -6,   -11,   -10,   -11,   -14,    -2,    -8,    -1,     2,    -1,    -8,   -17,    -4,   -21,     2,     0,    -3,     2,     5,    -2,     3,     2,    -8,    -9,   -18,    -1,     0,     8,     1,    -1,    -6,   -11,   -20,   -24,   -10,    -2,    -2,    -1,    -4,   -12,    -3,    -5,     8,     5,    -1,    -7,     5,    -4,   -13,   -13,    -5,    -9,   -12,    -3,     5,     6,    -9,    -8,     2,   -15,    -1,   -30,   -18,    -2,    -2,     0,    -3,    -1,    -3,     0,     1,     8,     4,   -21,    -1,    -7,   -15,     2,    -5,    -3,    -5,    -1,     0,     2,    -6,     0,     4,    -1,     6,   -26,    -7,    -1,     2,    -6,    -1,    -8,    -2,    -2,     0,     0,   -11,     1,    -2,    13,    -4,     9,    -1,    -7,     3,    -1,     7,    10,     4,    13,     7,    17,     3,     0,   -16,     0,    21,   -16,    10,     3,    -6,   -17,   -14,    -6,    -3,     0,    11,     0,     4,    -2,     2,    14,    13,    15,     3,    13,    13,    13,    13,     1,     2,   -13,   -23,    -7,    -2,    -1,    17,   -13,   -12,    -8,   -10,   -12,    -1,     6,     4,     0,     0,    -1,     7,     6,     9,     6,    -6,     2,    17,     8,    -2,     0,     4,   -19,   -10,    -3,    -4,    -3,    15,     8,   -15,    -8,     6,    -1,    -2,    -2,     2,    -4,    -6,    -3,     0,    11,     5,    12,     1,     0,     6,     7,     2,   -10,    -9,   -20,   -25,    -1,    -2,    17,   -13,    -3,   -28,     1,     4,     4,     4,    -8,    -6,   -12,   -11,     2,    -6,    -9,    -5,    -5,    -6,    -8,     1,    14,     3,   -16,   -21,   -20,   -16,    -2,    -1,     3,   -11,    -3,    -6,     3,     9,     7,    -1,     4,    -3,   -16,    -6,    -3,   -16,    -9,    -3,    -6,    -7,    -5,    -1,    10,    12,     0,   -11,    -5,    -9,    -7,    -2,     4,     0,     8,    13,     5,    18,    10,     0,     8,     0,    -9,    -3,   -14,    -6,   -15,    -4,     7,     2,     4,   -14,     5,     0,    -1,   -12,    -5,   -11,   -11,     1,     0,    -1,    -2,    21,    24,    25,    11,     8,    11,    13,     4,     0,   -10,   -12,    -2,   -12,    -1,     1,     6,    -5,   -16,     0,    -7,     6,   -16,   -22,     0,     1,     0,   -10,    -8,    15,    27,     8,    16,    18,    27,    16,    -5,    13,    -9,    -9,    -5,    -8,     0,    -2,    -5,    -2,   -11,     2,     4,    -1,   -12,   -23,   -12,    -2,    -1,    -6,   -19,    17,    18,    11,    11,    21,    23,     9,    19,    13,    -8,     3,     5,    -7,    -4,    -1,    -7,    -5,   -14,   -16,     9,   -17,   -26,   -33,    18,     1,    -1,    -6,   -24,     6,     7,    -5,    10,     5,    10,    15,    15,     0,    -8,    -3,    -2,    -1,     1,     1,     1,     0,   -16,     5,    -5,   -18,   -19,   -17,    25,    -2,    -2,    -4,   -27,     0,    -3,    -3,     1,    11,     5,     8,     2,     6,    -1,    -2,     1,    -5,    -8,    -7,    -6,    -7,    -6,     0,    -6,    -9,   -15,   -17,    -6,     1,     6,    -7,   -19,    -9,    -3,    -4,    -2,    -4,   -14,    -7,    -2,    11,     3,    -1,     0,    -5,   -10,    -3,     0,    -7,     1,     1,    -8,    -8,   -27,   -15,    -6,     1,     9,    -6,   -22,    -6,    -1,    -4,    -8,   -13,   -15,    -5,     4,    -2,     3,    10,     5,    -2,    -7,     0,    -7,    -7,    -5,    -5,    -5,    -9,   -24,     0,    -2,    -2,     2,   -19,   -13,   -14,    -3,     7,     3,    -6,    -6,    -5,    -4,     5,    14,    11,    13,    12,     3,    -6,   -17,   -14,    -6,     2,    -5,    -7,    -7,    16,     5,     0,     1,   -26,    -8,   -25,    -8,     0,     5,    15,    -1,     6,     6,    21,     8,    16,    14,     2,    -1,    -7,    -9,     1,     5,     9,    10,   -11,    -7,     9,     5,     1,    -2,    -7,   -26,   -21,    -5,     5,    -4,     0,    -6,     3,     3,     5,     6,    10,     2,     8,    -8,    -7,    -6,    -6,     6,    -4,    -9,   -11,    -8,   -19,     0,    -1,     0,    -3,    -6,    -3,     8,    -7,   -12,   -15,   -23,   -22,   -15,     6,    17,    16,    14,    13,    -2,    -6,   -24,   -17,    -8,   -12,   -14,    -8,     0,    -2,     2,     1,     2,     0,    -8,   -41,   -33,    -8,    -3,    -3,   -26,   -20,   -14,    -2,    -6,    -8,   -12,    -4,    -2,   -16,   -26,   -20,   -18,   -11,    -5,     1,    -1,     2,    -1,     1,     1,     2,    -1,   -21,   -18,   -26,    -9,   -12,   -21,   -20,   -10,   -12,   -12,   -21,   -18,   -12,   -29,   -28,   -13,   -18,   -20,    -9,   -11,    -4,    -1,     0,    -1,     0,    -2,     1,    -1,     1,     0,    -3,    -2,    -8,    -5,     1,     1,     1,    -7,     0,     0,    -4,    -5,    -6,    -6,    -3,    -9,   -10,    -8,    -1,     2,    -2,     2),
		    31 => (    2,    -2,    -1,    -1,     0,    -2,     1,     1,    -1,    -1,     1,    -2,     1,     2,    -1,     2,    -2,    -2,     2,    -1,     0,    -2,    -2,    -2,     0,     1,     2,     2,    -1,    -1,     1,     2,     2,    -2,    -1,    -2,    -1,     0,    -3,    -3,    -3,   -10,     4,     5,     1,    -6,    -3,     1,    -1,     1,     0,     0,     2,     3,     1,    -1,    -2,    -2,    -1,     0,    -2,     1,    -2,     2,    -7,   -12,    -8,    -8,   -16,     6,    -4,    -1,     6,     1,     4,    13,    13,   -22,   -18,   -11,    -4,    -5,     2,    -2,     0,     0,    10,     8,     0,   -10,   -15,     7,    11,    11,    -1,   -15,    -6,    -8,     1,    11,     2,     0,    -1,    12,    10,    -5,    -2,    -7,   -10,    -2,    -2,     0,    -1,    -2,    12,    10,     8,    13,     0,     1,     7,     2,     8,    -1,    -1,     7,    -1,    -1,     1,    13,    18,    12,    -2,    -2,     2,    -2,    -7,   -13,   -16,   -12,     2,     2,     6,     3,    13,    15,    11,    12,    -5,   -12,    -5,    -6,    -1,    -2,    -8,    -1,    -4,    -5,     1,    13,     5,    -4,    -4,     8,    -4,   -18,   -13,   -12,     1,    -2,   -10,     4,    15,    13,    14,    10,    -6,    -7,    -1,    -3,    -9,    -5,    -6,    -9,     2,     0,     2,     5,     3,    -8,    -8,     1,    -1,    -7,   -17,    -2,     1,    -6,   -17,    -7,   -24,     2,    13,    14,    -9,    -7,    -8,    -3,     1,     5,     4,     1,     2,   -11,    -1,     5,     5,    -3,     0,     9,    -3,   -14,   -32,   -18,     1,   -16,   -18,   -23,   -22,   -10,     5,     0,   -11,    -8,    -1,    -2,    13,    11,    13,    -2,    -3,    -5,     5,     2,   -10,    -5,     7,     1,    -3,   -13,   -45,    -9,     2,    -5,   -15,   -25,   -20,   -10,   -13,    -5,   -12,    -9,    -2,     4,    15,    16,    11,    -4,    -1,    -6,     1,     2,    -7,   -14,     1,    -5,   -11,   -13,   -20,   -11,     0,    -4,   -14,    -7,   -19,   -14,   -14,    -8,   -10,   -18,   -10,    -5,    18,    16,     9,    -2,    -3,     5,    -5,    -7,    -9,   -10,   -14,   -14,   -12,    -8,    -7,    -3,    -2,     3,    -1,   -11,   -12,   -15,   -20,   -19,   -18,   -12,   -14,   -11,     0,    13,     5,     8,    -6,    -3,    -5,   -10,     2,    -9,    -5,   -17,   -17,    -9,   -10,    13,     0,    -2,   -21,    -6,    -3,   -13,   -12,   -26,   -18,   -15,    -8,    -7,     1,    14,    -3,     1,    10,     2,    -5,    -4,     5,   -12,   -12,    -7,   -12,    -4,     2,    11,     1,     1,   -18,     6,    -5,   -15,    -9,   -15,   -12,    -9,    -8,   -11,     1,    -2,     5,     6,    15,    11,    -1,    -4,    -5,   -23,   -18,   -17,   -16,     2,     2,    -1,    -2,    -1,     4,     2,    -9,   -10,   -13,    -8,   -12,    -7,   -13,   -11,     4,    -2,     1,     4,     3,     3,    -5,   -14,    -5,   -16,   -12,    -9,   -12,   -12,    -5,    -1,     0,     0,     3,    -9,   -17,   -14,   -14,   -16,   -11,    -2,    -2,    -2,    -1,     5,     4,     2,     6,     6,     3,    -7,   -14,   -26,   -22,   -17,   -42,   -21,   -11,    -8,    -2,     0,     5,   -18,   -16,    -2,    -6,   -11,    -6,     4,    -5,    -7,    -3,     2,     2,    -1,     6,     0,    -3,    -4,   -10,   -18,   -10,    -8,     3,   -14,    -8,   -10,     2,     0,    -7,   -19,    -9,    -6,   -11,   -20,     4,     1,     6,     7,    -6,    -6,    12,     9,     7,     3,    -1,     0,    -4,     6,     5,    -3,     5,    -7,   -11,   -11,    -1,     1,     2,   -22,   -14,   -14,   -29,   -19,     0,     8,     9,    -4,   -11,    -7,     3,    15,    12,    -4,     3,   -14,    -8,    -4,    -3,     4,     5,    -1,   -10,     1,    -2,     0,    -4,   -23,   -25,     1,     1,    -1,     7,    11,    10,    -3,    -7,     3,     6,     6,     5,    -6,    -8,   -17,   -13,     0,    10,    10,    13,     6,   -12,    -3,    -2,     1,    -8,   -23,    -4,    13,    15,    20,     4,    13,    12,     1,     6,     9,     5,     3,     3,    -8,     3,    -4,     4,     6,    13,    11,    13,     1,    -4,     0,     7,     5,    -3,    -1,    -4,     7,    11,    14,    19,    19,     9,     0,     7,    17,     0,    -7,     3,    -6,     3,    -1,     7,     9,    10,     2,     3,     6,    -8,     1,     3,     4,    -6,    -2,    -3,    11,    13,    14,    11,    18,     8,     8,     7,    15,   -16,   -10,    -2,    -4,     3,     7,    13,     9,    -9,    -4,     7,     0,     2,     0,     1,     1,    -3,    -3,    -6,     4,     4,     0,     4,    18,    11,    10,    12,    -1,   -14,    -7,   -12,     5,    -5,    -4,     6,     1,    -4,   -11,   -13,   -10,    16,    -2,     1,    -2,     2,    -3,   -10,     1,    -5,     2,    -3,     6,     5,   -13,    -4,    -1,   -15,   -14,   -14,     3,    -3,   -13,    -5,     7,    -2,   -16,   -16,     1,     3,     2,    -2,     1,     0,    -4,   -11,   -18,   -11,   -25,     2,   -10,    -3,   -11,     8,     0,   -13,   -16,   -19,   -26,   -29,   -22,   -41,   -15,   -10,    -7,    -3,    -4,    -5,    -1,     0,    -2,    -1,    -3,   -13,   -27,   -38,   -41,   -29,   -27,     4,     1,   -16,   -16,   -16,   -16,   -11,   -21,   -11,    -3,    -7,    -8,    -2,    -3,     0,    -1,    -1,     2,    -2,     0,     0,     2,    -2,    -3,     0,     2,     1,    -2,   -16,   -13,     1,    -4,   -12,    -4,    -5,    -1,     0,     0,     2,    -2,    -1,     2,     1,    -2,     2,     2),
		    32 => (    0,     2,     1,    -1,    -1,     0,     0,     1,     0,    -1,    -1,    -2,    -5,    -4,     2,     0,     0,    -2,     0,     0,    -1,     2,     2,    -1,     1,     1,     2,     1,     0,    -2,    -1,     2,     0,     0,     2,     1,   -10,    -6,    -5,    -2,    -4,    -4,   -15,     1,     2,    -4,    -2,   -12,    -6,    -4,    -7,    -1,     2,    -3,    -1,    -1,     1,    -2,    -1,    -3,    -3,    -1,    -1,    -7,    -3,     2,     3,    -3,     3,    -4,    -2,    -6,    -7,    -9,     3,    -1,   -10,    -4,    -3,     1,     0,     4,     2,     0,    -1,    -2,    -1,    -4,    -9,     7,     4,     3,    -7,    -7,   -13,    -8,   -14,   -18,   -11,    -6,   -19,   -22,   -15,    -5,   -15,   -15,    -6,    -1,     0,    -1,     1,    -1,    -2,    -1,    -4,    -3,     9,    11,    15,    12,    12,     9,     0,     3,     6,    -6,    -7,    -4,    -4,   -14,    -4,    -2,   -11,   -11,   -15,    -7,    -5,    -4,    -7,     0,    -2,    -2,     3,     3,     4,    -1,     3,     3,     6,     9,     6,     5,    -2,    -8,   -12,   -16,    -4,    -2,    -9,    -8,    -6,    -4,   -11,    -8,    -1,     1,    -5,    -5,     1,    -1,    -6,     9,     9,     9,    15,    -1,    -3,     1,    -1,     1,    -6,    -5,    -6,    -7,    -1,     0,    -1,     0,    -9,    -4,    -3,   -10,    -4,    -7,    -4,     0,     1,     0,     2,    15,    15,     5,    15,     7,    14,    -1,    -6,    -1,     7,    -2,   -10,    -3,    -3,   -10,     0,    -4,    -5,    -4,    -8,   -22,   -14,    -7,    -9,    -3,    -6,     4,     0,     5,     7,     5,    13,    10,     7,     8,     3,    -2,     6,    -3,     7,    -4,   -15,    -6,    -9,    -4,    -5,   -13,     1,    -8,   -15,    -8,   -13,    -5,     2,    -3,    -2,    -4,     1,     8,     2,     3,    -3,    -5,   -16,    -9,    -6,    -7,     3,     1,    -4,   -11,    -4,    -1,     0,    -3,     3,    -4,   -14,    -7,     4,    -1,     0,    -2,     1,   -15,    -8,     0,     6,     1,    -4,   -14,   -11,   -27,   -25,   -11,    -2,     0,    -4,    -5,    -4,    -4,     4,    -9,   -10,    -1,    -6,    -6,    -7,    -1,     2,    -2,    -6,    -9,   -11,    -9,    -3,    -4,    -5,   -14,    -3,    -7,   -24,   -12,    -6,    -3,    -1,    -8,    -6,    -1,    -4,    -9,    -1,    -4,     0,     1,   -17,    -4,     1,    -1,    -2,     1,   -13,   -24,   -18,   -16,   -13,   -13,    -9,    -4,    -8,   -13,    -7,   -13,    -5,    -2,    -9,     1,    -7,    -6,     7,     2,    14,     4,    -3,    -3,    -2,     0,    -1,    -4,    -4,   -23,   -28,   -24,   -17,   -16,   -11,     1,    -1,    -2,    -5,   -15,    -9,   -10,    -7,     0,     6,    -3,    10,    15,    21,    12,     1,    -5,     2,    -5,    -5,    -3,   -11,   -19,   -27,   -19,   -15,    -9,     8,     3,    -6,   -13,    -2,    -8,   -11,   -15,    -4,    12,     2,     3,    10,     6,     4,     2,     6,    10,     2,    -7,     7,     7,    -8,   -18,   -15,    -3,     0,     4,     9,    -1,     4,     8,     7,     1,    -4,     2,     3,    20,    15,     8,     1,     9,    13,    12,     9,    15,    -1,    -3,     9,     1,    -6,   -19,    -3,     1,     0,     0,     4,     2,     2,     1,     0,    -5,   -14,     2,    11,    16,     3,    11,    11,    12,     3,    20,     6,     7,     2,    -2,    13,    -3,   -11,    -4,     4,    10,     5,    12,    -1,     0,    -8,    -8,     5,    -3,   -17,    10,    16,    -3,    -1,     7,    -2,    -2,   -13,    12,    -2,     9,     1,     2,     2,    10,   -15,     1,     7,     5,     6,    -2,    -7,    -5,     2,    -9,     1,    -6,     5,    13,     9,    -9,   -12,    -4,    -6,    -6,     5,    15,     2,    21,    -2,   -10,    -6,    -5,   -15,     0,     4,    10,     3,    -6,    -8,    -1,    -4,     1,    -5,    -1,     8,    10,     1,    -8,   -12,   -15,     2,    -9,   -14,     1,    14,    16,    -2,    -9,    -1,    -1,   -11,     0,     6,     5,     4,    -8,   -11,     0,     2,     7,    -5,     0,     3,    -3,    -2,    -8,   -12,   -12,    -9,   -12,   -17,    -2,     3,     1,     0,     2,     3,     2,   -16,   -10,    -3,    -9,     6,    -2,    -3,     3,     0,     3,    -1,     7,    10,     0,     2,    -6,     0,     2,    -7,     2,   -10,    -2,     4,    -2,     0,     1,    -1,     7,   -12,   -19,    -9,   -10,    -8,    -8,    -4,     9,     2,    12,    10,    -1,     0,     4,    -1,    -6,     3,     1,   -12,     1,     1,    -2,    -7,     0,     0,     1,    -2,     8,   -12,   -17,   -12,    -9,    -9,     1,     5,     4,    14,     9,     2,     2,     4,     7,    -5,    -4,    -5,    -3,     3,     5,     3,     5,    -8,     0,     1,     1,   -12,    -9,   -19,   -13,   -17,    -7,   -13,   -16,   -15,   -11,   -10,   -11,    -4,    -5,   -15,    -4,     2,     5,     3,    -5,    -1,     5,     8,    -1,     1,     1,    -1,    -2,     1,    -1,    -4,    -4,    -3,    -2,    -8,   -18,   -25,   -18,   -17,   -31,    -2,    -2,    -9,     1,    -5,     7,     7,     5,    -7,    -2,     3,     2,     2,     0,     1,    -2,     1,    -1,    -1,    -8,    -8,    -7,    -7,   -15,    -3,    -4,    -8,    -7,   -10,    -7,   -13,   -17,   -13,    -8,    -7,    -6,    -8,     1,     0,     0,    -1,     0,    -3,     1,     2,    -2,    -2,     1,     1,     0,    -3,     0,    -5,    -4,    -5,    -9,    -7,     2,     0,    -4,    -2,    -2,    -3,    -7,    -6,    -1,     2,     0,    -1,     2),
		    33 => (   -2,    -1,     0,     2,     1,     2,     0,     2,     2,    -1,     2,     0,     0,    -2,    -3,     0,     1,    -2,    -2,     1,     1,     2,    -2,     1,     0,    -2,     0,    -1,     0,     1,    -1,    -2,    -2,    -1,     0,     1,     2,    -2,    -3,    -1,    -2,    -3,    -2,    -2,    -1,    -4,    -1,     2,     0,     0,     0,     2,    -1,    -1,     2,     0,    -2,     1,     0,     0,     0,     2,    -2,     0,    -6,    -8,    -3,    -3,   -10,    -9,   -15,     0,    -5,    -3,    -5,    -4,    -9,    -4,    -4,    -5,     0,     2,    -2,    -2,     1,     2,     0,    -2,     1,     1,     1,    -1,    -1,     0,     1,     1,    -1,     0,     1,    -3,    -6,    -5,    -3,    -6,    -2,    -1,    -2,    -6,    -8,    -5,    -1,     0,    -1,    -1,     0,     8,    -2,    -2,    -1,    -1,    -2,     0,     0,     0,    -4,    -4,    -2,    -3,     0,    -1,    -6,    -4,    -6,    -4,    -1,     0,   -17,    -8,    -5,     1,     0,     0,     0,     3,     8,    -1,     2,    -2,    -5,    -9,    -7,    -8,   -10,    -3,    -9,    -3,     1,     6,     8,     5,     0,    -4,    -6,    -5,    -4,   -14,    -4,     0,    -1,    -1,     6,    -2,     6,     6,     2,     2,    -1,     2,     3,     2,     4,    -3,    -4,    -4,    -8,   -11,     1,     2,    -3,   -10,    -8,    -6,    -1,    -1,    -9,    -2,     0,     2,    11,     1,    -3,     6,     1,     6,     6,     7,     2,     6,     0,    -7,    -5,    -9,    -8,    -4,    -8,   -17,   -10,    -7,    -7,    -7,    -5,    -3,   -14,    -3,    -2,     4,     9,     8,     5,    -1,     7,     8,     7,    -4,     2,    -5,    -8,    -1,     3,     4,    -1,     5,     1,     0,    -8,    -5,    -3,    -2,    -3,    -7,   -12,     0,     2,   -10,    22,     5,     6,     0,    11,     4,     0,     6,     5,   -10,    -7,     1,     7,    -1,   -14,     2,     6,    -1,     0,     5,    -6,     0,   -12,   -13,    -6,     0,     2,    -9,    19,     6,    -3,    -6,     6,     0,    -6,   -12,    -9,    -8,     0,     1,    10,   -10,   -13,    -3,     3,    -3,     3,     4,    -1,    -2,   -11,    -5,    -1,    -1,     1,    -1,    -8,    -7,    -3,    -7,   -12,   -10,   -12,   -14,    -6,     0,     3,    -5,    -9,    -9,    -2,    -1,     3,     1,     2,     4,     4,    -3,    -5,   -11,    -4,     0,     2,     0,   -10,    -4,    -4,   -12,   -15,    -1,    -3,    -4,    -2,     0,    -6,   -18,    -8,    -1,    -1,     5,     6,    -2,    -1,     1,     0,    -4,    -4,     2,     0,    -2,     1,     1,    -6,    -4,    -1,    -6,    -9,     0,     2,     3,    -6,     1,    -5,     4,    -2,    -2,    -4,     6,    -3,    -4,    -8,     0,     2,    -4,    -6,    -5,    -6,    -5,    -1,     7,    -3,    -5,     1,    -1,    -4,    -9,    -5,    -6,     0,    -2,    -7,     2,     7,     4,     2,    -7,   -11,    -7,   -10,    -4,    -4,    -2,    -4,   -14,    -7,    -5,    -1,     3,    -2,    -6,     5,    -6,    -6,    -3,     0,    -4,     0,     0,     2,     3,     4,    -4,     1,    -1,    -7,   -10,    -5,    -5,     5,     0,    -4,     0,    -2,     0,    -1,     0,    -3,    -4,     1,    -6,    -1,    -5,    -2,     9,     2,    -2,    -2,     1,     1,    -4,     0,   -10,    -1,     0,    -3,    -1,     5,     0,    -3,     2,   -10,    -7,    -2,     3,    -2,     8,     1,    -2,    -1,    -3,     0,     7,    -2,     4,     3,    -2,    -4,     1,    -3,   -11,   -10,    -6,    -3,     0,     5,    -1,    -6,    -3,    -1,    -3,    -4,     1,     1,     6,     6,     5,     0,    -8,     0,     6,    12,    -2,     2,     9,    -2,    -4,    -5,   -11,   -11,    -5,    -2,     5,     8,     2,    -5,    -4,    -2,    -5,    -2,    -1,     2,     2,     8,     5,     2,    -3,    -2,    -1,     5,    -4,     4,     1,    -6,    -4,    -7,    -6,    -6,    -6,     3,     3,    11,     9,    -6,    -3,    -4,    -4,    -1,     1,    -2,     3,     3,     3,     5,    -3,    -6,     2,    -1,   -14,    -1,     7,     0,    -7,    -2,    -4,    -6,     1,    -3,     4,    10,     8,    -9,    -7,     0,    -3,     0,     0,     1,     4,     5,     1,    -1,    -9,   -12,    -2,    -6,   -13,   -13,    -8,   -11,    -3,     4,    -5,    -1,     1,    -1,     1,     0,     8,    -6,    -7,     0,     2,    -3,     0,     1,     3,     9,     2,     0,    -5,   -13,    -7,    -5,   -14,   -19,   -11,   -17,   -12,    -5,    -4,     9,    11,     5,    -5,    -1,     8,    -3,    -6,    -2,     2,     1,     2,     5,    -3,    -2,    -3,    -2,    -3,    -8,   -14,    -4,    -3,   -10,    -9,   -11,    -2,     8,     3,     5,    -5,     1,     2,     4,     1,    -5,    -7,     2,    -2,    -1,     0,    -5,     0,    -4,    -4,    -3,     4,    -8,   -10,   -12,    -2,   -14,    -5,     7,    16,    10,     0,    -5,    -3,     1,    -2,    -6,     4,   -10,    -5,    -3,    -1,     0,     0,     4,    -4,   -11,   -12,    -4,     2,     7,     0,    -4,    -4,     3,    16,    22,     3,     7,    -5,    -1,     1,     6,     0,    -9,   -23,    -2,     0,     0,     1,     0,     1,    -1,    -8,    -9,    -9,   -14,   -10,   -10,   -15,    -8,    -7,     8,    15,    11,    -2,    -5,    -5,    -4,    -5,    -8,    -6,   -12,     2,     2,     0,    -1,     2,     0,     2,     0,     2,     1,     0,    -3,     2,     2,    -8,    -8,    -3,    -5,    -5,    -4,    -9,     0,     1,    -3,    -2,    -5,    -5,    -1,    -1,     1,     1,     2,     0),
		    34 => (   -2,    -1,    -1,     1,     0,     0,    -2,     2,    -1,     2,    -2,    -1,     0,    -2,     1,     2,     1,     2,     0,     1,    -1,    -1,    -1,     0,     2,    -2,    -1,     2,    -2,    -2,     2,     2,     1,     0,    -2,    -5,    -5,     1,    -2,     1,     1,    -9,    -8,    -2,    -1,    -4,     0,     1,    -1,    -2,    -3,    -2,     0,    -2,    -1,     0,     2,    -2,    -2,    -2,    -6,     1,    -4,    -8,    -3,    -2,    -4,    -4,    -2,    -6,    -7,    -3,    -2,    -7,    -1,    -1,    -7,    -3,    -3,    -2,     1,     0,     0,     2,     2,    -2,    -1,    -2,    -3,    -3,   -11,    -6,    -9,    -5,    -2,    -3,    -4,    -9,   -14,   -14,    -9,     3,    -1,    -6,    -3,     0,    -2,    -2,     0,    -3,     0,    -1,     1,    -1,     0,    -3,    -5,    -1,    -5,    -4,    -2,    -3,    -4,    -5,    -6,   -12,   -17,    -9,    -5,    -5,   -13,   -11,    -2,    -8,   -10,    -2,     3,    -1,    -2,    -3,     1,     2,     2,    -3,    -4,    -1,    -5,    -2,    -6,    -8,    -2,   -10,   -16,   -10,     0,     6,    -3,   -21,   -18,     1,    -6,    -3,    -4,     7,     8,     1,    -7,    -2,    -1,     0,     2,    -6,    -4,     8,    -6,    -1,    -6,    -6,   -10,    -6,    -3,     0,    15,     1,   -31,   -37,   -12,     2,    14,     0,     9,    -8,     3,    -3,     8,   -13,    -2,   -14,     0,    -2,    -3,    12,    -2,    -2,     2,    -6,   -16,    -9,     6,     5,     6,   -25,   -33,   -25,    -4,     7,     3,    -2,     8,     5,     3,     3,     0,    -7,    -5,   -12,     3,    -2,    -2,     2,     2,     7,    -1,    -5,   -17,     2,     8,     9,   -11,   -14,   -28,    -7,     2,     1,     3,    -1,     8,     2,     6,    -1,    -5,   -10,     2,   -10,     4,    -2,     1,    -5,    -8,    -3,    -8,   -12,   -10,    12,     1,    -1,    -7,   -25,   -19,    -2,     4,     7,     4,     1,     3,     1,     2,    -5,    -1,    -5,    -2,    -2,    -8,    -1,    -1,   -12,   -10,    -2,   -10,   -11,    -2,    12,     0,    -8,   -16,    -8,    -5,    -4,    -3,     1,    -2,   -12,   -18,     1,   -12,    -1,    -4,    -4,    -2,    -1,    -8,    -5,    -8,    -9,    -5,   -11,    -2,    -4,     3,     6,     0,    -6,    -1,     7,    -4,     1,     0,     9,    -5,    -5,   -10,   -12,    -8,    -4,    -9,   -12,     2,     0,   -14,   -10,   -15,    -7,   -11,    -6,    -7,     1,     5,    -3,     1,     0,     3,    -3,     1,    -3,    -4,     2,    -3,     5,    -5,   -11,    -7,    -7,   -19,   -13,    -2,    -2,   -10,    -9,   -16,    -8,     0,    -4,     0,     1,    15,     4,    -4,     4,     6,     6,     7,    -3,    -9,     6,     6,     3,   -10,   -13,   -12,   -16,   -19,    -2,    -1,    -2,    -7,   -15,   -15,    -6,    -7,    -2,    -7,     1,     6,    -1,    -3,     3,    -2,     8,     7,    -8,     1,     5,    13,     5,   -10,    -3,    -8,    -8,    -9,    -1,    -1,     0,    -4,    -3,     2,    -7,   -10,     1,    -2,     2,    -2,    -4,    -2,    -2,    -1,    12,    -6,    -1,    -5,    10,    -8,     2,    -1,     4,    -8,    -5,    -3,     4,    -2,     2,    -4,     0,    -1,     3,    -7,     0,     5,     7,    -6,    -7,    -3,     3,     1,    -2,    -6,   -10,   -18,    -6,    -9,    -8,    -6,     2,     2,     0,    -3,    -2,     2,     1,    -8,    -2,    -5,    -6,     1,    -5,     5,    -2,   -10,    -3,    -6,    -8,    -5,    -1,     6,   -12,   -14,   -11,    -8,    -2,    -3,     4,    -1,     1,     0,    -4,    -3,     2,    -8,     3,     6,     0,    -3,    -1,   -13,   -14,   -11,    -1,    -5,    -5,    -2,    -3,     0,   -12,     0,    -1,     3,     0,    -4,     0,    -1,    -2,     1,    -2,     1,    -9,   -10,     3,    10,    -5,   -13,   -11,   -13,    -8,   -14,     0,     0,    -4,    -3,    -2,     0,    -8,    -2,     4,     0,    -6,    -8,     0,    -2,     2,     1,    -3,     0,    -2,    -2,    -4,     2,    -8,   -19,   -11,   -18,    -6,    -5,     4,    -6,    -7,    -9,   -15,    -6,   -11,    -6,    -5,    -6,    -6,    -2,     3,     2,    -6,    -3,     1,     1,     2,    -5,    -8,    -1,    -7,   -24,   -15,    -2,     0,     0,    -4,     0,    -4,    -8,   -10,   -18,   -10,     1,     1,    -5,    -9,     5,     3,     4,   -14,    -4,     1,    -2,     2,     2,    -6,    -7,     0,    -9,   -12,     1,     1,     4,     9,     2,    -4,   -12,    -5,    -9,    -5,     3,    -8,    -5,    -1,     2,     1,     2,     0,     1,    -2,    -2,     2,    -5,    -4,    -4,   -10,    -7,    -8,     3,    -4,     3,     0,    -8,   -15,    -9,    -3,    -5,    -3,    11,     7,   -11,    -1,     2,     7,     4,     2,     1,     0,     2,     2,     0,    -3,   -11,    -6,    -1,    -2,     3,     3,     8,     4,   -11,    -1,    -2,     5,     0,    -5,    13,    11,     7,     4,     6,     5,    -2,    11,    -1,     2,     0,     0,    -6,     1,    -9,    -2,   -11,    -6,   -11,    -9,     2,     1,     4,     3,     1,    -5,    -9,    -1,     9,    11,     3,     2,     9,     3,     4,    -2,    -2,     2,     1,     0,     1,    -2,    -9,    -2,    -6,    -7,    -8,   -10,     2,    -4,     4,    -3,   -12,    -5,    -2,    -5,   -12,    -6,    -6,   -19,   -17,    -1,    -4,     0,     0,    -2,     2,    -1,    -1,     2,     1,     0,    -4,    -1,    -1,    -4,   -15,   -15,   -11,    -9,   -12,    -1,    -6,   -13,    -4,    -9,    -6,    -5,    -4,    -3,    -2,     1,     2,    -1),
		    35 => (    2,    -1,     2,     2,     0,     1,    -1,     1,     1,     2,    -2,    -1,    -2,    -2,     2,    -1,     0,     1,     1,     0,    -1,    -1,     0,     1,    -1,     2,     2,     1,    -1,     0,     1,    -1,     1,     0,    -2,    -1,    -1,    -1,     1,    -4,    -3,    -3,    -2,    -5,    -8,    -7,    -3,    -5,    -1,    -3,    -2,    -2,     0,    -1,    -2,    -1,     2,    -2,    -2,    -4,    -4,     2,    -6,    -6,    -5,   -11,   -12,   -10,   -14,   -13,   -30,   -20,   -12,    -6,    -5,     4,     1,   -14,    -6,     2,    -6,    -4,     1,     1,     2,     2,    -1,     1,    -2,   -12,   -10,    -8,   -20,   -21,   -16,    -4,    -5,    -1,    -4,    -5,    -9,     5,    14,     6,    -8,    -4,    -5,    -8,    -8,    -2,     1,    -2,     0,     1,    -4,     3,    -8,    -4,   -13,     1,    -4,    -1,     7,    -4,   -13,    -5,     6,     8,    -3,    -6,     1,    -8,    -9,    -5,   -10,   -15,   -18,   -12,    -4,    -3,    -1,     0,    -3,    -2,    -8,     1,    -7,   -17,   -13,    -7,    -7,    -3,   -13,   -11,    -6,   -12,   -11,   -21,   -22,    -3,     4,    -9,   -10,    -3,   -12,   -15,     5,     3,    -1,    -1,     8,   -11,   -13,     6,    -7,   -10,    -3,    -9,     2,    -4,   -11,    -5,     1,    -6,   -10,    -8,    -3,    -3,    -1,    -2,     0,    -2,     0,   -14,    -2,     1,     2,    -3,     8,    -6,   -15,     6,   -13,    -6,    -2,    -2,    17,     4,    -5,    -1,    -1,     3,   -11,   -11,   -19,   -20,    -6,    -2,     2,     2,    -6,    -3,     0,     9,    -2,     0,   -10,     1,    -5,    -3,    -7,    -1,    -1,     2,     4,     6,    -4,    -4,     6,     5,     7,     5,     0,     8,     8,     9,    13,    13,    12,     8,    -8,     6,    -1,    -1,   -11,    -7,    -5,   -18,     4,     6,    -1,    -2,    -3,    -9,    -5,    -2,     6,     6,    14,    22,    16,    18,    12,    15,    13,     9,    21,    17,   -12,     2,    -1,    -2,    -2,    -8,    -1,    -4,     5,     4,    -4,    -1,     1,    10,    -6,    -1,     2,     4,     2,     8,    18,    16,    16,    20,    14,     6,    23,    17,     8,    12,     2,    -3,    -1,    -2,     4,     0,    -5,   -11,    -4,    -8,     5,    -3,    -5,    -9,   -18,   -15,   -13,   -13,   -10,   -16,   -11,     3,     2,     8,     2,    19,    17,     1,     0,    -3,    -1,     2,    -4,    -6,    -9,    -3,    -1,     6,     8,    12,     6,     0,    -9,   -12,   -19,   -17,   -34,   -55,   -35,   -23,   -24,   -14,   -11,    12,    18,    -6,     0,     0,    -3,     4,    -4,   -12,   -14,     5,     1,    -3,    14,     5,     9,     2,     3,     0,   -10,    -1,   -12,   -23,   -31,   -20,   -27,   -27,   -10,    -4,    12,    -6,     4,     1,    -3,    -4,     6,    -1,     5,     3,    10,     9,    -1,     1,    -2,    -2,    -3,    -1,    -5,     4,     0,   -19,   -21,   -16,   -14,    -9,   -10,   -13,    -4,    -2,     3,     1,   -10,     9,    17,     7,     3,    13,     8,    10,    -2,     1,     4,    -1,    -8,    -9,   -15,    -4,     6,     0,    -9,    -8,   -15,    -6,   -11,     5,    -4,    -7,     0,     1,    -9,     1,     6,    17,    -2,     9,     0,     6,    -1,    -6,    -5,    -2,   -14,    -6,    -9,    -4,     4,     0,    -1,    -7,    -6,    -8,    -5,     5,    -9,   -10,     2,    -2,   -17,     2,     5,     4,     3,    -7,    -4,     4,     2,    -3,   -11,   -11,   -10,    -1,    -5,    -1,    -7,    -1,    -6,   -10,    -4,    -3,   -17,   -19,   -18,   -18,    -4,    -3,   -10,   -18,    -8,    -5,     0,    -5,    -6,   -10,   -19,     8,    10,    -5,   -10,     2,    -8,     1,    -5,     1,     5,   -11,    -2,     9,     2,    -7,   -19,   -12,     1,     0,    -3,   -15,     7,    11,    -4,    -6,    -4,   -14,   -17,   -17,    -1,     7,   -11,    -9,    -4,     3,     2,     8,     1,   -12,     4,    16,    15,    18,   -17,   -13,    -1,     1,    -3,   -10,     8,     0,    -7,    -2,    -7,    -7,    -9,     1,     3,     6,   -21,    -7,     3,     0,     1,     7,     5,    -9,     3,     3,    18,    20,   -14,     0,     0,     2,    -3,    -7,    -4,     5,    -9,    -9,    -3,    -1,     2,     3,     4,     3,    -6,    11,    -3,    -1,    -2,    -1,     3,    -6,   -10,     0,    14,    24,    12,    -2,     0,    -1,    -7,    -2,    -4,     5,     6,    -8,   -13,    -1,     2,     4,     9,     2,     0,     7,     3,     7,     0,    -9,     2,    -2,    -9,    16,    27,    27,    27,     2,    -2,    -1,     8,    -2,     0,     0,    -5,   -12,   -11,     7,    11,    -5,     0,    -7,     3,     4,    -4,    -1,    -1,    -9,     1,    -8,    -1,    26,    27,    24,    32,    -2,     2,    -2,    -2,     0,   -13,   -17,   -13,    -9,    -5,    -7,     2,     4,     9,    -4,     9,    -3,    -3,    -4,    -6,    -5,     1,     7,    18,     9,     7,   -19,    -6,     2,     1,     1,    -1,     1,   -17,   -19,   -11,   -17,   -13,    -7,    -9,     2,    18,     9,    -2,   -11,    -8,    -7,     3,     0,   -10,     8,    10,    13,    14,    -2,    -3,    -2,    -1,     0,    -1,     0,   -10,   -21,   -29,   -27,   -25,   -24,   -21,   -14,   -15,   -23,   -36,    -9,    -2,    -6,    -3,     3,    -1,     4,    -1,   -11,    -6,     1,     2,     0,     1,     1,     2,     1,     0,    -5,    -2,    -6,    -5,    -3,    -2,    -5,    -6,    -4,   -20,   -10,    -4,    -8,   -11,    -7,    -5,    -8,   -19,   -13,    -2,     2,    -1,     0),
		    36 => (    0,     2,     0,     1,     0,    -1,     1,     0,    -2,    -2,    -2,    -1,     3,     2,     0,    -1,     1,    -2,    -1,     2,     1,     1,     1,    -1,    -2,     0,    -2,     0,    -2,    -2,     2,    -2,     1,     2,     8,     8,     8,     6,    12,     2,    -1,     5,    -7,     0,     1,     5,    11,     7,    21,     9,     8,     8,     2,     1,    -1,     2,    -2,     1,     7,     4,    11,     9,    11,    13,     8,    -4,    -6,    -8,   -11,   -11,     2,     6,     9,    18,    10,     5,     3,    20,    18,    14,     9,    13,    -2,    -1,    -1,    -1,   -15,     2,    -5,     7,    13,    13,     1,    -6,    -7,   -19,   -25,    -1,    11,     8,    -9,    -6,     3,    -6,    -6,    -1,   -10,     3,   -15,    -7,   -11,    -2,     1,     1,   -20,    -3,     7,    16,    12,    -5,   -13,   -11,   -14,   -25,   -33,   -14,   -17,    -9,    -1,    -7,    -4,    22,    14,     3,   -17,   -19,   -30,   -22,    -9,     6,     0,     0,    -9,   -12,     6,    13,     6,    -4,    -6,    -5,    -9,   -28,   -19,     1,     3,    -9,    -5,     0,     6,     6,    11,     8,    -6,     1,   -14,   -21,     1,     2,    -2,    -1,     9,     3,     3,    12,    12,    -1,    -4,   -14,   -16,   -11,    -7,    -9,    -7,    11,     8,     2,     1,    -1,     1,     1,     4,    -8,    -6,   -17,    -8,    -2,     0,    -1,    -1,    -4,    -4,     2,    -6,     0,    -9,   -17,   -29,   -22,    -7,    -9,     5,     8,    -8,   -11,    -4,   -20,     2,    -3,     9,   -11,   -25,   -23,    -5,   -10,     0,     0,   -10,    -8,    -5,     2,     8,    -9,   -14,   -27,   -27,    -4,    -1,    -2,    -3,     3,     0,    -9,   -23,     0,    -9,   -11,   -10,   -27,   -23,   -11,    -9,   -13,     1,     0,    -9,    -7,    14,    -4,    -2,    -2,   -15,   -14,    -8,    -1,    -4,     3,     8,     4,   -11,   -18,   -24,   -30,   -37,   -35,   -32,   -30,   -23,   -13,   -14,    -4,     2,     1,    -9,    -4,    -9,   -10,   -12,   -11,   -24,    -7,     3,     0,     2,     4,     0,    -2,   -10,    -3,    -5,   -21,   -22,   -21,   -26,   -29,   -21,   -17,   -12,   -10,    -1,     0,     2,   -15,    -6,    -2,    -3,    -6,     3,     0,     3,     4,     7,     6,    -3,   -15,   -13,    -6,   -10,    -3,    -6,   -11,     0,   -25,   -26,   -24,   -16,   -13,     2,    -2,    -3,   -10,   -10,    -3,    -2,   -10,    -1,     2,     9,     7,     3,    15,    -5,     2,   -11,     7,    -2,     0,    -4,    -9,     4,     3,   -10,   -24,   -24,   -12,    -2,     1,    -3,   -13,   -10,    -5,   -10,   -12,     3,     2,     5,    16,     4,     8,     0,     1,    -4,     5,    16,     0,     2,     1,    16,    14,   -14,   -27,   -13,    -1,    -1,     1,    -1,   -15,   -10,     3,   -14,     0,    -5,     6,     9,     3,     0,    -6,    -5,    -1,     0,   -21,     4,     8,    -1,    14,    10,     1,     4,   -10,   -12,     0,     1,     2,     0,   -13,    -2,     3,    -8,     0,     6,     5,     6,   -11,    -4,    -5,     0,   -15,   -12,   -15,     4,    11,     6,    17,     6,     3,   -13,   -18,   -22,   -13,     0,     2,     0,    -5,    -4,     5,    -2,     9,    -3,     6,     1,     7,    11,     8,     7,     0,     4,     0,     1,    -2,     7,    15,     8,    -2,   -17,   -20,   -21,   -16,     0,    -1,    -1,     1,     3,     5,     1,     3,    11,    -1,     4,     7,    -6,     1,    -4,    -7,    -6,    -2,    -1,     1,     6,    13,    -5,    -4,   -16,   -13,     0,   -17,     0,    -3,     1,     0,    12,    -3,    -7,    -4,    -3,    12,     8,    -6,    -4,    -6,    -1,    13,    -2,     6,     9,     5,     3,    -3,   -24,   -19,   -14,   -12,    -2,    -7,     0,    -6,    -7,     3,     9,    -9,    -4,     0,    -7,     3,     6,    10,    -1,   -19,    -7,     5,    -2,    -2,     8,    -5,    -4,    -9,   -26,   -10,    -5,    -5,    -9,    -3,    -2,    -6,    -5,   -15,    10,     4,    -3,    -3,    -3,    -6,     3,    10,     9,    -5,    -2,    -3,   -14,    -9,   -14,    -4,    -1,    -2,    -4,   -12,    -7,    -8,   -11,     2,     1,    -2,    -8,    -7,    -7,    -9,     0,    -3,    -1,     0,    -4,    10,    -5,    -3,    -5,   -13,    -4,    -8,    -5,    -9,    -3,     2,   -10,    -8,    -8,    -8,    -8,    -2,    -2,    -1,    -3,    -5,   -10,   -14,   -15,    -8,   -10,    -5,     1,     2,     5,     7,    -1,     3,    -5,   -11,    -5,    -9,   -17,   -14,    -4,    -9,   -19,    -9,     2,    -3,     0,     2,     2,    -3,    -6,    -9,   -10,   -17,   -11,   -14,     0,     6,     5,    -1,     5,     8,   -10,   -19,    10,    15,     9,    -2,    -1,    -3,    -4,    -2,    -4,    -2,    -2,    -2,     1,     2,    -4,    -1,    -2,    -6,   -10,   -16,   -18,   -18,    -8,    -4,     3,    12,    15,     0,    -2,   -19,   -12,    -4,    -4,     0,    -1,    -1,     2,     2,     1,    -1,     2,     2,     2,    -2,    -6,    -8,    -5,    -2,    -8,     4,    11,     2,    -2,     0,    -3,    -2,     0,    -3,    -8,    -2,     1,     0,    -3,     2,    -1,     2,     1,     0,    -2,    -2,     0,     0,     1,     0,     0,    -1,    -1,    -1,     1,    -2,     0,    -3,    -3,     1,     0,     2,     0,    -4,     0,    -3,     0,    -1,     2,     0,     1,    -1,     2,     0,     0,     1,     2,    -2,     1,     1,    -3,     0,    -2,     0,    -3,     0,     1,    -3,    -3,     1,     1,     1,     1,     0,     2,     0,     2,     0),
		    37 => (    0,    -2,    -1,     1,     1,     1,     1,     0,     0,     1,    -1,    -2,     0,    -1,     2,     0,     1,    -1,    -1,    -2,     1,     1,    -2,     1,     1,     2,    -2,    -2,     0,    -2,     1,     1,    -1,     0,     1,    -1,    -2,    -3,    -1,    -8,   -10,    -7,    -5,    -8,   -10,    -8,    -3,     1,    -1,     0,     2,    -1,     1,     2,    -2,     1,    -2,     1,    -1,    -6,    -6,     0,    -2,    -7,   -12,    -5,    -1,   -11,    -4,    -1,     0,    -1,     0,    -3,    -3,     1,    -1,     0,     1,    -2,     2,     0,     2,     1,    -2,     2,    -2,    -4,    -4,    -3,    -7,   -18,   -17,    -6,   -10,    -8,    -6,    -8,    -4,    -5,    -5,   -12,    -5,    -8,    -3,    -3,    -4,    -1,    -2,     1,    -2,    -1,    -2,     0,     2,    -3,   -12,    -9,    -7,   -11,   -19,   -18,   -18,   -21,   -21,   -10,   -18,   -15,   -10,   -10,   -11,    -3,    -6,    -7,    -8,    -8,    -9,    -3,     1,     2,    -1,     2,     1,   -15,   -23,     3,    -7,     6,    21,     7,   -13,   -19,   -11,     8,    -6,    -3,   -22,   -27,   -19,   -28,   -23,   -12,   -12,   -12,    -3,   -11,    -2,    -2,     1,     1,     4,     4,    -2,     1,    -1,   -10,     0,    -4,   -17,   -10,   -11,   -13,    -5,    -9,   -22,    -2,     6,    -2,     0,    13,     1,   -11,   -17,    -2,   -18,    -5,     1,     3,     3,     7,     7,     2,     6,     9,     1,     0,     2,   -13,    -7,    -4,    -7,   -15,   -13,    -2,     0,   -25,   -14,    -4,    -3,    -7,   -15,    -8,    -8,    -4,    -6,     3,    -9,     2,     8,    10,    16,     6,     2,    14,    -2,     2,     5,     1,   -11,    -7,    -7,    -6,     7,   -12,    -5,     0,    -5,     3,     0,    -8,   -14,    -4,     1,     5,     0,     4,    21,     0,     3,    -1,    -2,     2,   -10,     5,    13,     7,    10,     6,    -8,    -7,    -1,    -5,     2,    10,     9,    18,     3,   -11,    -9,    10,     0,    12,     7,     9,    23,    10,    10,    -8,     1,     7,     0,     8,     2,     0,     8,    10,    -2,    -1,    -3,    -1,    -4,    -3,    20,     7,   -14,    -1,    -7,    10,    -1,     8,    19,    16,    20,     3,    -7,    -1,    -6,    -1,     3,     8,    -1,     3,     3,     4,    -8,    -6,    -5,     2,   -10,     6,     6,    -6,   -22,   -19,    -5,    16,     2,     3,     3,    22,    10,     4,    -3,    -3,    -4,    -4,    -3,     2,     2,    -5,     4,     4,     2,    -7,     5,     3,    -2,     8,    11,   -13,   -11,     5,    -5,    12,     2,     8,     9,    20,     8,     5,    -7,    -6,   -11,    -9,     6,     5,    -3,   -14,     5,   -10,     1,    -3,    -4,    -5,    17,    11,     4,    -3,    -2,    13,    -6,    -6,    -3,     5,    21,    21,    -2,     9,    -6,   -11,    -8,    -2,     9,     7,    -9,   -25,    -5,    -5,    -1,     7,     0,    12,     8,     9,     5,    18,    17,    -8,    -9,    -3,    -1,     2,    12,    10,    -8,     1,     3,     0,    -5,     1,    10,     0,   -13,   -15,    -1,    -9,    -9,     3,     3,    17,     7,     3,    11,     8,     6,   -12,    -6,    -4,     0,     0,     5,     3,    14,     5,    -6,     6,     5,    14,     1,    -3,   -24,   -11,    -8,     1,    -4,     1,     2,     7,     1,    15,    21,    19,     8,   -30,   -13,     1,    -2,    -1,    -5,    -1,     8,     4,    -8,     1,     7,     6,    -9,   -13,   -20,   -18,     6,     5,     2,    -4,    -2,    -4,     5,     8,    21,    10,     0,   -29,    -8,   -19,     9,     2,     7,   -22,     0,     1,    -7,     4,     7,     3,    -8,   -18,   -39,   -15,    11,     8,     2,     0,    -2,    -9,     2,     6,    11,    -3,   -15,    -7,    -1,    -6,     0,     8,    -3,   -20,    -5,     2,     9,     3,     1,    -4,   -24,   -44,   -36,   -11,    14,     1,    -6,     3,    -9,    -4,    -7,   -19,   -28,   -14,   -11,   -12,    -1,    -1,    -1,     5,    -2,    -4,     4,    13,    10,    10,     1,   -24,   -33,   -45,   -12,    -5,     1,     1,    -3,    -6,    -8,   -10,   -12,   -14,   -20,   -19,    -2,   -10,     1,     1,     0,    -2,    -2,    -4,   -11,     8,     3,     4,   -12,   -23,   -28,   -22,     0,   -10,     3,     6,     8,    -8,    -8,    -9,   -13,    -7,   -10,   -18,   -18,    -6,    -2,     1,     0,     1,    -2,    -3,     0,    -1,     3,    -5,   -16,   -15,   -24,   -12,    -4,    -5,     5,     0,     0,     1,     2,     4,     3,    -6,   -10,   -11,    -8,    -7,   -11,     2,    -2,     1,    -5,    -5,     3,     4,    -2,    -6,   -15,   -14,   -21,   -12,     3,    -3,    10,     5,    -1,     1,    13,     1,    -1,    -9,   -11,   -16,     0,    -5,    -8,    -2,    -2,     2,    -3,    -1,     2,    -2,    -1,    -7,   -12,   -14,   -18,    -8,     3,    -6,     0,    -3,    -3,     4,     2,     8,    -1,    -2,    -4,   -16,    -1,     0,    -2,     2,     0,     1,    -5,     0,    -1,    -2,     2,    -3,   -10,   -11,   -21,   -11,   -12,    -7,     8,    -2,     9,     9,     6,     9,     3,     2,     4,   -20,    -1,    -6,     1,    -2,     1,     0,    -2,     0,     1,    -3,    -1,     3,     5,     3,    -4,   -21,   -13,    -7,   -19,    -8,     7,     6,     7,    14,     2,     4,     4,    -4,    -5,     2,     0,    -1,     0,    -3,    -2,     1,     1,     7,    -8,    -7,     1,    10,     9,     0,    -3,   -13,   -16,    -7,     8,    10,     2,   -11,     2,    12,     7,    10,     2,     1,    -1,     1),
		    38 => (   -1,     0,     0,     1,     2,     2,     1,     0,    -1,    -2,    -1,     1,     1,     1,     0,    -1,     1,     2,    -2,     0,    -2,    -1,    -2,     1,    -1,     2,     2,     2,    -2,     2,     0,     2,    -2,     2,    -2,     2,    -2,     1,     1,    -2,     2,    -3,    -4,    -9,   -11,    -6,    -5,     0,    -4,    -2,    -4,    -2,    -2,    -1,    -2,     1,     1,     1,    -4,    -1,     0,    -2,    -1,     0,    -4,    -5,   -10,    -8,     1,    -2,     1,    -6,    -3,    -6,    -3,    -2,    -8,    -9,   -12,    -5,    -1,    -4,     0,    -1,     1,     1,    -4,    -1,    -1,    -9,    -4,   -13,   -12,     1,    -1,    -8,    -8,    -9,     1,     8,     8,     6,     3,    -5,    -6,    -3,    -1,     2,    -2,    -1,    -6,    -1,    -2,    -2,     2,    -5,   -14,    -6,    -1,    -1,     1,    -2,    -4,    -2,    -6,    -9,    -3,     3,     4,     2,     3,     2,    10,     7,    -7,    -4,   -14,    -6,    -2,    -5,    -2,    -1,    -3,   -12,   -14,    -5,    -1,    -4,    -7,   -10,    -8,   -10,   -11,   -11,    -9,     4,    -3,    -3,     5,     6,     7,     1,    -1,    -9,    -5,     0,     0,    -8,    -1,     1,    -5,    -7,    -1,     3,    -6,    -3,    -5,   -10,   -15,   -16,   -13,    -8,     1,     3,     0,     0,    -3,     7,    -5,     8,     2,     1,    -9,    -2,    -2,     0,     2,    -9,    -7,    -4,     3,    -1,    -1,     1,     4,    -2,     3,    -3,    -3,     7,     2,     5,    -1,    -7,    -5,    -1,    -1,    -8,     0,    -3,    -7,     5,     9,     4,    -4,    -6,    -4,     1,     1,     2,     1,     2,    -4,     6,     6,     0,     1,    -1,    14,    12,     3,     1,    -7,     0,    -7,    -4,    -8,    -2,    10,    18,    13,     5,     2,    -5,    -1,     2,    -3,    -5,    -5,    -2,   -11,   -10,    -2,    -7,    -3,    -1,     5,     9,     2,    -9,   -10,     1,    -6,    -2,     3,    11,    12,    12,     4,   -16,     1,    -2,     0,    -1,    -4,    -6,    -7,    -6,    -6,     3,    -6,   -13,   -11,    -7,     1,    -2,    -3,    -5,   -13,    -7,    -2,    12,    11,     4,     0,   -17,    -9,   -15,     0,    -1,    -3,    -1,    -4,    -6,    -8,    -5,    -9,    -2,    -3,   -11,    -6,    -6,     5,    -4,     3,    -8,    -3,     3,    -8,    -2,    12,     0,    -5,   -10,     5,   -10,     2,     1,    -1,    -8,    -3,    -8,    -5,   -11,   -15,    -1,     2,     0,     2,     2,    -2,     5,    -3,     3,     5,     2,     8,     6,    -1,     0,    -1,   -14,    -8,   -16,     0,    -2,    -8,   -13,    -3,    -5,   -15,   -12,    -8,    -6,    -9,    -3,    -5,     3,     1,     1,     5,     9,    -5,    -3,    -9,    -8,     2,    -1,     1,    -7,    -2,     3,    -1,    -1,    -2,   -16,    -6,   -10,     8,     5,    -7,   -20,   -16,     2,    -1,     8,     6,     3,     6,    -8,    -9,   -18,    -5,     2,     1,     3,     0,     1,    -4,    -6,    -2,    -2,     0,    -2,    -4,    -2,    14,     5,    -9,    -9,    -3,     5,     6,     5,     0,    -2,    -2,   -11,   -20,   -10,    -6,    -2,     1,    -8,   -10,     1,    -8,    -5,     2,    -1,    -3,    -5,    -3,     5,     7,     2,     4,    10,     6,     8,     4,    -9,   -14,   -10,    -1,   -15,   -22,   -14,    -9,    -4,    -7,   -12,    -9,     0,   -15,    -7,     2,    -4,    -1,    -3,    -1,     5,    13,    21,    16,    12,     8,     0,   -11,    -7,   -10,    -7,   -13,    -2,   -11,    -8,    -8,   -15,    -8,    -9,    -6,    -3,     1,    -3,     1,    -2,     1,    -2,    -1,     7,    13,    12,    11,     6,    -6,   -11,   -17,     1,     8,    -8,   -11,    -2,     1,    -3,    -8,   -13,   -12,    -5,    -2,    -4,     0,    -7,     0,     1,    -2,    -9,     4,    16,     7,    -3,     2,    -8,   -18,   -10,    -6,     4,     1,    -3,    -8,     2,     4,   -12,    -7,   -13,   -11,    -7,    -2,     0,    -7,    -5,    -1,    -2,    -1,   -10,    -4,    14,    -3,     4,     3,   -10,   -12,    -9,   -11,    -5,    -6,    -4,    -6,    -5,    -6,   -12,   -15,   -12,   -11,    -3,    -4,    -1,    -7,    -1,    -7,    -5,    -4,    -9,    -1,    11,     1,     1,     6,    -8,    -3,     2,    -9,    -8,    -7,   -11,    -9,    -6,   -14,   -18,   -17,   -14,    -5,    -3,    -1,     0,    -7,    -1,    -7,    -5,    -2,    -6,     3,    -1,     1,     2,     7,    -4,    -2,     1,   -11,    -9,    -5,   -12,    -2,    -9,   -11,    -9,   -14,   -12,    -6,    -3,    -5,    -2,    -7,    -1,     0,     1,     1,    -8,    -4,    -7,    -9,     3,     0,     5,     2,    -1,    -5,    -2,    -7,     0,     3,    -7,   -16,   -12,   -13,    -8,    -1,    -3,    -2,    -3,   -12,     0,     0,     1,    -3,    -3,    -9,    -4,     8,    12,    10,    15,     6,     3,     3,    -2,   -10,     2,    -6,    -8,    -8,    -7,    -3,     0,     0,     0,    -5,    -4,    -4,     0,     0,     0,    -3,    -3,    -5,   -10,    -1,     7,     6,     2,    -3,     1,     5,    -4,     6,     1,    -3,    -6,    -3,     0,     1,     1,     2,    -1,     0,    -3,    -6,     1,     0,     0,     1,   -10,    -2,    -8,   -11,   -10,     3,     1,     2,     0,     3,    -5,    -7,    -8,    -1,    -3,    -2,    -2,   -10,    -5,    -6,     1,     1,     2,     2,    -2,    -2,    -1,    -1,    -1,     0,    -5,    -2,    -2,    -2,    -2,    -1,    -1,     1,    -4,     0,    -2,    -1,    -2,    -3,     1,     1,     0,    -2,     2,    -2,     2,    -1,     1),
		    39 => (   -1,    -1,     0,     0,     2,    -2,    -1,    -1,     1,     0,    -2,     1,    -2,    -1,     1,    -2,    -2,    -1,    -2,    -2,    -1,     2,     1,    -2,     0,    -1,    -1,     1,    -2,     2,    -2,    -2,    -1,     1,    -1,    -2,    -1,     1,    -2,    -1,    -9,    -8,     0,    -5,    -5,    -4,    -8,    -4,    -1,    -3,    -2,    -1,    -2,     0,     2,    -1,     2,     0,     2,    -2,     2,     2,     0,    -1,    -3,    -7,    -6,    -6,    -3,     1,    -7,     0,    -1,    -2,     1,     1,    -2,    -4,    -6,     1,    -1,     2,     1,    -1,    -2,     0,     1,    -5,    -4,    -2,    -3,    -5,   -11,   -16,    -9,   -16,    -7,   -10,    -6,    -9,    -5,    -3,    -4,    -4,   -13,    -9,    -3,     1,    -6,    -3,     1,    -2,     2,     2,     0,    -4,    -9,   -12,   -22,    -3,   -10,   -10,     0,    -3,    -6,   -12,   -15,   -18,    -9,   -10,    -3,    -5,    -6,    -2,    -3,    -1,    -2,   -15,    -2,     1,     2,     2,     2,    -2,     0,    -2,    -8,    -8,   -14,     3,     8,     1,    -1,     6,    -9,   -15,    -7,   -12,   -23,   -10,    -9,   -13,    -3,    -5,    -2,    -5,    -4,     0,    -2,     1,    -1,    -8,   -10,   -19,     2,    -6,     7,     8,    11,     4,     1,    15,     1,   -10,   -16,   -11,   -21,    -8,   -20,    -8,     5,     2,   -11,    -3,    -1,    -2,     2,    -4,   -11,   -10,   -14,   -16,   -12,    -7,     1,    12,     5,     2,     0,     4,    -4,   -16,    -6,   -16,    -7,   -13,   -23,    -8,     4,    -1,    -7,    -5,    -6,    -3,    -6,    -4,   -10,   -10,   -11,    -8,   -10,    -6,    -2,    -5,    -2,    -8,     1,     5,     8,    -5,   -12,    -7,   -14,    -7,   -11,   -13,     1,    -1,    -5,    -7,    -2,     0,     0,    -2,   -14,    -3,    -1,    -4,     3,    12,     5,    -7,   -10,     5,     2,     6,     5,    -4,    -6,    -4,    -8,   -14,    -8,   -16,    -9,    -9,   -13,   -12,    -3,    -2,     0,    -6,   -10,     0,    13,    -5,     8,     0,     5,    -8,    -2,    -2,    -5,    -3,    -7,     4,     2,    -4,    -2,   -13,   -10,    -3,   -23,   -25,   -13,    -9,     0,    -7,    -1,   -14,    -6,     8,    -3,    -2,    17,    11,    -7,   -13,    -7,   -10,    -4,     4,     4,     8,     3,     9,    -7,     1,    -4,    -9,   -19,   -14,   -11,   -21,    -2,    -8,    -2,   -13,    -8,     5,    -2,    10,    11,    -6,    -6,    -3,    -9,   -17,    -6,    -3,     7,     6,    -3,     6,     1,    -5,    -1,     5,   -10,    -8,    -2,   -14,   -11,    -5,    -2,   -12,    -5,    -1,    -9,    12,     0,    -2,     1,    -2,     5,   -12,    -6,    -3,     2,    -8,    -4,    -1,     5,    -2,     6,     5,    -2,   -11,     1,   -11,    -6,    -3,    -4,    -3,    -3,    12,     1,     4,     2,    -2,    -3,     9,    10,    11,     2,     4,    -6,   -17,   -10,     2,    10,    -2,    -5,     6,     3,    -2,     5,   -15,    -6,     1,    -2,    -1,    -4,    11,     5,     8,     7,    -9,     3,     3,    -2,     5,    10,   -10,    -3,   -12,   -18,    -5,     5,     3,     4,    -2,    -3,     0,     4,   -15,   -10,    -6,    -2,    -2,    -9,     3,    14,   -10,     7,    -3,    -2,    -5,    -4,    -3,     2,    -5,   -14,   -17,   -12,     1,    12,    11,    -3,    -3,   -10,    -2,     7,     0,    -8,   -14,     2,    -2,    -8,     2,     3,    -5,     2,    -7,     0,    -4,    -2,     1,     5,     5,    -6,    -7,    -3,     5,    -1,    10,    -3,    -5,   -17,    -5,    -6,   -12,   -10,   -12,    -2,     1,    -8,     3,    -6,     6,     6,     4,    -5,     0,     5,     9,    -1,    -1,     8,    10,     7,    -7,     2,     5,     5,   -17,   -11,    -7,    -5,   -11,   -13,    -9,     1,    -1,    -7,    -1,    -6,    -4,     3,     7,    -1,     7,     6,     6,    14,     8,     2,     0,     0,   -14,   -10,     3,     3,    -5,    -5,     3,     1,   -15,   -10,    -4,    -2,    -4,    -4,    -2,     3,    -2,   -12,   -13,     3,    -8,     1,    -9,   -11,    -9,    -8,   -15,   -14,   -15,    -4,    12,     3,    -4,    -5,     4,    18,     1,   -16,     0,     2,    -1,    -8,    -2,     2,    -2,    -3,   -14,   -24,   -24,    -9,    -7,   -12,   -12,   -17,   -18,   -22,   -12,    -7,     9,     2,     0,    -6,     1,    11,    -8,   -21,    -1,    -3,     0,    -9,     6,    -3,    -4,    -4,    -6,   -15,   -19,    -6,     7,    -3,     6,    -2,   -12,    -5,   -11,    -1,     2,     5,    -2,     2,     1,     8,   -14,   -10,    -2,     1,    -2,    -1,     9,     3,     2,    -4,    -6,    -9,   -10,    -6,    -7,     1,     4,     1,    -2,    -9,    -6,    -3,    -5,     4,     2,    -3,    13,    15,   -11,    -7,    -1,     1,     1,    -7,    -1,    -2,     1,    -4,    -5,    -7,   -13,    -9,   -10,     0,     0,     1,    -7,    -4,    -1,     5,    10,    19,     4,    14,    22,     5,     5,     0,    -2,     1,    -1,     8,    -4,    -5,     3,    -2,    -7,    -9,    -8,    -2,     2,    -1,     3,   -14,   -17,   -17,   -14,    -3,    11,     7,     5,    -1,    -8,    -7,     1,    -3,     1,     1,     2,     2,     5,    -1,     1,     5,     2,     3,     1,     0,    -6,    -4,     5,     4,    -5,   -12,   -10,   -13,   -11,     1,     1,     5,    12,     8,    -2,    -1,     1,     0,    -2,    -2,    -2,    -3,    -5,     2,    -1,     1,    -1,    -2,    -1,     4,     5,     5,    -1,    -6,    -7,     5,     4,    -6,   -13,    -1,    -7,     1,     2,     0,    -2),
		    40 => (   -2,     0,     0,    -2,    -2,     1,     1,    -1,    -2,    -1,     2,    -1,     2,    -1,    -1,     0,     0,     2,    -2,     1,    -1,     0,     1,     2,     1,     1,    -1,     0,    -1,     0,     1,     0,     1,     1,     2,     0,     0,    -2,    -4,     2,     5,    -1,    -1,     4,     7,     7,     0,     0,     2,     1,     0,     2,    -2,    -2,    -1,     0,    -1,     0,     2,     6,     5,    -1,     1,     1,    -7,   -14,   -12,    -8,   -13,   -19,   -15,   -19,    -4,    -9,    -8,   -12,   -12,    -2,   -11,    -6,    -4,    -2,    -1,     1,     1,    -2,    -2,     4,     0,    -4,    -9,    -4,    -5,     0,    -2,    -6,    -6,     0,     0,    -3,    -5,   -10,   -18,   -20,    -4,    -6,   -12,   -10,    -7,    -3,    -9,     0,     2,     0,    -2,    -4,    -1,   -15,   -13,    -6,    -4,     7,    -1,    -5,   -13,    -1,     0,    -4,     3,    -9,   -11,    -7,    -8,    -6,     5,   -12,    -6,    -7,   -11,     0,     0,     1,    -5,     6,    -2,    -7,    -2,     1,     8,    -6,    -2,    -7,    -7,     4,    -2,    -7,    -3,     4,    -1,    -9,   -13,    -9,    -2,    -8,    -5,    -6,   -10,    -9,     2,     1,    -4,    -4,     8,     7,     2,     2,   -15,   -13,    -1,    -5,    -6,     6,    -4,    -8,     3,     4,    -9,     7,    -2,     8,     3,   -16,    -8,   -17,    -9,    -5,     2,    -1,    -4,    -5,     8,     8,     2,    -6,   -18,     2,    -3,    -7,     0,    -4,    -1,     1,     3,     9,    15,    14,     3,     4,     2,     6,   -12,    -7,   -18,     6,    15,    -8,    10,     1,     6,     5,    -4,     1,    -1,     0,    -4,    -4,    13,     0,     6,     4,     6,     8,    11,    -8,     1,     6,     3,     9,   -15,   -20,   -17,    -3,    -1,    -3,    11,    -1,   -14,    -1,    -3,    -5,     3,     1,    -8,    -7,     0,    -5,     6,    -1,    -9,     3,     6,    -3,    14,    -5,    -1,    -2,     1,   -21,   -18,     0,    -1,    -1,    11,     0,    -9,   -11,     0,    -6,    -2,    -2,    -9,   -13,     2,     0,     8,     0,    -3,     4,    -1,    -5,    12,     7,    13,    -3,     0,   -14,   -17,     0,    -2,    23,    -8,    -2,   -11,   -13,     9,    12,     3,     5,    -3,    -3,     3,    -3,     3,    -7,    -8,     3,   -10,    -4,     7,    11,     9,    -8,    -9,   -14,   -14,    -1,     2,     3,    -3,    -3,   -10,    -9,    14,    10,     5,     6,    -1,     3,     1,    -6,   -10,    -8,   -18,   -12,    -4,    -3,     5,    12,     3,     2,    -1,    -4,   -16,     1,     0,     5,     6,     7,    -4,     4,    10,    10,    17,     7,    -3,     3,   -13,   -11,    -5,   -20,   -14,   -17,     5,     1,     3,     8,    11,     8,     2,     8,    -8,    -3,    -1,     2,    -2,     3,     3,    15,    12,    22,    13,     5,     1,     3,    -5,    -2,   -11,   -13,   -20,    -9,    -3,     7,     5,     0,     1,    12,    -3,    -2,   -12,     2,    -1,     1,    -5,    -6,    -1,    10,     1,     9,    19,     8,    -2,    -1,    -5,    -8,   -13,   -13,    -6,   -14,    -3,     0,     7,    12,     9,    17,    12,     2,   -20,    -5,    -1,    -2,    -4,    -9,     8,    -1,    10,    15,     6,     4,     5,    -6,   -11,   -11,   -15,   -13,    -1,    -3,     4,    -9,    -5,    11,     7,     0,     6,    -7,   -22,    14,    -1,    -2,    -6,   -15,     3,    -6,    -2,     2,     9,    11,    -1,   -12,   -19,   -13,    -4,     7,    -1,    -4,    -9,    -8,     3,    -9,    13,    -5,     4,   -11,   -16,    15,     2,     2,    -5,   -15,    -4,   -12,    -3,     9,    20,    12,     4,    -9,   -19,   -10,     7,     3,     0,    -4,     0,    -2,     4,     1,     7,    -8,    -1,    -1,   -10,    -6,     1,     7,    -7,    -6,    -4,    -9,    -6,    -4,    18,     7,     4,   -14,    -7,    -9,    -7,    -4,     1,    -6,    -2,   -10,    13,    -3,     6,    -2,    -1,   -19,    -2,    -1,    -1,     5,   -12,     1,    -3,     2,    -4,    -2,     7,    11,    21,    -8,    -1,    -6,    -4,    -9,    -7,    -6,    -8,    -4,   -11,    -8,    -5,   -15,   -14,   -10,     5,     2,    -1,    -2,   -16,    -7,    -4,     0,    -7,    -8,     4,    -3,    -1,    -7,    -8,   -11,    -8,     0,     4,    -6,   -16,   -11,    -8,    -5,     9,    -5,    -8,    -7,     8,     4,     1,    -2,   -15,    -4,   -14,    -3,     1,     2,    11,     9,     7,    -8,    -3,    -3,    -4,    -2,   -10,   -13,   -10,    -1,    -8,     2,     3,    -5,    -6,     2,     8,     5,     0,     2,    -2,   -18,   -14,    -9,     1,     1,    -1,     4,     6,     7,    -5,     0,    -5,    -5,    -7,    -8,   -16,    -8,   -16,    -4,   -10,    -9,   -11,    -3,    -7,    -1,    -2,    -2,    -2,     2,     2,     7,    -9,   -10,    -2,    10,     7,     7,     8,    -6,    -2,     3,    -9,   -16,   -10,   -11,    -9,   -11,   -14,   -11,    -2,     4,     0,    -1,    -2,     2,    -3,    -2,   -13,   -20,   -17,   -14,   -14,   -12,   -18,   -18,   -22,   -11,    -9,   -25,   -25,   -23,   -27,   -19,   -15,   -11,   -10,    -6,    -3,     1,    -1,     0,     1,     2,    -1,    -1,    -5,    -8,   -19,    -9,    -9,   -16,   -17,   -20,   -14,   -13,   -11,   -14,   -10,   -19,   -19,   -12,   -16,   -14,    -6,    -8,     0,    -1,     1,    -2,    -2,    -1,    -1,    -1,     2,    -2,    -2,     2,     0,    -1,     0,     1,    -2,    -8,    -4,    -5,    -5,    -4,    -2,     1,     1,    -8,    -5,    -5,    -1,     0,     1,     1),
		    41 => (    2,    -1,     1,     2,    -2,     0,    -2,    -1,    -2,     1,     1,     1,     0,     1,     0,     2,    -1,     2,    -1,    -1,    -2,     2,     2,     1,    -2,    -1,    -1,    -2,     0,    -2,     0,    -1,     2,    -2,    -1,    -2,     2,     0,    -3,    -2,    -5,    -6,     2,     6,     0,    -5,    -1,     1,     2,     0,     1,    -1,    -1,    -2,    -2,     0,     0,    -2,     2,    -2,     0,    -2,     1,     0,    -4,    -5,    -7,    -5,    -6,    13,    16,    21,    19,    11,    11,    21,    16,   -14,   -15,   -10,     1,     2,     0,     2,     2,    -1,     8,    15,    -1,    -7,   -11,     9,     7,    -2,   -20,   -20,     1,     2,     3,     9,    19,     8,     8,    10,    16,    14,    -8,   -10,    -5,    -4,     2,     2,     2,     1,     2,    10,     1,     3,    -4,   -12,    -9,    -5,     2,    -6,   -14,   -16,     3,    14,    14,     6,    10,     3,     4,     9,    -8,    -7,    -4,   -11,   -10,    -8,    -3,     0,     7,     6,     1,    12,     4,   -13,    -9,   -10,    -5,    -5,   -15,    -8,    -2,     8,    13,     3,     0,    -5,    -5,     8,    -8,    -2,    -5,    -9,    -9,    -5,    -1,    -1,   -10,     1,     1,     3,    -9,   -12,    -6,    -7,   -11,   -10,    -4,     2,     2,     8,    12,    -3,    -3,    -7,    -2,    -6,    -6,     1,     2,     0,    -7,    -6,    -2,    -3,   -13,    -3,    -6,   -17,   -18,    -2,     7,     6,    -6,     1,     1,    -6,    11,     3,     2,     3,   -22,   -12,    -2,    -8,   -11,    -4,    -1,    -1,    -9,    -9,    -2,    -4,   -13,     0,    -7,   -18,    -9,    -8,     3,    23,    -2,    -6,    -4,    -4,     4,     7,    -2,    -5,    -3,   -12,    -1,    -7,    -7,    -5,    -4,    -2,    -9,    -5,     0,     0,   -15,    -3,    -6,   -10,    -1,     3,    11,     8,     3,    -8,    -8,    -4,     5,     8,     7,   -18,    -7,   -19,   -10,   -10,    -5,    -6,    -4,    -4,    -3,    -6,     2,     0,   -15,    -2,   -10,   -16,    -9,     9,    -7,    -8,    -4,    -2,     0,    -7,     0,    -2,     0,     0,    -8,    -8,    -9,   -10,    -4,    -2,    -2,    -4,    -6,     7,    -1,     3,     1,    -2,    -6,    -9,     0,    -5,   -15,     2,    10,    -1,    -1,   -12,     0,    -1,    -3,    -8,   -18,   -10,   -11,    -5,    -7,    -1,    -7,    -3,   -10,     2,    -1,     2,    -1,    -2,    -1,    -4,    -5,    -9,   -11,     8,     0,     9,    -7,   -19,    -1,     0,     3,   -15,    -7,   -15,    -9,    -3,    -5,    -1,    -1,    -2,     1,     2,    -1,     1,     2,     0,    -8,    -4,    -4,    -8,    -3,    11,     3,    -1,    -5,   -32,     1,     5,     1,    -7,   -23,   -14,    -9,   -11,    -7,   -15,   -12,    -1,    -1,    -1,     0,     2,    -1,    -2,    -8,   -10,   -12,   -15,    11,     7,     2,   -12,   -32,   -17,     8,     1,    -5,   -15,   -22,   -17,   -15,   -12,   -12,   -10,    -2,    -4,     5,     1,    -2,     0,     3,     3,   -11,   -13,   -16,   -12,    12,     8,    -9,   -19,   -25,     2,     3,    -2,    -1,   -18,   -24,   -20,   -16,    -9,    -9,   -13,    -9,    -4,    -2,    -6,    -1,     1,     1,    -5,    -8,   -13,    -9,    -7,    -5,    -4,   -29,   -23,   -34,    -3,    -8,   -10,   -15,   -23,   -30,   -19,   -13,   -10,    -8,   -18,     5,    -9,   -11,    -4,     1,     1,    -2,    -8,    -1,     4,    15,    -3,   -10,    -7,    -3,   -19,   -23,    -8,    -2,   -11,    -8,   -13,     2,    10,     4,     1,    -2,   -16,     1,   -21,    -6,    -7,    -1,     0,    -2,    -2,    -6,    14,    -1,    -4,     5,    -4,    -1,   -21,   -24,    -6,     1,    -2,     4,     0,     2,     7,    12,     1,    -4,    -4,     0,    -7,   -12,    -2,     1,    -2,     2,    -4,   -10,    -4,     1,     1,     5,     6,    -3,    -5,   -13,    -3,     0,     2,    12,     1,    -5,     7,    11,    -3,     1,     6,    -2,    -9,   -11,    -8,     0,    -1,     2,    11,    10,   -26,    -4,   -10,    -2,    21,     4,    -2,     0,     6,     8,     6,    12,     5,    14,    11,     7,     4,    18,     9,     1,    -5,    -4,     3,     7,     7,    -3,    16,    14,     7,    -3,     7,     7,     9,    14,    -8,    -4,     7,    -2,    -1,     3,    -3,     6,     2,     9,    11,     1,    -5,     4,     6,    -7,     0,     5,     5,    -7,     9,     6,    22,    14,     2,     5,     5,     0,    -2,     2,    -1,   -12,     0,    -1,    -2,    -2,     0,     5,     8,     8,    11,    12,    11,     5,    -1,     2,    -1,     1,    -3,     0,     6,    16,    -8,   -13,     5,     1,    -6,     0,    -2,     2,     4,     0,    -4,   -14,   -35,   -29,   -21,    -5,   -10,   -11,   -10,     6,     2,     0,    -2,     1,    -4,    -3,    -8,    -5,    -6,    -4,     5,     3,    -4,     2,     0,     4,     0,   -12,   -16,   -10,   -18,   -10,     0,    -8,    -8,   -15,    -4,     3,     1,     1,     1,     0,    -1,     1,     0,    -3,     0,     4,     4,    -2,     0,    -3,   -16,     2,     4,   -10,   -30,     0,    -4,    -9,   -11,   -10,    -7,    -1,     1,     2,     2,     2,     0,     1,     1,    -5,    -8,    -3,    -2,    -7,    -7,    -1,     0,   -17,   -16,     2,     7,     8,    -9,    -2,     1,     1,    -3,    -2,     2,     2,     0,    -1,    -1,     1,     2,     2,     2,     0,    -1,     0,     0,     3,    -2,    -6,    -6,    -2,    -5,     2,    -5,    -8,    -1,    -1,     0,     0,     2,     1,     2,    -2,    -1,     0,     2),
		    42 => (   -2,    -2,     2,     1,    -2,    -1,     1,    -2,     2,     1,    -1,     1,    -3,    -3,     3,     4,     0,     1,     0,    -2,    -1,     1,     0,    -1,    -2,     0,    -1,    -1,     1,    -1,    -1,     2,    -1,    -1,     0,     0,     2,     0,    -6,    -5,    -5,     1,    -6,    -6,     2,     1,    -2,   -17,    -6,    -5,    -4,     1,    -2,    -2,     0,     0,     2,     0,    -2,    -6,    -4,    -1,    -1,    -3,    -2,     0,    11,    13,     1,     3,     7,     7,    12,    14,     4,    -1,     0,    -4,    -6,    -4,     1,     2,    -2,     0,    -2,     1,    -1,    -9,   -11,    -5,    -2,    -6,     6,     6,    15,     1,    -4,    -2,    -5,    -2,     3,    13,    -9,    -1,    -2,     7,    -1,    -6,    -3,    -4,    -1,     2,     0,    -2,    -5,    -8,     0,    -3,    -5,    -1,    11,    21,     9,    -1,    10,    -4,    -4,    -1,     7,     3,     4,    -3,   -12,    -8,    -3,    -9,   -10,    -7,   -16,    -9,    -2,     0,    -3,     0,    -2,     1,     3,     6,     1,     2,     7,    16,     5,    12,    11,     6,    12,    -3,    -3,     7,     4,     0,   -10,    -9,    -9,    -3,   -22,    -8,     2,     1,     4,    -7,    -3,     7,     8,    14,     6,     3,     6,     4,    -2,    -5,     3,     8,    10,     4,    10,     0,     5,    10,    -6,   -23,   -23,    -2,   -18,    -3,     2,    -1,     8,    -4,    -3,     6,     8,    10,     5,     2,    -5,    -3,     9,     7,    -1,     8,     8,     4,     0,    -6,    -3,     3,   -11,   -13,     1,    10,   -27,   -11,    -6,     9,    10,    -3,    -1,     2,     4,     2,    -5,    -1,    -6,     4,    -5,    -5,    -4,    -9,     2,    -6,    -8,    -4,   -13,    -6,    -2,    15,     7,    -4,   -18,   -11,     1,   -11,    11,     3,     1,     1,     3,     0,     1,     6,     8,     1,    -6,    -8,   -10,    -4,    -4,    -2,   -13,   -10,    -4,     3,    -4,     9,    -2,   -14,    -6,    -4,    -2,    -5,    13,     0,     4,     1,    -1,    -1,    -6,    -1,     2,     4,    14,    -1,    -3,    -1,    -1,     4,    -9,    -8,    -6,    -5,   -12,   -11,    -5,    -8,    -4,    -9,     0,    -6,    -4,    -8,     0,     4,     1,    -3,    -2,   -10,     0,     3,     7,    -9,     0,     5,     1,    -4,   -13,    -2,     4,     0,    -7,     3,    -5,     7,   -11,   -14,     1,    -6,   -15,    -4,     0,    -2,     1,    -6,     6,    15,     8,     4,    10,    -9,     2,     1,    -3,    -2,     0,    11,    -4,     7,    13,     9,    -2,    -1,     0,     0,     0,    -3,    -8,    -9,    -2,    -1,     8,     8,    11,     5,     0,    -5,     0,    -1,     0,    -5,     1,     5,    11,    13,     9,     9,     9,     5,    -5,    -7,    13,     1,    -1,    -8,    -2,    -1,   -11,   -13,     3,    17,    12,     2,    -6,    -3,    -7,    -9,   -12,    -6,    -5,     0,    17,    12,     8,    13,    15,    18,    15,     3,    10,    10,     2,    -5,     9,     3,   -10,    -5,     0,     4,    13,     5,    -7,     4,    -4,   -18,   -15,    -5,    -4,     2,     2,    13,    15,    12,     7,    12,     2,     2,     1,     9,     1,    -1,    10,    -7,   -10,   -10,    -4,     9,     6,     6,     3,     6,    -9,   -12,   -11,     9,     2,     5,    17,    18,    15,    20,    11,    24,     7,    10,    14,     7,     0,    -1,    10,    -2,   -12,    -5,    -6,    -3,     9,    14,    13,     9,     5,    -3,     1,     5,    -8,     0,    13,    22,    12,     4,     4,     4,    -4,    -8,    10,     8,    -1,     0,     1,    -5,    -6,    -4,    -1,     1,     5,    11,    20,     9,    -1,    -4,    -8,    -3,    -1,    11,    19,    24,    18,     6,     3,     5,     6,   -11,    -5,    12,     1,    -4,    -7,    -1,    -3,    -1,    -2,     3,     5,    14,    11,     6,     5,   -14,    -1,     2,     1,    31,    33,    29,    11,     7,     9,     3,     3,   -11,    -1,     8,     0,    -5,     2,     4,     2,   -10,   -12,     1,     7,     2,    10,     8,     9,    -3,    -8,     5,    23,    21,    23,    15,     8,    -1,    -9,     1,    -3,    -2,    -6,     0,    -1,    -1,     8,     0,    12,    -4,   -12,     1,     0,    -6,    -5,     0,     0,     3,    -2,    16,    26,    24,    18,    18,     5,    -3,    -3,    -6,   -11,    -5,     1,     1,    -1,    -2,    -3,     1,    -5,     1,   -10,    -6,    -1,    -6,    -5,    -1,    11,    -2,    -3,    16,    34,    22,    29,    10,     7,    -2,    -2,    -4,     1,     8,    -1,    -1,     0,     2,    -2,    -1,    -6,    -1,    -5,     0,     7,    -7,   -20,   -13,    -1,     2,    13,    27,    37,    30,    23,    11,     0,     7,    -9,    -1,     5,     6,    -9,     2,    -2,     2,    -6,    -9,   -27,   -27,    -8,    -6,    -2,   -18,   -15,    -9,    -7,    12,    17,    13,    27,    26,    19,     5,    -1,     0,    -6,    -4,     6,     0,     4,     2,     2,     2,    -1,    -5,   -11,   -17,    11,     3,    -3,    -7,     0,    13,    20,    24,    27,    25,    18,     8,     9,     5,    -3,    -5,   -16,    -2,     2,     6,     4,     0,    -1,     2,    -1,     0,    -5,   -13,   -19,   -18,   -18,   -19,   -21,   -10,   -15,   -13,   -18,   -13,   -13,   -13,   -12,   -16,    -7,    -6,   -19,     0,    -2,    -1,     2,     2,    -2,     0,     1,     2,    -4,    -2,    -2,    -3,    -3,    -2,    -4,    -4,    -2,    -4,    -5,    -2,    -3,    -3,    -4,    -1,   -11,   -15,    -3,    -3,    -2,     1,    -2,    -1),
		    43 => (   -2,    -1,    -2,     1,    -1,    -1,    -1,     2,     2,     1,    -1,     1,     0,     0,    -3,     0,     1,     0,    -2,     1,     1,     1,     2,     1,    -1,     0,    -2,     0,     1,    -1,    -1,     0,    -2,    -2,     1,     1,    -2,    -2,    -4,    -5,    -4,    -9,    -7,   -16,   -22,   -24,    -9,    -3,     0,    -2,     0,    -2,     2,     0,     0,     1,    -1,     1,     0,    -2,    -4,     1,    -5,    -9,   -16,   -16,    -3,     0,    -2,    -2,     0,     0,     4,    -2,    -9,    -7,   -10,   -12,   -12,   -15,    -5,     0,     0,     0,     0,     0,     0,    -6,    -3,     3,    -1,     4,    10,    -4,     0,     4,    14,    -2,    -1,    15,    16,    12,     5,    -9,     1,    -7,   -12,   -26,   -22,    -9,     2,     0,     0,    11,   -17,     4,     5,    -5,   -12,   -13,     4,     8,    12,    -3,     1,     0,    -2,     2,     8,    -4,    -7,   -12,   -10,    -2,    13,   -13,   -26,   -24,    -6,     0,     0,     1,    -4,     3,    -5,    -1,     4,     5,    -2,     1,    -2,     1,    -1,     5,     2,     5,     7,    -4,   -15,    -2,     7,    -5,    -7,    13,    -3,   -27,   -10,    -1,    -1,     2,   -11,    -5,   -11,     1,    10,     8,     2,     2,    -3,   -12,   -12,     0,     6,     9,     7,    13,     8,     6,     5,    11,     4,     5,    16,   -25,   -21,   -10,     1,    -1,    -3,     2,     2,     0,     1,     4,     0,    -1,    -7,    -4,    -2,     3,     5,     1,    -5,     8,     9,     3,    -5,     3,    -3,    21,     9,   -34,   -19,   -11,    -8,    -3,     5,     8,     2,     0,    -5,     2,    -2,    -5,     4,    -2,    10,     9,    -7,   -11,    -3,     4,     6,    13,     2,    -9,     9,     9,     2,   -37,   -24,    -1,     0,   -14,     0,    -4,     7,    -1,   -10,   -13,   -12,    -1,   -13,    -2,    23,    16,     6,     3,     8,     3,    -2,     3,    10,    -1,    15,    11,   -19,   -29,   -26,   -10,     1,   -14,     3,     5,    -7,    -8,   -16,   -17,   -19,   -19,   -23,    -5,    14,    21,    26,     8,    -7,    -4,    -8,    -6,     1,     5,     2,     5,   -19,   -12,   -19,   -10,    -1,    -8,    -2,    11,     1,    -9,   -22,   -20,    -9,   -15,   -29,    -6,     4,    21,    13,    12,     4,     1,    -1,    -7,    -4,    -7,   -10,   -19,   -48,   -24,   -15,    -2,     1,    -4,     1,     1,    -4,     0,    -9,   -17,    -6,   -26,    -5,   -11,     5,    12,    30,    15,    -3,     6,     6,    -7,     0,    -4,   -29,   -33,   -35,   -18,   -13,    -2,     0,    -2,   -30,    -6,    -8,    -9,    -4,    -8,    -2,   -11,   -13,    -7,     2,     9,    21,     8,    18,     4,     5,     4,     2,    -9,   -20,    -8,   -21,   -21,   -14,    -2,    -3,     7,     1,   -17,   -19,   -12,    -8,   -10,    -8,    -4,   -14,    -4,     0,    10,     8,    12,     5,     0,   -11,    -9,   -10,   -14,    -7,     2,   -17,   -19,   -11,    -3,    -1,     4,     0,   -11,    -3,    -3,     3,    -2,     4,   -17,   -16,     4,    16,    16,    12,    15,    -4,   -16,   -18,    -8,    -5,    -2,     9,     9,     7,   -14,     3,    -7,     0,     2,     5,     9,     2,    -5,     0,     1,     0,    -8,    -3,     8,     6,     3,    12,    -5,   -19,   -11,    -5,    -3,    -9,    -9,    11,     2,     7,   -27,   -18,    -8,     0,     3,     6,     8,     5,   -10,    -4,    -4,   -13,    -9,    -2,    12,     2,     6,    -1,   -13,   -16,   -10,    -9,    -3,   -13,    -3,     1,     1,     1,   -21,    -5,    -7,    -5,     2,     8,    11,     0,    -3,     3,     8,    -7,    -4,     9,    15,     0,     1,    -6,    -7,    -5,     1,    -6,     2,     4,     7,    -6,    -6,   -11,   -18,    -4,   -10,     0,    -8,     6,    19,     9,    13,    -7,     9,    -1,     5,    12,     3,   -11,    -7,   -15,     3,     2,     6,     6,     1,     4,     4,    -9,    -5,    -7,   -14,   -18,   -10,     0,    -7,   -13,     4,    -1,    -9,    -9,     5,     8,     2,     8,     4,   -13,    -4,    -4,     8,     9,     4,    -1,    -3,    -2,     4,    -6,    -1,    -9,   -12,    -3,     0,    -2,    -3,    -8,     4,     1,   -14,     0,    10,    10,    -3,    -8,    -7,    -6,     2,    -3,     1,    -2,     1,    -1,     1,    -7,    -6,     0,    -9,   -22,   -14,    -6,    -2,     0,     0,    -4,     5,   -10,    -6,    11,     1,    -9,    -5,    -3,    -4,    -1,     1,     0,    -1,    -3,     3,    -4,    -4,    -3,     2,     0,   -16,   -20,   -26,    -2,    -1,     0,     1,     5,    15,    -4,     1,    13,     4,     8,     2,    11,     6,    -7,     6,    -9,     0,     8,    -1,     8,    -3,    -6,    -9,   -10,   -13,    13,     2,    -8,     2,     1,    -2,     6,    15,    -3,     0,     4,     1,    -7,    -8,     1,    21,   -12,    -1,    15,    -4,    -3,    -7,     1,     1,    -1,    -2,    -7,    -7,   -14,   -12,    -5,     2,     2,     0,     2,    -8,    -9,    -8,   -12,     3,     5,     1,    18,    17,    26,     8,    -1,    -8,     7,     0,     3,     9,   -11,   -22,   -25,   -28,   -13,    -3,    -4,     1,    -1,     2,     1,    -8,   -18,    -8,   -10,    -4,    -2,    -5,     8,     5,    10,     2,   -15,    -9,    -1,     2,     4,    -8,    -7,   -15,   -20,   -13,    -1,     0,    -2,    -1,    -2,    -1,     1,     2,    -4,    -7,    -5,    -5,    -5,   -14,   -15,   -16,   -13,   -24,   -10,   -11,    -7,    -4,    -4,   -15,   -16,    -7,    -1,     2,    -1,     1,    -1,    -1),
		    44 => (    1,     2,     2,     2,    -2,    -1,     2,     2,     1,     2,     1,     1,     0,     0,    -2,    -2,     0,     0,    -1,     2,     0,     1,    -1,    -1,     2,     2,     1,     2,    -1,     1,     2,    -2,     0,    -2,    -2,    -4,     0,    -2,   -12,    -5,   -17,   -13,    -1,    -8,    -6,    -1,    -2,    -1,    -8,    -1,    -3,    -5,    -2,    -2,     0,     2,    -2,    -2,    -2,   -13,   -13,   -15,    -6,   -11,    -9,    -8,    -4,   -15,     4,     2,    -8,   -18,   -12,   -10,   -10,    -4,    -4,    -6,    -8,    -2,    -1,    -2,     2,    -2,    -2,    -2,     0,   -16,   -25,   -14,   -14,   -13,   -16,   -10,     8,    -6,   -15,   -31,   -18,    -2,    -4,    -1,   -13,   -14,    -3,    -4,   -10,    -5,     0,    -6,    -1,     2,    -2,     1,    -3,   -10,    -5,     3,     4,     1,    -3,     0,   -13,   -23,    -2,     3,   -20,   -26,   -28,   -25,   -14,    -4,    -2,     0,     5,     8,    11,     3,    -7,    -4,     0,     2,    -3,    -2,    -3,     0,    -5,    -4,   -14,   -22,   -18,     1,    14,    -5,   -10,    -4,   -12,   -48,   -25,     3,    11,     4,     1,     1,     1,    -1,    -6,    -4,    -2,    -1,     0,    -9,     7,    24,    -3,   -16,    -9,    -7,   -12,     4,    11,     4,    -8,    -9,   -35,   -37,   -15,    11,     8,     3,     0,     8,    10,   -23,     7,   -20,    -1,   -17,    -2,    -8,     3,    21,   -11,    -6,    -5,    -2,     4,     7,    -1,     7,    -3,   -19,   -41,   -38,    -2,    13,     6,    -4,     1,     6,    -4,    -6,     8,   -21,    -7,   -15,     3,    -5,     0,     5,    -8,     4,    -8,     0,    -7,    -1,     7,     6,     2,   -19,   -49,   -15,     6,     6,     3,    -4,    10,    -9,     1,    14,     6,   -13,     1,   -13,     2,    -7,    -3,     4,    -7,    -5,    -5,     2,    -1,     1,    12,    12,     8,   -25,   -25,     7,    12,     5,     6,     4,     5,     4,    13,   -13,   -12,    -8,     2,    -8,   -12,     3,     7,    12,     1,    -7,    -1,     4,    -4,    -4,    -2,    16,    -6,   -27,   -18,     4,    13,    11,     1,    -2,     5,     8,     4,   -23,    -7,    -2,    -2,    -5,    -6,   -16,    -7,     5,    13,    -2,     6,    -5,     3,    -1,    12,    -6,   -18,   -27,   -16,    -6,     2,     2,   -12,     9,     0,    -3,     9,   -11,   -11,    -9,    -2,     0,   -12,   -15,   -21,    -6,     3,    10,     8,    -8,    -3,     8,    11,     6,   -23,   -13,    -3,    -2,    -4,     8,     0,    11,     3,     9,   -14,   -12,   -23,   -13,     1,    -4,   -13,   -15,   -17,    -9,    -3,    -3,     5,     5,     8,    11,     3,     4,     1,     3,     4,     8,    -6,     8,     7,     4,    -2,    -5,   -23,   -19,   -18,     0,    -2,    -2,    -3,   -16,   -12,    -1,    -2,     0,    -3,     7,     2,     8,     2,    -3,     8,     2,    -1,     1,    -4,     7,     3,    -5,    -6,    -3,   -11,   -13,   -15,     0,    -1,    -1,    -2,     5,    -1,     0,     0,    -2,     6,     2,     7,     6,     0,     3,     5,     1,    -4,    -2,     0,    13,   -24,    -7,    -4,    -3,   -12,   -18,   -13,    -1,    -1,    -2,    -6,     4,     0,    -4,   -17,    -1,     2,     1,     0,     0,    -3,     0,    -7,     1,    -3,    -5,    -4,    -5,   -18,   -10,    -6,   -10,   -14,   -20,   -19,    -4,    -1,     0,    -8,     4,    10,    -2,   -12,    -6,    -8,    -4,    -4,    -4,    -1,     0,    -3,     1,    -7,     3,    -3,   -13,   -20,     3,    -4,    -4,   -15,     1,    -3,    -5,    -9,     2,   -10,    17,    22,   -10,    -6,   -12,    -9,   -11,   -22,    -1,    -8,     1,     2,    -2,     3,   -10,     0,    -5,     2,     9,     4,     5,     0,     8,    -1,    -2,    -1,   -11,    -5,    14,     7,   -10,   -14,    -8,    -5,   -12,   -13,    -3,   -11,     1,    -2,    -6,    -1,     2,    -4,    -5,    -3,     4,     3,     4,     9,     6,    -2,    -5,     2,     0,    -4,   -17,   -16,   -19,   -16,   -10,   -13,     0,    -7,    -7,   -10,     0,    -3,    -6,     3,    -2,    -6,    -6,   -17,   -14,   -10,    -5,   -15,   -23,    -4,     1,     1,     0,    -4,   -10,   -17,    20,    -2,     3,    13,    16,    -5,    -2,     1,    -2,    -5,    -4,    -2,   -17,   -14,     2,     2,    -2,     2,     6,    -8,   -30,   -10,    -2,    -2,     2,     1,   -11,   -19,    11,    13,     8,     7,     0,     8,     1,     0,    -1,    -6,    -3,     1,    -7,   -13,    -6,     0,     2,    -1,     8,   -10,    -9,     4,     2,     2,     1,     0,   -11,   -16,   -32,     5,     8,     6,     6,     4,    -1,     5,    -3,     3,     4,    10,    -7,    -6,    -4,    -2,     5,     2,     5,    -6,     2,     6,     2,     1,     1,    -1,    -4,   -25,   -21,    -3,   -10,     0,     4,     6,    -3,     2,     0,    -1,     9,     4,   -11,   -27,    -6,    -5,     7,     4,     7,   -10,    11,    -8,    -2,     2,    -2,    -4,    -1,     0,   -15,   -13,     0,    -2,    -8,     0,     2,     4,     7,     1,    -9,   -10,   -23,   -14,   -10,    -2,    -4,     6,    14,    -3,    -6,    -1,     0,     1,    -1,    -1,   -12,     1,   -14,   -13,   -22,   -11,   -13,   -14,   -10,   -18,   -26,   -30,   -40,    -8,   -11,   -17,    -8,   -10,   -11,    -8,     6,     0,    -2,    -1,    -1,     0,    -1,     0,     1,     2,     0,    -7,   -10,    -9,    -7,   -14,   -16,    -2,    -9,   -14,    -1,   -11,   -15,    -8,    -7,     1,    -2,     1,     0,    -1,     2,     2,     1),
		    45 => (    0,    -2,    -1,     0,    -2,    -2,     0,    -2,     2,    -2,     1,     2,     1,    -1,    -2,     1,    -2,    -2,     2,     1,     0,    -1,    -1,     0,    -1,    -1,     2,    -2,     0,     0,     1,     0,     0,    -2,    -2,     0,     2,     0,    -2,    -5,    -4,    -5,    -7,   -10,   -11,    -9,   -13,   -12,   -12,   -10,    -1,     0,     1,    -1,    -2,     2,    -1,    -1,    -4,    -5,    -5,    -1,    -2,    -2,   -13,    -3,    -7,    -5,    -9,   -12,   -13,   -12,    -3,    -7,    -8,    -8,    -7,   -10,   -10,     6,   -17,    -2,    -1,    -2,     2,     0,    -2,    11,    23,    -4,   -10,   -11,    -3,     5,    -4,   -15,   -13,   -20,   -17,    -8,     6,     1,     2,    -2,     1,     4,   -16,   -13,     0,    20,    18,     1,     1,     2,    -7,    19,    -1,    -1,   -11,   -10,    -9,    -2,    -1,   -18,   -20,   -14,   -10,    -7,   -13,   -12,    -1,    12,    -1,     0,   -12,     1,    15,    13,     1,    -5,     2,     0,   -13,    20,    -5,    -4,    -6,   -12,   -11,    -5,     1,     0,   -16,    -6,    -5,    -3,    -7,    -3,    -2,     8,     2,    -3,    -6,    -4,    -6,     4,    -1,    -5,    -1,     0,   -10,    -3,    -6,    -5,    -7,   -13,    -7,    -2,    -2,   -11,    -1,     1,    -3,     1,    -2,    -9,    -1,    -5,    -6,   -10,    16,    12,     8,    16,    18,     1,     1,    -3,     2,    -5,    -4,   -10,    -7,    -9,     2,    -4,    -1,    -1,     6,     7,     7,     4,     8,    11,    -2,    -8,    -1,     6,     5,     7,     4,    -1,    21,     5,    -6,    -2,   -11,    -3,    -5,    -8,    -5,    -4,    -4,     0,     1,    -3,    -3,     1,     7,    -2,    -3,     2,     2,    18,    21,    10,    15,    12,     4,    -3,     7,    10,     2,    -4,   -20,   -15,    -7,    -7,   -10,    -5,    -3,    -6,    -7,    -1,     5,     0,     4,     0,    -1,     3,    -5,   -11,     7,     3,     6,    10,    26,    21,     4,     5,     0,    -2,    -9,   -10,   -11,     6,    -5,     0,     2,    -6,    -8,    -1,     8,    -1,    -1,     4,     9,   -12,   -41,   -43,   -24,   -21,   -22,    -8,     0,     5,     3,     8,     0,     2,     0,     9,     4,     5,    -4,    -5,    -9,   -18,    -4,   -11,   -13,    -9,     1,    -2,     2,    -3,   -22,   -25,   -37,   -34,   -35,   -27,   -22,    -5,    -1,    -5,     1,     0,    -1,    11,     5,    -2,   -13,   -17,   -15,   -11,    -3,   -11,   -15,    -1,     7,    -3,    -5,     4,     0,    -4,   -16,   -29,   -25,   -45,   -29,   -14,    -2,    -8,    -1,    -2,     0,    14,    -2,    -6,    -4,    -6,    -9,    -1,    -5,     0,    10,     2,     4,     5,    -2,     3,     7,    13,     8,     9,    -1,   -17,   -24,    -7,     1,    -9,     3,     0,    -4,     8,   -10,   -15,    -1,   -10,   -12,    -3,     0,     6,    -2,     1,     2,     9,     8,    -8,     0,     4,    12,    -3,     0,    11,     5,    -7,    -4,    -8,     2,    -1,    -9,     1,    -8,     0,     6,    -2,    -5,   -13,    -4,    -6,    -6,     7,     1,   -10,    -6,    -1,    -5,    -4,    12,    -1,    -3,     9,    16,     0,    -1,    -2,    -2,    -7,   -19,     1,     3,   -13,    13,     3,     1,   -19,   -16,   -17,   -11,    -4,    -2,    -7,     6,     4,     0,    -1,    14,    10,     0,    -8,     2,     6,    -4,    -4,    -2,    -8,   -23,    -8,    10,    -3,    11,    21,     9,     1,     2,   -12,   -22,   -10,   -12,   -10,     0,     0,    -2,    -6,     8,     0,   -18,   -14,    -3,    -3,    -7,    -4,    -2,    -1,   -18,    -1,     2,     4,     6,    17,    10,     2,     4,    -6,    -1,    -7,     0,     0,    -1,     1,    -6,    -8,    -6,    -4,    -9,   -18,   -12,    -5,   -14,   -13,     1,    -3,    15,   -16,    -6,    -3,     7,    13,     9,    14,     6,    10,    10,     8,     4,    -1,    -4,    -6,     4,     6,    -4,    -7,    -9,   -12,    -8,    -6,    -8,   -10,     2,    -3,    12,   -21,   -14,    -1,     0,    -9,     3,     5,     7,     5,     5,    -1,     2,     0,    -2,    -1,    -1,    -5,    -4,    -8,    -4,    -4,    -4,    -4,    -2,    -2,    -2,     1,    -7,     0,    -9,     6,    -5,    -2,   -13,    -9,    -6,     5,    -5,    -3,     4,     0,     4,     3,     3,    -6,   -10,     0,    -2,    -3,    -4,    -4,    -2,    -2,    -1,    -1,   -20,     6,     8,    -1,   -10,     1,   -13,    -6,    -5,    -2,     0,    -4,     3,     2,     0,     0,    -1,    -8,    -1,     6,     2,    -1,    -3,    -2,    -1,     2,     1,    -2,     2,     4,    12,    15,     2,    -8,   -11,   -10,    -1,    -1,    -9,   -12,    -1,    -6,     0,     7,     9,     1,     0,     6,     4,    -1,    -9,    -4,    -3,    -2,    -1,     1,    -9,     0,    -3,    -3,   -11,   -21,   -18,    -7,   -21,   -25,    -9,    -3,    -7,   -10,   -13,    -9,     2,     7,     6,    -1,     5,     1,     3,   -12,    -5,    -1,     1,     2,     0,     4,    -8,    -5,     1,    -5,   -13,    -3,   -23,   -22,     2,    -6,    -7,    -3,    -1,    -3,    -2,    -2,    -3,    -8,     3,     1,     2,     1,    -3,    -2,     2,     2,     2,    -3,    -4,    -5,    -9,    -5,    -7,    -5,    -4,    -5,    -4,     8,    18,    17,    14,     7,    -1,    10,     1,    -5,     0,    -2,    -2,     2,     2,     0,    -1,    -2,     2,     2,    -1,    -3,    -1,     1,    -1,     0,     1,    -1,    -1,     0,    -2,     0,     0,     1,    -5,    -5,    -4,    -4,   -13,    -2,     0,     0,     2,    -2),
		    46 => (   -1,     1,    -2,    -1,    -2,    -1,     0,    -1,    -2,     0,     2,    -1,     1,     1,    -2,     2,     0,     1,    -2,     2,    -1,    -2,    -2,    -2,     2,     0,     2,     1,    -1,     1,     0,    -1,    -1,     0,     7,    10,    13,    14,     7,     5,     2,     5,     4,     2,     0,    -1,     3,     3,    17,     5,     3,     5,    -1,     1,    -1,     0,     0,    -1,     2,     2,     3,     1,    10,    14,    15,     7,    -5,    -4,    -4,     0,    -2,    -1,    -3,    -6,    -2,     9,     8,     3,     3,     9,     8,     3,    -2,     0,     1,    -1,   -11,    -8,     1,     2,     6,    11,     4,     8,     1,   -10,   -12,    -4,    -2,    -2,    -1,    -2,    -2,     4,     1,     8,    -1,     9,    11,     0,    -5,    -1,    -1,    -2,    -6,    -3,     1,     3,     3,     1,     2,     3,    -8,    -7,     0,    -6,    -3,     7,     5,     0,    -3,     0,    -2,     5,     0,     4,     3,     1,     5,     7,    -2,     1,     2,    -4,     2,    -5,    -2,     2,     2,    -6,   -10,     2,    -1,    -6,     4,    -4,    -8,     2,     2,     2,     4,     0,     2,     5,     6,     1,    12,     8,     1,     0,     1,    -1,    -3,    -1,    -5,     2,     0,    -4,     2,    -2,     2,    -7,    -7,   -10,   -13,    -1,     3,     5,     6,    10,     7,     5,     0,    -7,     4,     5,    -1,     0,     2,    -4,    -1,    -3,    -6,    -7,     3,     2,     1,    -3,   -11,    -5,     4,     1,    -6,    -3,    -7,    -1,    -1,    -2,    -3,    -2,     5,    -4,     2,     3,     1,     2,    -1,    -8,    -3,     0,    -4,    -8,     3,     3,    -2,   -11,    -7,    -3,    -3,    -7,     4,     6,    -6,    -6,   -10,    -4,   -15,   -12,    -9,    -9,    -3,   -10,     1,     2,    -1,    -2,    -5,   -10,     0,     0,     7,     1,    -4,    -8,    -8,    -8,    -3,     4,     1,    -2,    -7,   -13,   -14,   -11,   -18,   -13,    -4,    -7,     2,    -3,    -1,    -1,     0,    -5,    -2,    -7,     0,    -3,     6,    -8,    -8,   -12,    -6,    -8,    -1,     5,    -1,   -11,   -12,    -6,   -11,    -9,   -12,   -13,    -5,    -4,    -4,    -6,     0,     0,    -1,    -2,    -1,     3,     7,    -1,     2,    -7,   -13,    -8,    -3,     0,     6,    -1,   -12,   -13,   -10,     0,     1,     0,    -3,    -4,     2,    -7,    -5,     0,     2,    -1,     0,    -1,    -7,     4,     2,    -4,    -2,    -5,   -12,    -5,    -5,     3,    -3,    -8,    -7,     6,     4,    -1,     3,     5,     4,     3,     4,   -10,   -11,    -2,    -2,     1,    -3,    -2,    -4,     6,    -2,     2,     6,    -9,   -11,    -6,     3,     3,    -9,    -3,     0,    -1,     4,     5,    -2,    -2,     0,     5,     7,    -7,    -7,     1,    -2,    -2,     1,    -1,    -3,    10,    -3,     3,     2,    -8,    -8,     8,     5,    -3,    -8,    -1,     2,     9,     9,     8,    -1,    -8,    -2,     5,     6,    -3,    -5,    -6,     1,     2,    -3,    -3,    -2,     6,    -2,     0,     0,    -3,    -9,    -2,    -5,   -10,    -4,     4,     8,     7,     8,    10,    -2,    -4,    -3,     7,     8,    -5,    -6,   -11,    -2,     2,    -2,    -5,    -1,     3,    -3,    -9,     2,    -5,    -5,    -4,    -9,    -2,     3,     2,     4,     8,     1,    -6,    -1,    -3,    -1,     1,     0,    -3,    -5,    -9,    -1,     1,    -5,    -1,    -1,    -7,     0,   -10,     3,    -1,    -3,   -14,   -13,    -1,     5,     1,    -1,     1,    -2,    -5,     6,     5,    -1,    -2,     0,     1,    -4,   -10,     0,    -1,    -4,     0,    -3,    -7,   -11,    -5,     6,     4,    -3,    -7,    -4,     4,     0,     3,    -1,    -6,    -4,    -4,     7,    -1,     0,    -6,    -5,     0,   -11,    -8,    -1,    -2,     0,     0,    -1,    -7,    -1,    -2,    -2,     1,    -6,     3,     0,    -4,     2,    -6,    -1,    -5,    -1,    -4,     5,    -2,    -2,    -2,    -3,    -4,    -4,     0,     1,    -1,     1,    -6,     2,    -4,    -5,    -2,    -1,    -5,     5,    -1,    -8,    -5,     2,    -3,    -9,    -4,    -2,     2,     6,     4,    -5,    -8,    -2,     3,    -4,    -1,    -2,     2,    -1,    -3,     1,    -5,    -6,     2,    -2,     3,    -2,     0,    -7,    -8,    -3,    -5,    -3,    -5,    -1,     2,     5,    -3,    -9,    -4,    -6,     2,    -2,     0,     0,    -1,     1,    -1,     0,    -1,     4,    -1,     0,    -3,     0,    -5,    -2,    -4,    -7,     0,     1,    -2,    -7,    -4,    -6,    -3,   -10,    -6,    -4,    -5,     3,    -1,    -2,     1,     0,    -4,     1,     0,    -4,    -4,     3,     3,     2,     3,     7,    -6,    -3,    -6,     4,    -2,    -7,   -11,    -6,    -9,    -4,    -3,    -5,     1,    -4,     1,    -2,    -1,    -2,     0,    -3,     0,    -4,    -6,    -4,    -6,    -4,    -1,    -1,    -5,    -5,    -7,     0,     1,    -2,   -10,   -11,    -2,    -2,    -3,    -1,    -2,    -1,     2,     0,     0,     0,    -2,     2,    -1,    -5,    -3,    -2,     1,     1,     0,     0,    -1,     0,    -1,    -3,    -3,     0,     0,    -7,    -2,    -3,    -8,    -2,    -2,     1,     1,    -1,     2,    -1,    -1,    -1,    -2,    -2,    -3,     0,     1,     1,     0,     2,    -2,     1,     0,    -2,    -1,    -2,    -1,    -2,    -5,    -1,     1,     2,     2,     2,     1,     2,     2,     1,     2,     0,     1,     1,     0,     1,    -1,     1,    -3,     1,     1,    -2,    -2,     0,     2,     2,     2,    -1,    -2,     0,     0,    -2,     1,     1,     1),
		    47 => (   -1,    -1,     1,    -2,     1,     0,    -1,     2,     1,     0,     0,     2,    -1,     1,    -2,     0,     1,     0,     0,    -2,    -1,    -2,    -1,     2,    -1,    -1,     2,    -1,    -2,     0,     1,    -2,     2,     2,     2,     0,    -2,     2,    -2,   -13,    -9,   -11,    -3,    -2,    -5,    -4,     1,     1,     2,     1,     1,    -2,     0,    -2,     1,    -1,     2,    -2,    -1,    -1,    -1,    -2,    -1,    -1,     1,    -2,    -3,   -10,   -14,    -9,    -7,    -6,    -3,     1,     0,    -3,    -3,     0,    -3,    -1,    -2,     0,    -2,     2,     0,     0,     2,    -5,    -5,    -2,    -4,    -8,    -7,    -5,     0,    -4,    -7,    -4,     1,   -11,   -11,    -7,    -5,    -2,    -4,    -1,    -9,    -2,    -3,     1,    -1,    -2,     2,    -2,     2,    -2,    -1,    -8,    -9,    -8,   -12,    -5,    -8,   -12,   -14,   -11,    -7,    -9,    -8,   -10,    -6,    -1,    -5,    -4,   -13,    -7,    -5,    -5,    -3,     0,    -1,     2,    -1,    -7,    -5,   -13,   -16,   -10,    -3,    -3,   -12,    -2,     3,     0,    -9,   -20,   -22,   -14,   -20,   -25,   -23,   -14,   -13,   -13,   -10,    -4,     0,     2,    -2,     0,     2,     3,    -6,   -14,   -18,   -23,   -19,   -29,   -24,    -7,     8,     9,     3,    -7,   -14,     4,     7,     0,     5,    19,     5,    10,   -11,    -4,   -11,    -3,    -2,    10,     7,    10,     5,    -3,    10,    -1,    -9,   -25,   -22,   -21,   -16,    -4,    -3,   -13,     0,     0,     5,    -8,   -16,    -8,    -6,    -4,    -3,     2,    -6,    -5,    -6,    12,    -5,    -1,    -2,     1,    10,    10,    -8,   -19,   -19,   -19,   -10,   -15,   -17,   -18,   -12,    -8,     4,    -9,   -10,   -16,    -6,     9,     5,     0,   -18,    -6,    -5,    11,    -6,    -5,     0,     3,    17,    -1,     3,    -6,   -15,    -6,    -9,   -15,    -2,    -3,    -2,     1,     2,    -8,    -7,    14,     9,    19,    12,     4,   -12,     1,    -3,     6,     2,    -3,   -15,    -5,     7,     1,    -9,    -5,     0,    -1,     1,     7,     3,     0,    -4,    10,     7,     6,    -1,    10,     8,    -1,    -9,    -3,   -14,     4,    -1,     3,     2,     1,     0,     3,    -4,    12,    -4,     0,    -1,    17,    12,     8,     9,     0,    -7,    -6,     1,     6,     3,     6,     3,     6,    -3,    -7,    -3,    16,     0,    -1,     4,    10,     8,     9,    -9,     9,    11,     0,     3,    11,    15,     3,    -8,    -8,     7,    11,     2,    -3,    -1,    -4,     8,    -1,    13,    10,    19,    19,     1,     3,     9,    11,     9,     4,     4,   -12,    -4,     1,     8,     3,     1,    -8,    -9,    -9,     5,    -3,    -3,    -1,    11,     6,     9,   -14,    13,    13,     7,    -3,    -4,     9,    16,    12,     3,    20,     1,   -13,     5,     6,    10,    -3,   -19,   -26,    -7,    -7,    -4,    -7,     9,     3,     6,     6,     4,     2,     1,    -4,   -11,    -2,     2,    -2,     0,    16,   -11,     5,    -3,     8,     0,    11,    10,   -10,   -32,   -27,   -15,    -2,    -1,     5,     0,    11,     9,    -1,    -3,   -15,   -13,    -3,    -1,     0,     1,    -3,    -1,     8,    18,     1,     3,     4,    -1,    -1,    -9,   -38,   -44,    -9,    -5,     0,    -2,     1,   -10,     3,     9,     7,     3,   -10,   -17,   -21,     1,    -9,     2,    -1,    10,    -1,    11,    -1,    -3,    -3,    -1,   -10,   -26,   -32,   -26,    -1,    -5,     2,    -8,    -3,    -6,    -8,    11,     7,     3,    -8,   -13,   -15,     2,   -13,     5,     1,     9,   -15,     1,    -3,     0,     8,    -2,   -22,   -32,   -14,    -8,     1,     4,     1,   -14,     0,    -5,    -5,    11,     5,     1,   -12,   -13,     1,     2,     0,    -1,    11,     2,   -16,    -4,    -1,     8,     2,    -8,   -23,   -27,   -10,    -5,    11,     1,    -3,    -2,     6,    -7,     5,    -3,    -7,    -5,   -13,   -11,     3,    -2,     1,    -1,     2,    -1,    -7,    -3,    -4,    -3,    -8,   -11,   -18,   -13,    -3,     3,     1,     3,    -6,   -10,     5,    -3,    -1,    -5,    -2,    -5,    -9,    -8,    -2,     0,    -1,     2,     2,     0,   -11,   -14,    -9,   -15,   -22,   -12,    -9,     2,     5,    -2,     1,    -1,    -7,    -8,    -2,     5,     4,     0,     3,    -4,   -11,    16,     0,    -2,     2,     0,    -1,    -3,   -16,    -7,    -8,   -11,   -16,   -11,     1,    -4,     1,     4,     6,    -3,     5,    -4,    -8,     4,    -8,    12,    -4,     0,   -12,     2,     2,    -1,     0,    -2,    -1,    -3,   -12,     0,     2,   -14,    -7,    -3,    -8,     6,     2,     3,     0,     0,    -8,    -2,     1,    -4,     0,     6,    -9,    -2,   -11,     5,     0,    -2,     2,     0,     0,     0,     3,     6,     1,    -8,     1,    -1,     9,     0,     7,     4,   -13,     6,    -2,    -3,     0,    -7,   -14,     6,     2,    -4,   -15,     2,    -8,     2,     1,     1,     0,    -1,     1,    -4,     5,     4,     3,    -2,    -1,     5,    12,     8,     2,    14,     5,     9,     0,    -4,     3,    -4,     3,     0,   -15,     5,    -3,     2,    -1,     0,     2,    -1,    -3,    -2,    -7,     2,    -7,     0,    -1,   -11,     0,    15,    10,    -3,    -6,     1,     3,    -6,   -10,     1,     6,     3,     3,    -3,    -2,    -2,     1,    -2,    -2,     0,     1,     3,     6,    -3,     4,    10,     9,    -3,     1,     3,     8,    -3,    -6,     4,    10,   -13,    -2,     0,    15,    14,    13,    -2,     0,    -2,     2),
		    48 => (   -2,    -2,     0,    -1,     1,     2,     1,    -2,    -2,    -1,    -1,     2,    -1,    -1,     0,    -2,     2,    -2,     0,    -2,     2,     1,    -2,     1,     0,     1,     2,     2,     2,     0,     0,     2,    -2,    -1,     0,    -2,     0,    -2,     0,    -1,    -1,    -1,    -4,    -2,    -6,    -3,    -4,     0,     2,     0,    -2,    -1,     2,    -1,     1,    -1,     2,     2,     0,     1,     0,     0,    -1,    -2,    -8,    -9,   -14,   -11,     2,     1,     1,    -7,    -7,    -1,    -3,     2,   -10,    -9,    -8,    -4,    -5,    -2,     2,    -1,    -2,    -2,    -2,     1,    -4,    -7,   -11,   -10,    -7,    -7,    -8,     3,     7,     5,     2,    -5,     0,    -3,     9,     3,     1,    -2,    -2,    16,     2,     2,    -4,     2,     2,    -1,     2,    -6,   -10,   -15,   -11,   -12,    -5,     2,    -4,    -3,    -6,    -9,     0,    -8,    -3,    -4,    -7,     8,    20,    23,     6,   -14,   -15,    -5,     7,    -2,     0,     0,    -5,    -4,   -13,    -7,    -6,    -2,    -2,    -6,    -4,     2,     0,    -8,    -1,   -20,   -14,   -10,   -14,     3,    12,    16,     8,    -6,   -10,    -4,     2,    -2,    -1,     0,    -5,   -17,    -3,    -6,    -2,     1,   -10,    -3,    -3,    -3,    -4,    -4,    -5,    -9,    -4,    -3,     1,    -4,    -3,    -1,    -2,    -5,   -12,    -8,     0,     3,     0,    -4,    -3,   -10,    -1,     0,     0,    -2,    -1,    -6,    -6,    -9,   -12,     0,     1,     3,     2,    -7,    -1,    14,     2,     0,     4,    -3,   -12,    -6,     4,     6,     0,    -9,    -3,     4,     3,     3,     3,    -1,    -2,    -7,   -10,   -15,   -13,   -12,    -4,     4,    -5,     5,    -2,    -6,     2,    13,    11,    -2,    -9,     2,     5,    12,     0,    -6,    -8,    -4,     5,     0,     3,     5,    -3,     3,    -1,   -10,   -14,   -22,   -10,    -6,    -5,    -3,    -1,    -2,     1,     6,    -2,    -3,    -3,    -5,    -3,    -1,     2,    -5,   -10,   -10,     1,     6,     0,    -1,    -5,     6,    -3,    -4,   -12,   -15,    -7,    -2,     6,     4,    -3,     8,    10,     1,    -2,    -3,    -4,   -13,    -1,    -5,    -1,     0,    -6,     7,    -5,     1,     4,    -4,     2,     5,     6,    -3,    -3,     0,    -4,   -15,    -3,    10,    -3,     1,     5,    -3,    -9,    -8,   -12,    -7,    -1,    -4,     1,     2,    -6,    -6,    -4,    -2,    -5,    -7,   -12,    -3,     5,    12,     2,    -9,   -13,   -12,    -1,     6,    -6,    -4,     2,     0,    -6,     1,     2,    -4,    -7,    -6,     0,     0,    -8,    -7,   -12,    -4,    -4,    -1,     0,     6,     3,    12,     6,     4,   -11,   -10,     2,    -4,   -18,    -6,    -6,    -4,    -1,    -2,    -9,    -7,     1,    -2,    -2,    -3,    -5,   -10,    -7,    -9,   -17,   -11,     3,    -8,    -3,     4,     3,     6,    -4,    -7,     2,   -10,   -13,   -14,   -13,    -5,   -10,    -7,   -13,    -4,   -15,    -6,    -3,    -1,    -4,     4,     0,    -1,   -13,   -11,   -10,    -8,   -15,    -3,    -4,     7,     6,     6,     4,     0,   -13,   -16,   -12,    -3,    -8,    -5,    -4,    -2,   -11,   -10,    -2,    -3,    -5,     6,    -1,    -6,    -8,   -10,    -2,    -9,    -6,    -2,    -6,     5,    -8,    -3,    -3,     0,   -12,    -6,    -9,     4,    -9,    -7,    -5,    -6,   -13,   -10,    -2,    -3,    -7,     7,    -2,    -7,   -11,   -10,   -20,   -20,    -4,     0,     6,     7,    -9,    -6,   -12,     1,     1,    -8,     5,     6,    12,    -2,    -8,    -1,    -1,    -6,    -4,    -2,    -3,    -3,    -3,    -6,   -14,   -13,   -13,    -8,    -2,     5,    13,    -4,     0,     5,    -5,     8,     2,     2,    -3,     0,     5,    -3,    -6,    -4,    -4,    -4,     1,     2,    -3,    -4,    -2,    -5,   -13,   -11,   -10,    -5,    -5,     1,    12,    -7,    -1,     6,   -10,    11,    10,     3,    -4,    -4,     2,     4,    -8,    -3,    -9,    -4,     2,     2,    -4,    -2,    -8,    -6,   -17,   -13,    -7,    -1,     7,    10,     8,    -6,    -7,     2,   -15,    12,    -6,     7,     3,    -1,    -1,     2,    -4,    -4,   -11,     0,    -4,    -1,    -3,    -2,    -7,    -9,   -19,   -17,    -9,    -4,     6,     7,     2,    -9,    -4,    -1,     0,     0,     0,     7,    -1,     2,     4,     2,   -14,    -3,    -9,     2,    -3,     1,    -4,    -2,    -4,    -9,   -24,   -19,   -17,   -13,     1,     1,    -3,     3,    -6,     2,    -5,   -12,    -5,    -1,     1,    10,     2,    -9,    -8,    -1,    -7,    -3,     1,     2,    -5,    -6,    -2,    -6,   -10,    -8,   -14,   -10,    -3,   -10,    -1,    -3,    -1,     3,    -1,     5,    -6,    -1,    11,     3,     9,    -2,     1,    -2,    -5,     0,    -1,     1,    -1,     0,    -2,    -6,   -14,   -14,   -15,    -7,    -2,    -5,   -10,   -15,   -10,    -5,    10,    -8,     2,     1,    13,    -2,    -5,    -5,    -9,    -4,    -2,    -2,    -2,     0,    -6,    -1,    -6,    -7,    -5,   -14,   -13,   -12,    -8,   -10,    -8,    -9,    -2,    11,    14,     7,     8,     4,     4,    -5,    -2,    -2,    -2,    -1,     0,     2,     0,    -2,     1,    -9,     0,    -5,    -8,    -3,    -2,    -8,   -15,    -8,    -7,   -10,   -17,   -13,    -9,    -4,    -2,   -16,   -18,    -6,    -8,    -3,    -2,    -1,     1,    -2,    -2,    -1,     1,     0,    -2,    -1,    -2,    -2,    -3,    -3,    -3,    -5,     1,     1,    -6,    -4,    -7,    -8,     0,     0,    -1,    -2,     0,    -2,     2,     1,     2,    -1),
		    49 => (   -1,    -1,     1,     0,     1,     1,     2,    -2,    -1,     1,     0,     1,     0,     0,     0,    -1,     1,     2,     1,     1,     2,    -2,    -1,     1,    -2,     2,     0,     2,     1,     0,     1,     1,     0,     0,     2,    -1,    -2,    -2,    -3,    -7,    -6,    -6,    -1,   -18,   -17,   -14,    -5,    -2,     2,    -3,     0,    -2,     2,     0,    -1,    -2,    -2,     1,    -1,    -4,    -3,     0,    -3,    -7,    -7,    -4,    -4,   -11,    -5,    -6,   -14,    -6,   -13,    -3,    -1,    -3,    -9,    -2,    -2,    -6,    -2,     2,     1,     0,    -1,     2,    -1,   -20,    -6,    -6,    -3,   -11,   -12,   -16,   -15,   -15,   -29,   -20,   -23,   -22,   -21,   -10,     3,   -11,   -11,    -8,    -5,    -2,    -4,    -4,    -2,     2,     0,     1,    -6,    -7,    -7,   -15,   -20,   -15,   -11,   -20,   -15,   -27,   -32,    -7,   -19,   -13,    -8,     2,     6,   -34,   -18,   -22,   -13,    -3,    -3,   -14,   -12,    -3,    -2,     2,    -4,    -7,    -1,    -7,   -15,   -13,   -14,   -13,    -8,     2,    -5,     7,    -8,    -3,   -12,   -11,   -10,    -9,    -6,    -7,   -21,   -18,   -11,   -11,    -9,     1,    -2,    -3,    -5,   -18,   -22,   -44,   -22,    -3,     0,    18,     4,     8,    -2,    14,    -2,     2,     3,     7,     9,     0,     6,     5,   -13,   -14,   -21,   -19,   -12,    -8,     2,   -11,   -15,   -19,   -34,   -43,    -3,   -13,    -5,     3,     7,     8,    13,     3,    -4,    10,    -2,     6,     3,     0,    -2,     0,    -7,   -19,   -19,   -16,   -12,    -5,   -19,   -13,   -12,   -12,   -21,    -1,    -2,   -13,     2,    -5,    -3,     0,     0,    -9,    -1,    -7,    -1,    -2,     6,    -6,    -1,     7,    -7,    -8,   -12,   -19,   -17,    -8,    -4,    -7,    -1,    -6,   -20,    -2,    -3,     0,    -5,    -9,    -1,     4,    -1,    -3,    -6,    12,    -4,    -6,    -6,     3,     0,     6,     0,    -3,    -7,   -18,   -18,    -7,    -2,   -13,   -20,    -1,     4,     2,    -8,    -7,    -4,     5,    -3,     5,     4,    -7,    -9,   -10,    -4,     6,    -3,     4,     7,     3,     5,    -4,    -9,    24,   -19,   -13,     1,   -31,     9,    -3,    10,    -3,    -6,    -4,     5,    -3,    12,     2,     2,     3,    -8,    -4,     1,    12,     3,     4,     8,     9,    17,    -9,     2,    24,   -15,   -15,    -3,    -7,     5,     5,    19,     4,     2,     7,     1,    13,    -1,     6,   -13,   -15,     3,     1,     4,    12,    15,    17,     6,    11,    13,    18,   -19,   -37,   -22,    -4,     1,   -14,   -11,     2,    25,    19,     7,    14,    13,     8,     9,     1,     4,     4,     8,     6,    15,     0,     6,    10,    14,    10,    27,     5,   -32,   -20,   -14,     0,    -5,   -12,    -7,     4,    19,    15,     4,     6,    16,     5,    11,    -5,    -7,     4,    -3,     0,    10,     2,     7,    12,    -2,     5,    30,    -2,   -45,   -30,    -3,    -2,    -2,    -2,   -25,     5,    17,     2,    -8,     7,    19,    10,     1,   -11,    -8,     3,    -6,    10,     9,    16,    11,    10,    -5,   -11,    -1,   -11,   -40,   -23,     9,    -4,     2,    -2,   -22,   -13,     3,   -11,    -1,    -2,    -2,   -10,    12,   -10,    -5,    -5,    -5,    -1,    -2,     1,    -2,    -6,    -4,   -19,    -5,   -10,   -34,   -18,    -4,   -12,     2,     0,   -25,    -1,    -9,   -10,    -9,     2,    -1,    -6,    -5,   -15,    -4,    -7,    -7,     4,     2,     5,    -8,   -10,   -10,   -10,   -10,    -8,   -27,    -1,    -4,    -9,    11,    -1,   -24,     3,    -9,   -14,    -7,    -3,     1,    -2,     2,    -3,    -9,   -17,     0,    -4,    -3,    -1,     4,    -2,   -13,     2,    -2,   -21,   -46,    -5,   -12,    -7,     2,    -3,   -13,    16,    -7,   -17,   -14,   -16,   -11,   -12,   -11,    -9,   -13,   -28,    -5,    -2,    -8,    -7,    -4,     5,    -1,    -7,     8,   -11,   -21,    -2,   -10,    -4,     2,     0,   -23,    12,    -7,    14,    -8,   -33,   -26,   -15,   -19,    -4,   -16,   -18,     4,    -6,     2,     2,    -7,     5,   -14,    -9,    -5,    -4,     3,     8,    -6,    -2,    -1,     0,   -23,    15,     4,    14,    -7,   -14,   -15,   -13,   -19,   -16,   -16,    -1,   -20,    -8,     2,    -7,   -12,    -7,   -16,    -4,    -7,   -16,    -8,     6,   -39,    -2,     2,    -3,   -21,    13,   -11,    -5,     3,    10,    11,    -1,     5,    -8,    -3,     0,     1,     4,    -5,    -9,   -12,   -18,    -6,    -3,    -3,   -18,     2,    -6,   -23,    -5,     1,     1,   -16,    11,    -3,    -8,    -7,     3,     0,    -8,     1,    -9,    -7,     0,    -1,   -11,    -9,    -7,    -6,    -4,    -1,     7,     8,    -5,     0,    -1,    -4,     2,     0,     1,   -16,   -17,    -3,     8,   -11,     6,    -4,    -2,     4,     9,    -4,    -7,   -16,    -2,     2,   -10,     2,     5,    -7,     2,    11,    14,     0,    -6,    -8,     0,    -2,     2,    11,   -11,    14,     6,   -19,   -22,    -7,    -4,   -15,   -11,     4,    -2,    15,     0,     7,    12,    11,     7,    17,    20,     4,    -3,    -6,    -1,    -9,     2,     0,     1,     0,     9,    11,     0,     4,     1,     3,     4,    -9,    -2,    11,     3,    16,     3,     7,    17,    22,     6,    16,    15,     9,     9,     9,     2,     2,    -1,    -2,    -1,    -1,     0,   -12,   -14,     5,     3,     7,     5,    -2,     4,     2,    -7,    11,     9,     6,   -20,    -7,    11,     1,   -12,     4,   -12,     2,    -2,     0,     1),
		    50 => (    0,    -1,     1,     2,     2,    -1,     0,     0,     2,     1,    -1,     1,    -1,     2,    -2,     1,     0,    -1,    -1,    -1,    -2,    -2,     2,    -2,     2,     2,     1,    -2,     0,    -2,     2,     2,     2,     1,     1,     2,     2,    -2,    -1,     1,     2,     3,    -1,     1,    -2,    -2,     0,     2,    -2,    -2,     2,    -2,    -2,    -1,     2,     1,     1,    -1,     0,     4,     6,    -4,    -4,    -3,    -5,    -6,    -9,   -15,   -16,   -17,    -9,   -12,    -9,   -10,    -4,     2,     2,     0,   -10,    -2,     1,     1,    -2,     0,     2,    -2,     1,     2,     0,     3,    -6,    -4,   -17,   -16,    -6,     0,     0,     6,    -1,   -13,   -17,    -8,    -5,    -1,    -4,    -2,    -4,    -2,    -1,    -2,    -2,     2,    -2,    -2,    -1,     2,    -4,   -14,     9,    -2,    10,    10,     6,     7,    -3,    -1,    -2,   -11,    -2,     5,     6,     1,   -12,   -16,    -4,    -1,    -2,    -1,    -5,    -1,     1,     2,     0,     4,     2,    -9,     0,    -4,   -14,    -3,     3,     7,     3,     7,     4,    -1,     6,     2,     4,    -3,    -4,    -4,    -1,    -2,    -8,   -10,    -8,   -10,     1,     1,    -7,    -3,     5,    -4,     0,    -6,    -6,    -3,     3,     3,     0,     0,     1,     3,    10,     4,     6,    -4,    -3,   -11,    -4,    16,    10,   -12,   -13,    -3,     1,    -3,    -6,    -4,    -5,     7,     6,     4,    -3,     5,    11,     3,     3,     0,     5,     1,     0,     7,    -1,    -4,   -11,    -9,    -6,     6,     8,    -9,   -10,     4,     3,     0,     2,    -7,    -6,     0,    -1,     1,     9,    10,    -3,    -2,    13,     7,     8,    -5,     2,    -7,    -1,    -6,    -1,    -5,     3,     1,     2,   -10,   -14,    -6,    -1,     0,     0,    -4,   -11,    10,    -9,    -1,    -2,     4,    -1,     0,    -4,    -1,     1,     2,    -7,   -11,    12,    11,    12,     5,     9,     0,    14,   -16,   -13,    -2,     2,    -2,     0,    -4,   -16,     2,     0,    -2,     5,     3,     8,    -2,   -15,    -6,    -2,    -2,    -8,     5,     7,    -4,   -10,    -5,    14,     3,    12,   -10,    -9,    -2,     0,     6,    -7,    -9,   -13,    -1,     2,    -1,     1,     2,     7,   -13,   -14,   -14,   -12,   -15,    -4,    -2,     0,   -11,    -7,   -10,    -7,     2,     8,    -5,    -2,    -2,     3,     1,     1,    -6,    -1,    -9,     3,    -4,     1,    -3,    -9,    -3,   -11,   -10,   -10,   -12,    -8,    -5,   -10,     2,    -3,    -5,    -2,   -14,     2,    -5,   -10,    -4,     0,     5,     2,     2,    12,    -1,     0,    -1,    12,     3,    -8,   -22,   -20,   -29,   -24,   -16,   -12,   -11,    -2,    -8,     0,    -2,     2,    -9,    -1,    -3,    -5,    -4,    -2,     1,    -1,    -7,    -6,    14,     7,    11,     5,     3,    -8,   -29,   -21,   -25,   -10,   -14,   -21,   -16,    -4,     1,    -7,     2,    -5,     6,    13,    -1,   -10,     1,     2,     1,    -1,   -16,     4,    12,    13,    -4,     2,     7,     7,   -17,   -32,   -19,    -6,    -9,   -13,   -12,    -9,    -1,    -3,     4,     2,    -4,     3,     0,    -1,    -8,     2,     0,    -2,   -19,    10,    12,     1,    16,    -8,    -3,     3,    -9,    -8,   -17,    -1,   -10,   -24,   -20,   -16,   -14,     5,    13,     2,    -1,    -2,    -5,    -7,    -1,    -1,     1,    -5,    -3,     7,    10,     6,     1,    -4,    -6,     6,    12,     6,     4,    -6,   -26,   -33,   -18,   -23,   -11,    -4,    -2,    -4,     2,    -7,    -8,   -13,     2,     0,     1,    -3,     6,    -9,     9,    15,    10,     3,     3,    -4,    -4,     1,    -9,   -15,   -21,   -26,   -11,    -5,    -2,    12,     6,     6,     3,     3,    -6,    -9,    -4,     0,     0,     2,     3,     1,     8,    -2,     2,     2,    -4,    -3,    -3,     6,    -4,    -4,   -10,     0,     8,   -11,     0,     6,     9,    10,     0,     1,    -7,    -1,    -3,     0,     1,    -2,     3,    13,    17,    -7,    -1,    -6,   -12,    -9,     2,     5,    -3,    -1,     0,     3,     5,     2,    -2,     5,     6,    -6,    -2,     3,    -8,    -2,    -2,     1,    -4,     0,    12,    18,     4,    11,     3,   -10,    -3,    -7,    -2,    -8,    -3,     8,     8,    -6,    -1,    -1,    -1,     0,     8,    11,    -3,    -3,    -3,     0,     6,     0,    -1,    -2,    -3,     3,     8,     9,    13,     9,    -3,     2,    -4,    -1,     0,     4,     3,     4,     4,     0,    -4,     2,    -2,     5,     3,    -8,     1,     0,     3,     0,    -2,    -2,   -12,   -12,     2,    -5,    -8,     0,    -1,     3,     1,     9,     0,    -3,     7,     0,     9,     1,     0,   -11,   -11,    -5,    -4,   -18,     1,    -4,     0,     1,    -2,    -1,    -3,    -7,     1,     5,     4,    -2,    10,    12,     2,     4,     9,    -7,     5,    -2,    10,     6,     9,   -10,   -12,   -12,    -6,     4,     4,     0,    -2,    -2,    -1,     1,    -1,    -1,    -4,    -3,    -3,    -5,    -1,    -3,   -12,    -9,    -8,   -13,   -20,   -22,   -22,   -28,   -19,   -14,   -17,   -10,    -1,    -5,    -2,     2,     2,     2,    -2,    -2,    -2,    -3,    -5,    -6,    -4,     2,    -6,    -5,    -7,    -3,   -13,   -11,   -20,   -14,   -12,   -17,   -17,   -13,   -15,    -9,   -10,     2,    -2,    -2,    -2,     1,     0,     1,    -2,    -2,    -2,    -2,     1,    -2,    -1,    -1,     0,    -3,     2,    -1,    -1,     0,    -3,    -2,    -3,    -2,   -10,    -9,   -11,    -2,     2,     2,    -2),
		    51 => (   -2,    -2,    -1,    -1,    -1,     2,     1,     0,     1,     1,     1,     0,     1,    -2,     0,     0,     0,    -1,     0,     0,     2,     1,     2,    -1,     2,    -1,    -2,    -1,    -2,     0,     2,    -2,    -2,     0,     2,    -2,    -2,    -2,    -2,    -1,     0,    -2,     4,     2,    -2,    -1,    -3,     1,     0,    -1,     1,     0,     1,    -1,    -2,    -1,     0,    -1,    -1,     0,     1,    -1,    -2,    -1,    -4,    -7,   -15,   -14,   -10,     3,   -11,    -3,    14,     4,   -14,   -14,    -4,    -9,    -7,    -4,    -2,     2,     0,    -2,    -1,    -1,    23,    13,     0,   -10,    -6,    -2,    -6,    -7,   -13,   -20,   -11,    -2,    -9,   -12,    -5,    -6,    -3,    18,    15,   -14,    -3,    -7,    -3,    -2,     2,    -2,     1,     1,    20,    21,    -1,   -11,    -6,    -5,    -6,   -14,   -17,    -7,    -2,    11,    10,     0,   -11,   -18,     9,     4,     6,    -5,    -3,    -5,     0,    -3,    -9,    -8,    -2,     0,    19,    10,     3,    -2,    -1,    -8,   -22,   -25,    -5,     2,    -7,     5,     1,     2,     7,   -14,    -7,    -4,   -11,    -8,    -5,    -1,    -3,    -2,    -8,    -8,     0,    -1,    -8,     2,     1,    -4,    -9,    -1,   -21,   -27,   -14,     0,     4,    13,     5,    -8,     2,   -16,    -5,   -16,   -14,    -4,    -2,     2,     0,     0,    -6,    -6,     1,    -3,    -9,     2,    -1,   -11,   -13,    -5,   -29,   -18,     1,     5,     9,    13,     3,    -4,   -10,   -12,    -5,   -28,   -12,    -7,     0,    -2,    -1,    -4,   -16,    -7,     1,    -3,    -8,     3,    -4,    -8,   -12,   -11,   -28,   -14,     1,     0,     2,     9,    16,     9,   -12,   -10,    -7,   -28,    -8,    -6,     6,     0,    -2,    -1,   -10,    -3,     1,    -4,    -9,    -4,    -3,     1,    -7,    -5,   -15,    -1,     5,    -3,   -13,     0,    17,    13,   -10,   -19,     0,     2,   -11,    -1,     4,    -2,    -8,    -5,    -9,   -14,     0,    -3,    -4,    -3,    -7,    -3,   -14,    -7,    -6,   -14,    12,    -1,    -5,     6,     9,    -2,    -6,   -15,   -12,    -1,    -4,   -19,     2,     7,   -11,    -5,     3,    12,     0,     2,    -1,    -4,    -3,    -8,   -17,    -9,   -16,   -11,    -3,     6,    -6,     1,    14,    -3,     0,   -10,   -15,    -5,     7,    -2,     6,     8,   -10,    -6,    -5,    20,     2,     0,   -19,     7,     1,    -1,    -6,    -6,    -5,    11,     4,    -2,     3,     1,     8,    -6,    -2,   -17,   -18,    -9,    15,     1,     3,    10,   -11,     2,     1,    15,     1,    -1,   -18,     1,     1,    -3,    -2,     4,    12,     8,   -19,     4,     4,    -8,    -5,    -7,    -3,   -10,   -12,     5,    17,    -7,    -8,   -15,   -12,    11,     8,    -2,     0,     0,    -1,     2,    -2,   -10,     1,     6,    -4,    -7,   -17,   -11,     4,    -1,    -2,    -8,     2,     1,     0,     2,     4,    -7,   -14,    -2,    -1,    -3,    12,     2,    -2,     0,     2,     6,     0,   -11,    -9,     0,    -4,    -7,    -7,    15,     9,    12,     5,   -13,     1,    -2,     9,    -4,    11,    -5,   -12,    -4,   -12,    -7,     1,    -6,     1,    -1,     2,    -7,    -1,    -6,    -4,     1,    -4,    -9,    -6,     7,     4,     0,     4,    -9,    -9,    -2,     3,   -10,     2,    -6,    -9,    -9,     0,   -11,     0,    -3,    -1,     2,     1,    -4,    -3,   -12,    -9,   -12,    -4,    -7,    -8,    -5,     2,     2,     2,    -5,    -7,   -10,     2,   -10,   -13,    -8,     5,     6,    -6,   -10,    -3,     2,    -2,     0,    -3,    -2,    -6,     0,    -9,    -4,   -12,    -7,   -25,    -5,    -8,    14,     7,    -1,     2,    -3,     7,   -16,     5,    -2,   -14,   -13,   -12,     1,     0,    10,    -2,    -1,     2,    -2,    -3,    -1,    -3,    -8,     5,   -13,   -13,    -5,    -3,     6,    12,     7,     0,    -9,    -5,   -21,    -6,    -7,   -18,   -11,    -5,     6,     8,    11,     2,     2,     0,    -7,    -6,    -4,    -8,   -15,    -4,    -5,    -4,    -3,    11,     4,     5,     4,     2,    -4,    -5,    -9,     1,   -15,   -23,    -8,     0,    -2,    11,    -2,     4,     3,     2,    -6,    -6,    -3,   -10,   -23,    -1,     0,    -6,     0,     1,     2,    -3,     1,    -4,   -14,    10,    -4,     5,    -5,   -17,   -15,    -7,     4,    -4,    -1,     6,     2,     2,     2,    -4,    -3,    -4,   -19,     2,    -1,    -3,    -8,    -6,    -1,     2,    -3,    -4,    -5,     6,     2,     9,    -1,   -14,    -6,   -12,    10,     8,    -1,     2,     0,    -3,    -7,    -2,     2,     9,    -6,     3,    15,     1,     8,    -2,     1,     0,     1,     3,    14,    12,     4,     8,    -5,    -3,    -8,    -9,    -3,    19,     2,    -2,    -2,    -2,    -3,    -3,    -2,    12,     2,    -2,     2,    10,    14,    -2,   -13,   -12,   -17,   -22,    -8,   -16,   -10,   -10,    -6,   -15,    -1,    -9,    13,    10,     2,     2,    -1,    -2,     0,    -1,    -2,    -1,    -2,    -4,    -7,   -32,   -26,   -18,   -16,    -4,   -20,   -19,   -21,   -18,   -18,   -30,   -12,    -9,    -8,    -1,    -1,    -2,     1,     2,    -2,    -1,    -1,    -7,   -15,   -11,   -10,    -9,    -8,    -6,    -9,   -15,   -16,   -17,   -16,   -12,   -12,    -3,    -7,    -1,    -8,    -1,    -1,    -2,     1,     0,     1,    -2,    -1,     2,     0,    -2,     2,     0,     1,    -2,     2,    -1,    -2,    -1,    -2,    -3,    -3,     0,     0,     1,    -1,     0,     1,     0,     0,    -2,    -2,    -1,    -2),
		    52 => (    1,     1,    -1,    -2,     1,     1,    -2,     2,    -1,     0,     2,     2,    -3,    -3,     2,     5,     1,     2,     2,    -1,     1,    -2,     1,    -2,     1,     2,     1,    -1,     1,    -1,     2,    -3,     2,     2,    -2,    -2,    -1,     2,     2,    -2,     2,     2,    -5,    -3,     3,     3,    -2,   -11,    -5,    -1,     1,     1,     2,     1,     1,     2,    -1,    -1,    -4,    -4,    -4,     2,    -3,    -4,    10,    15,    18,     9,     7,    -5,     0,    -7,   -18,   -13,    -1,     5,     1,     5,    -5,     4,     8,     5,    -2,     1,    -2,    -2,    -4,   -15,   -12,   -14,    -4,    -7,     5,     5,    -2,    -3,    -6,     3,     7,    -3,    -1,    -2,    -3,    12,    -4,    -3,    -4,   -18,    -9,     4,    -5,     0,     0,    -1,    -3,    -4,    11,    -3,    -2,     2,     0,     3,    -4,     0,     7,     3,    -1,     5,    -8,     4,    -9,    -3,     6,   -10,    -5,   -17,   -18,     8,   -13,    -6,    -2,    -2,     0,    -6,     2,   -14,   -16,   -21,   -10,    -2,    10,     1,    -7,     6,     4,     3,    -6,     3,    -2,    -1,     0,     3,    -1,     8,   -14,    15,   -11,    -1,    -1,     0,     0,    15,    12,   -13,   -10,    -5,     5,    10,    10,     1,     2,    11,     3,     0,    -5,     3,     1,    -2,    -4,   -10,    -4,    -2,     1,   -12,   -12,    -2,     1,     0,    -4,    19,    15,    10,    -4,     2,    -3,     1,    -2,     4,     3,     6,     1,     7,     9,     8,     3,     7,    -4,    -7,    12,     1,   -10,   -12,   -10,    -8,    -7,    14,    -2,    14,     9,     8,   -10,    -4,    -5,     7,     0,    -2,    -4,    -7,    -3,     2,     7,    11,    -2,    12,    -8,     0,    11,    10,   -28,   -17,   -12,    -8,     3,    -5,     4,     3,    -4,     3,    -7,    -7,    -4,    10,   -10,     1,     5,   -14,    -4,     2,     6,     3,    -2,    12,     1,    -7,    -7,    10,   -23,   -15,    -7,    -3,     0,     0,     1,     8,   -16,    17,     9,    -1,    -3,     1,    -9,   -11,     0,     6,    -4,    -4,    -3,    -5,    -1,     3,     6,    -1,    -5,    11,    -5,    -5,     2,    -3,     1,    -7,    -2,    10,     2,     4,     8,     1,    -4,   -10,   -22,     0,    -7,   -13,   -15,   -12,     1,    -5,   -12,    -2,    -6,    -1,    -6,     5,    -2,     1,   -11,    -2,    -2,     0,   -14,    -1,     3,   -15,    -6,   -11,   -14,   -10,   -12,   -12,    -5,   -19,   -23,    -6,     0,    -2,   -13,    -3,    -8,    -4,    -2,    -7,    -3,     6,    -1,    -6,    -1,     2,     1,    -2,    -2,    -6,   -22,   -19,   -32,   -19,   -14,   -18,   -24,   -14,   -11,    -5,    -4,   -10,    -9,   -11,    -9,   -11,     4,    -9,    -2,     6,    11,    -5,     2,    -7,    -9,    -3,   -13,   -23,   -25,   -26,   -40,   -25,   -13,   -13,    -4,    -8,     0,    -5,   -14,    -5,    -5,    -4,   -11,   -17,    -2,   -20,    -2,     1,    13,     7,     2,    -7,    -1,    -6,   -24,   -13,   -12,   -17,     3,    -2,    -6,     6,     0,     8,     2,   -12,     2,    -2,   -15,   -17,   -17,   -10,   -19,   -10,     4,    -6,    15,    21,     0,     0,    -9,   -15,   -27,   -10,   -11,    -8,    -4,     4,     5,     5,    -9,     4,     4,    -5,    -8,    -3,    -7,   -15,   -11,    -4,     7,    -6,     6,    14,    19,    13,    -2,    -1,     1,   -11,    -9,   -12,    -1,    -3,    -1,     1,     6,     2,    -8,    14,     9,     0,    -2,    -3,    -2,   -13,    -8,    -5,    -4,    -5,   -11,    25,    14,    12,    -1,    -2,    -4,   -21,    -7,    -6,     7,    10,    -4,    -6,     2,    -1,     5,    -1,    -2,    -3,    -2,     6,    -8,   -10,   -13,     8,    10,     9,    18,    30,    -2,    16,    -1,    -5,     4,   -10,   -13,    -4,    10,     6,    -6,   -10,     5,     3,     1,    19,    16,     5,     8,    -2,    -4,    -8,     1,    10,     4,     9,    -3,     9,     8,    16,     1,    -2,    10,    -1,    -1,    -7,    23,     8,     5,     7,    16,    13,    10,    26,     9,     7,    14,    -1,    -3,    -2,    15,    14,     6,     4,     3,    12,     5,     0,     2,     5,     5,    12,     4,     3,    11,     8,    -3,     7,     5,     6,     1,    19,    15,    12,     8,    10,     5,     7,     8,     7,    12,    25,    12,    12,    12,    -3,     1,    -1,    -1,     0,    -1,    12,    18,     9,     2,    10,     2,     4,     3,     1,     6,     5,    -5,   -11,    -1,   -10,     4,    11,    19,    22,    18,    -2,   -17,    -5,    -2,    -2,     2,   -12,    -6,     3,    13,     7,     5,    12,     5,    16,    12,     9,     3,    -3,   -10,    -7,    -8,     0,     9,    13,    23,    16,    13,     2,    -8,     1,     1,     0,   -13,    -9,    -3,    -7,     1,     7,    17,    -5,     1,     1,    11,    -5,     7,     3,   -12,    -4,    -1,     0,   -14,    -8,    -1,    13,    26,    15,     8,     1,     2,    -1,    -8,    -1,   -10,   -25,    12,    -4,   -13,   -26,   -33,   -10,    -5,    -2,    11,     8,    -8,     3,   -17,   -22,    -2,     3,   -18,    -8,     5,    14,     9,    -1,     2,    -2,    -2,     0,    -9,   -16,   -18,   -11,   -11,   -17,   -29,   -23,   -13,   -15,   -15,    -9,   -22,   -21,   -17,    -2,    -7,    -9,    -6,     1,    -2,     0,    -2,     2,    -2,     2,    -2,     1,    -1,     0,    -3,     0,     2,    -1,    -8,   -13,    -1,    -5,    -1,    -1,     1,    -3,    -2,     1,    -5,    -9,    -4,    -1,    -1,     1,     0,     0),
		    53 => (   -1,    -1,     1,    -1,    -1,    -2,     2,    -3,     1,     1,     0,    -2,    -2,    -2,    -1,    -1,    -2,    -1,    -1,    -1,     2,    -2,    -2,    -1,     2,    -1,     0,     0,    -1,     0,     2,     0,    -1,    -1,     2,    -1,     2,    -2,     1,    -1,    -2,    -2,    -5,    -1,    -6,    -2,     0,    -2,     0,     0,     2,     1,     2,     2,     1,    -2,     2,     2,     1,    -2,     1,     2,     1,     0,   -10,   -12,     8,    10,     7,    -4,   -10,   -10,   -15,   -15,   -10,    -5,    -2,    -7,    -8,   -11,    -3,    -2,    -1,     0,    -1,     0,    -1,    -6,    -2,     0,    -4,     5,     2,    -3,     8,     8,     6,     6,     1,    -6,     4,     8,     9,    -4,    -4,    -6,    -2,   -18,    -8,    -2,    -1,     0,    -2,     4,     1,     0,    -3,     2,     3,     7,     3,    -2,    -5,    -8,   -11,   -12,     0,    -5,    -6,   -15,    -7,     0,   -10,    -8,    10,   -20,   -17,    -9,    -3,    -1,     0,     1,     2,    -4,    -2,     7,    10,    16,     2,   -11,   -16,    -8,    -6,    -7,     0,    -3,    -2,    -2,    -3,     2,    -3,    -7,    -9,    -8,    -7,    -2,    -7,    -2,     0,     4,     0,     5,     2,     0,     2,    -2,   -13,    -9,     8,    -2,     1,    -5,    -7,    -5,    -2,     0,     0,   -10,    -8,    -4,    -3,    -3,    -3,   -16,    -9,    -3,     2,     5,     7,   -10,   -23,    -9,     0,    -7,   -12,    -5,    -5,     2,    -4,     0,     1,     1,    -2,     5,    -1,   -10,     2,    -7,    -2,    -9,    -6,   -13,    -9,    -4,     0,    -2,     6,   -14,   -19,     0,    -6,   -10,    -6,     4,     4,    -3,     1,    -7,     2,    -6,     1,     1,     8,     2,     4,    13,     8,   -18,   -29,   -10,   -13,     0,    -2,   -11,    -9,   -11,     2,     1,     7,    -1,    -3,    -4,     6,     9,    14,     7,     6,    -4,    -7,    -5,    -8,    -5,     9,     5,     5,   -14,   -35,   -14,   -14,    -2,     0,   -12,    -5,     8,     4,     3,    15,     1,    21,    10,    11,     9,     0,    -1,    -2,    -6,   -18,    -1,     7,     8,     5,    -3,     7,    -4,   -33,    -3,   -10,     1,    -1,   -13,    -5,    18,    17,    16,     4,    10,     6,    14,     5,   -10,   -21,   -20,   -17,     6,     4,     5,     8,    11,    16,     3,     4,    -1,   -19,   -18,    -4,    -2,    -1,   -12,   -11,    19,    11,     7,     0,     4,   -12,   -11,   -16,   -36,   -26,    -6,     9,    16,     5,     2,     8,    -1,    -4,    -8,    -6,   -12,     0,     2,     0,     2,     1,    -8,   -24,     8,   -12,    -8,    -6,    -8,   -16,   -33,   -34,   -22,    -4,     6,    12,     2,     3,    -1,    -7,    -9,    -6,    -4,   -18,   -14,    11,    -6,    -6,    -2,    -4,     3,    -4,    -6,   -16,   -19,   -27,   -25,   -25,   -13,    -6,   -10,     5,     9,     5,     4,    -3,     2,   -13,    -8,   -11,    -8,   -19,    -4,    16,    -4,    -9,    -6,    -1,     8,     4,     2,    -5,   -10,   -21,   -28,   -20,    -1,     5,    -4,     6,    13,    22,     0,     7,    -3,    -3,    -1,    -4,     1,    -9,    -5,    12,    -5,    11,     2,     0,     2,     6,    12,     3,    -8,   -11,    -8,   -17,   -11,   -12,   -23,    -3,     2,    -4,   -11,     7,     5,    -7,     1,     2,    14,    -3,   -10,     7,   -13,     5,     1,     0,     1,     3,     3,     1,    -1,    -4,   -11,   -21,   -27,   -34,   -38,   -46,   -37,   -24,   -15,     9,    -2,   -11,     8,     7,    14,     5,   -10,    -4,   -17,    -2,    -1,    -5,     2,    14,     4,    18,     2,    -8,     0,    -3,   -18,   -16,   -25,   -36,   -28,   -17,   -16,    -1,    11,     8,     9,     3,    -2,     6,    -4,   -22,    -6,     1,    -6,     0,    -7,    -9,    -8,     5,     8,     0,     0,    -6,     5,    -3,    -8,    -6,     0,     1,    -5,    -5,     1,    -6,     0,     2,     1,    11,     0,    -7,     4,    -3,    -5,     1,    -2,    -9,    -1,     5,     8,    10,     7,     2,    11,    10,    14,     6,     0,    -5,   -13,    -5,   -10,    -8,     2,     9,    -2,     3,    -8,   -10,    -7,    -2,    -3,    -1,     6,    -4,     1,    -4,     5,     2,    10,    11,     4,     1,     0,     2,    -5,     1,   -10,    -9,   -14,    -3,     4,     7,     0,    -5,    -7,   -12,    -5,    -4,     0,    -2,     1,    -6,     1,     1,    -3,    -6,    -8,    -1,    -2,     2,     1,     3,     3,     4,    -2,    -1,     1,    -1,     9,    -1,     2,   -14,   -12,   -11,    -5,    -3,     2,     0,     1,     7,    10,    11,     8,    -3,    -5,    -3,    -2,   -12,    -5,    -9,    -4,    -4,     7,     2,     6,     7,     0,     3,     6,   -14,   -11,    10,     6,     0,     1,    -1,    -1,    -1,     8,    10,     0,    -9,    -5,     1,     6,     0,     2,     5,     1,     1,    -4,     9,     8,    -5,   -14,    -3,    -5,   -10,   -16,   -10,    -6,    -3,     0,    -1,     2,     0,   -11,    -8,     3,     6,     3,    -6,    -5,   -18,   -15,   -12,   -23,   -15,    -1,     0,   -12,   -12,   -12,    -7,    -8,    -7,   -14,     0,     0,     1,     0,    -2,     0,     1,    -8,   -19,   -17,   -13,   -14,   -19,   -17,   -24,   -20,   -17,    -9,    -7,    -7,   -10,   -25,   -23,   -19,    -1,    -8,    -2,     0,     1,     1,     0,     1,    -1,    -2,    -2,    -2,    -2,    -4,    -3,    -4,    -4,   -12,    -9,   -11,     0,    -8,    -8,   -10,    -8,    -8,    -8,   -11,    -5,    -3,    -2,     0,    -1,    -1,     2,     1),
		    54 => (   -1,    -1,    -1,     2,     1,    -1,     1,     0,    -1,    -3,     1,     0,    -3,    -3,    -3,    -2,     2,    -2,    -2,     0,    -2,    -2,     1,    -2,    -2,    -2,     1,     2,    -1,     2,     2,     2,     2,    -1,   -11,    -9,    -3,     0,    -5,    -1,    -4,     3,     9,    -2,    -2,    -1,    -2,    -1,    -5,    -3,    -3,    -2,    -2,     2,     0,     0,    -2,     0,    -1,    -4,   -15,    -1,    -6,   -11,   -16,    -5,    -3,    -3,    -5,   -10,    -8,   -14,   -19,    -8,    -5,    -2,   -12,   -10,    -1,    -3,    -2,    -7,     0,     0,     0,     0,    -4,    -7,   -12,    -4,    -9,   -11,    -5,    -2,    -6,    -3,     1,    -5,   -10,    -1,     2,     7,    -9,    -7,    -9,    -3,    -5,     0,    -1,    -5,     1,     0,     2,     1,    -4,    -3,    -5,    -7,   -12,     7,    15,     8,    -6,   -18,   -24,   -15,   -12,   -11,   -20,   -25,   -26,   -16,    -7,    -6,     2,    21,    16,     9,   -18,    -3,    -2,    -2,    -6,     2,    -7,    -1,    -6,     5,    22,     6,   -13,   -23,   -16,    -9,    24,    13,    10,    -4,   -24,   -30,   -11,   -10,    -2,     7,     4,    -7,    -3,    -3,     1,     1,    -2,    -9,     9,    12,    -4,     9,    10,    -9,   -27,   -32,    -5,     3,     4,    11,    10,     3,   -23,   -44,   -39,    -4,    13,    14,     9,   -20,     5,   -14,    -1,    -8,     0,    -9,     6,     9,     5,     7,    -2,    -5,   -15,   -10,   -14,    -1,    11,    11,     7,     7,   -33,   -46,   -21,     6,    19,    21,     2,   -25,     1,   -17,    -5,    -8,    -1,   -11,    -1,    11,     7,     8,    -3,    -3,   -11,   -15,   -19,     1,     8,    18,    -6,   -22,   -41,   -21,    -3,    10,     6,    -3,    -2,    -9,     5,   -13,    -1,    -3,    -4,   -12,     3,     1,     7,    16,     0,    -8,   -10,   -19,    -7,    -1,    14,     7,    -3,   -22,   -20,    -8,     7,     8,    -3,     4,    -3,    -6,     5,   -11,     1,    -5,   -11,   -13,    -5,     0,     3,     2,   -13,     4,    -4,   -16,     6,    -1,    12,     4,    -3,   -13,   -13,     0,     5,    -1,     1,    -8,     2,     6,    -2,   -10,    -2,     1,   -11,    -7,    -9,     5,    -3,    -4,     2,     7,    -1,     3,     4,   -12,     1,     1,    -7,   -13,    -9,    -3,     0,     1,     4,     0,    -9,    -1,    -8,   -17,     1,    -1,    -8,   -26,    -8,     6,    -4,     1,     3,     2,     7,   -10,     3,     3,    -2,    -7,    -8,    -7,   -13,     2,     5,     2,     2,   -11,    -2,    -7,   -20,   -14,    -1,     2,    -8,   -18,   -12,    -2,     0,     5,    -1,     6,    16,     0,   -11,     7,   -11,    -8,     5,     0,    -3,     6,     1,     1,     1,    -3,   -12,   -16,   -19,    -1,     2,    -1,    -8,   -16,    -5,     0,     9,     1,     1,     6,     8,     1,     1,     9,     5,    -5,     0,     8,    -4,     1,     2,     6,     6,    -7,    -1,   -11,    -5,     1,    -2,    -1,     0,   -16,    -2,     3,     5,    13,    10,     8,     7,     5,     6,    -1,     4,    -2,    -8,     2,     2,     2,    -5,    -6,     2,     0,    -6,    -8,    -3,     3,     2,    -1,    -2,   -12,    -7,     4,    12,    14,     7,     0,    -7,    -3,    -1,    -2,     1,    10,     5,     2,    -3,     1,     5,    -4,   -10,    -9,    -3,    -6,   -14,    -5,    -1,     1,    -4,    -7,    -4,     1,     4,     1,     8,    -6,    -1,    -6,     1,    -2,     9,     4,     3,    -3,    -5,    -6,    -6,    -3,    -1,    -6,   -13,   -12,    -7,    -6,    -7,    -2,    -1,    11,     9,    -3,    -8,    -9,    -7,     3,   -16,   -16,    -8,     1,     9,    -2,    -5,    -6,    -5,   -10,   -17,    -8,    -9,   -10,    -6,    -9,    -4,    -6,    -2,    -6,    -7,    16,     5,   -22,   -16,    -8,    -4,    -2,   -22,   -13,    -8,   -12,     1,    -3,    -5,    -4,     5,    -8,   -14,   -15,   -13,   -14,    -1,    -7,    -5,    -5,     0,     0,     0,    -7,     0,    -7,    -7,    -8,   -14,     3,   -10,    -1,     1,   -11,    10,     1,    -6,    -1,     9,    -9,   -22,     1,    -5,    -4,     7,   -11,    -3,     2,     1,    -1,    -5,   -20,   -11,     1,   -11,   -15,     3,     5,    -1,     3,    -3,   -19,     0,    -6,    -2,    -5,     2,    -3,   -16,    -2,    -6,     3,     2,   -13,    -6,     1,     0,    -1,     2,   -12,   -11,     2,    -3,     4,     8,    -8,    -3,    -1,    -6,   -11,    -4,    -6,     2,    -7,     2,    11,    -3,     1,     6,    -3,     7,     1,     2,     2,    -2,     0,     0,    -7,    -9,   -17,    -5,     4,     4,     1,    14,     6,     4,   -11,    -8,   -12,   -12,    -9,     1,     4,     8,    -2,    -6,     0,     5,     7,     0,     1,    -1,    -2,     1,     0,   -14,   -13,     6,     4,     4,     2,     2,    13,     9,    -8,    -2,    -2,   -19,     0,     4,     5,    10,     1,    10,     5,    -1,    13,     1,    -1,     1,    -1,    -2,    -2,   -10,   -21,     4,     0,    -1,    -1,     7,     8,   -18,   -27,    -8,     1,   -16,     4,   -10,   -16,     1,     1,     8,     1,    -2,    -4,    -1,     1,     1,    -1,     2,   -11,    -3,   -11,   -14,    -6,    -8,   -10,   -15,   -11,   -13,   -17,    -4,     1,    -4,     3,   -13,   -17,   -17,   -20,   -14,    -1,    -2,     1,     1,     2,    -1,     1,     1,     1,    -1,    -2,    -5,    -6,    -7,    -4,   -12,   -10,    -8,    -9,   -16,    -2,    -7,   -13,   -11,   -10,   -13,    -8,   -10,    -2,     0,     0,     1,     0),
		    55 => (   -2,     0,     1,    -1,     0,     2,     0,     2,    -1,    -2,     2,    -1,     1,    -4,     1,     1,     2,    -2,     0,     0,     2,     1,     2,    -1,     0,    -2,     1,     1,    -1,     0,    -2,     0,     0,     0,     0,    -3,     1,     0,    -2,    -8,    -4,    -3,   -10,   -12,   -11,   -13,    -9,   -10,   -15,   -14,    -5,    -1,     0,     1,    -1,     0,    -2,    -2,    -8,    -8,    -4,    -4,    -8,    -7,   -13,   -20,   -18,   -21,   -25,   -32,   -16,     5,     7,     9,     5,    -4,    -1,   -11,   -12,    -3,   -10,    -8,     2,    -1,     1,     2,    -4,     0,    -3,   -12,   -23,   -15,   -30,     6,    11,    -2,     4,     0,    -8,   -14,   -12,    -1,     7,    15,    -2,    12,     0,   -11,    -6,     7,    20,     0,    -1,    -5,   -10,     0,   -13,    -2,    -1,     3,     0,    -3,     5,    -1,     5,    -6,    -3,    -8,   -13,    -8,     9,   -11,   -10,    -2,    -6,    -5,    20,    13,     3,    -6,    -1,     1,   -10,     0,   -10,    -3,    -8,     1,    -7,     1,     0,    17,    14,    -4,     6,    11,    -2,    -9,   -23,    -4,    -2,     0,     2,    10,     0,    12,     4,    -1,     2,     0,    -1,   -14,   -14,    -7,     0,     6,     6,    -1,     0,    12,    17,     2,     2,    -6,    -9,   -11,   -12,    -2,    -5,    -4,     4,    16,    16,    19,    -2,     2,     2,    -8,     2,   -24,   -22,    -9,     7,    16,    14,    12,    12,     5,    -2,     2,     7,     0,     9,     3,   -13,    -3,     3,     0,     1,     0,     4,     4,    -5,     9,    -2,    -6,   -18,   -31,   -15,    10,     0,   -11,    -2,     4,     5,    -1,    -1,     2,     9,    10,    -1,     6,   -11,   -20,    -5,    -6,     2,    -1,    22,     8,   -16,     4,     0,    -2,   -14,   -22,    -9,     9,     5,   -13,     3,    -7,     2,    17,    10,    15,    21,    13,     1,    -6,   -22,   -24,   -24,   -12,     4,     0,    12,    13,    -8,    -6,     0,    -1,   -18,   -37,    14,    14,     9,     4,    -7,    -5,     7,    13,    24,    17,    16,    18,     1,   -22,   -12,   -16,   -15,    -9,   -31,   -26,    10,    14,    13,    -8,     2,    -4,    -2,    -8,     4,     8,     6,    -3,    -4,    -5,    -1,     5,    11,    12,     4,    13,     6,    -2,    -7,   -19,   -11,    -9,   -31,   -36,    -2,    -2,     6,     2,    -1,    -2,    -3,    -5,    10,     4,     0,     2,     0,    -1,     0,   -11,     2,     2,    -2,     2,    -7,    -9,     0,    -4,   -13,    -4,   -23,   -15,   -35,   -15,    14,   -15,     0,    -1,    -6,    -2,     0,     8,    -6,     0,    -2,    -2,     0,     5,     2,     2,    -2,     3,    -4,   -12,    -1,     6,     2,     2,    -5,   -18,   -29,   -22,     0,   -10,     3,    -2,    -2,     2,   -15,    -2,    -5,    -3,    -7,    -2,    -2,    -6,     0,    -9,     2,    -7,     7,    -1,    -6,     2,     6,    -2,     0,    17,     1,   -14,    -9,    -5,     1,     1,    -8,    -5,     2,     0,    -1,    -2,   -18,   -12,     3,    -1,     1,    -6,    -1,     1,    -4,    -2,     1,    -6,    -9,   -18,    -1,    16,     7,   -14,   -14,   -15,     1,    -5,   -17,    15,     2,     5,   -21,   -30,   -15,   -16,    -8,    14,    -2,    -2,    -3,    -9,    -4,    -9,     0,     5,    -5,    -6,    -1,     7,    -5,   -30,   -18,   -17,    -1,    -4,   -27,    27,     6,     1,    -6,   -27,   -19,   -14,    -6,    -1,   -10,    -6,    -7,    -6,     3,     9,     3,    11,     0,     0,     2,     6,   -17,   -30,   -25,   -25,    -3,     2,   -18,    26,    26,    14,    -2,   -16,   -22,   -30,    -4,   -13,    -8,   -13,    -1,    -1,     6,     7,    -2,    -6,     5,     8,     8,    14,    -2,    -4,   -27,    -8,     0,    -7,    14,     1,    21,    19,     6,   -10,    -4,   -17,    -7,    -9,    -2,    -2,     0,     7,    -5,     4,    14,     0,    16,     1,    10,    15,    16,     9,   -17,   -18,    -2,    -7,    11,    -3,     9,    11,     2,     0,     1,    -3,   -11,     0,    -2,     8,    -3,    -5,     8,    11,     2,    -9,     8,    -3,    19,     8,     8,    15,   -14,     0,    -2,    -3,   -13,   -24,    -2,     9,    -5,    -9,    10,     9,     0,    -4,    -5,    -1,     5,    12,    11,     6,    11,    10,     3,    11,    -2,    13,     5,    21,     8,    -3,    -3,    -1,   -20,    -8,   -15,   -14,    -8,     2,     3,     5,     6,    -2,     0,     4,    -3,     0,     4,     0,     3,    10,    -7,     0,     0,    22,    23,    28,    18,     0,     1,     2,     4,     5,    -7,    -4,     2,    -3,   -12,     1,    -3,    -2,    -5,     4,     4,    -2,     4,     3,     9,     9,    -4,     4,    -6,    16,    15,    19,    13,    -1,     2,    -2,   -13,    -4,   -10,    -6,    -8,     5,     7,    17,    12,    11,    -3,    -7,   -13,     3,    -4,    12,    10,    13,     5,    -7,     4,     0,    18,   -12,    -7,     1,     2,     0,     0,     9,   -19,   -24,    -8,    -4,     3,    -8,   -12,   -12,     1,    -7,   -15,     0,    13,    19,    17,    12,     3,    13,    21,    18,    18,    -7,    -2,    -1,     2,     2,    -2,    -5,    -8,   -18,   -23,   -22,    -8,    -2,     5,     4,     0,    -4,   -20,     6,    -4,     6,     5,    20,     5,    -1,    -5,   -10,    -6,     2,     2,     1,    -1,     2,     2,    -1,    -4,    -4,    -2,    -5,    -5,    -5,     2,     2,     3,     2,   -25,   -19,    -5,    -8,    -6,   -11,   -14,   -16,    -9,    -2,     2,     2,     1,     1),
		    56 => (    0,    -1,     0,    -1,     1,    -1,     2,    -1,    -1,     1,     0,    -2,     4,     5,    -1,     2,    -2,     2,     1,     0,     2,     1,     1,     0,     0,     1,     1,    -1,     2,     1,     0,    -2,    -2,    -2,     5,     6,    12,     7,     5,     4,     2,     8,    -1,    -4,    -3,    -2,     0,     2,    14,     7,     5,     1,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,     8,     0,     4,    13,    11,    10,     6,    -4,    -6,    -6,    -6,    -2,     0,    -2,    -2,     6,     8,    11,     8,    13,     5,     5,    -2,    -2,    -2,    -2,   -11,   -11,    -2,     9,     8,     6,     4,     7,    -2,    -9,   -12,   -23,   -10,    -6,    -1,   -10,     4,    14,     8,     6,     3,    13,     9,     2,    -1,     1,     2,     0,   -13,   -14,    10,    14,     9,     2,    -5,     4,     1,   -12,   -16,   -23,   -15,    -1,    -3,    -7,   -15,     1,     1,    -5,   -10,     1,    10,     8,    16,    17,    -2,     2,    -7,   -13,    20,    12,     5,     3,     3,     1,     0,    -6,    -9,   -17,    -7,     6,    -3,     3,    -6,    -7,    -7,    -3,    -6,     3,     6,     8,    17,    12,    -1,     0,     4,    -3,    15,     4,     8,     3,    17,     7,    -7,   -16,   -17,   -18,    -4,    -5,   -14,    -6,    -1,   -13,    -8,    -1,    -3,    -1,     2,   -10,     4,    20,     0,    -1,     1,    -5,    16,     6,    -3,     9,     7,    10,    -5,   -14,   -19,   -11,     0,   -13,   -17,    -1,    -1,    -2,    -3,    -8,    -9,   -11,   -10,    -4,     7,    17,     0,     1,     1,    -5,    12,     4,    -3,     7,     2,    -1,   -11,   -19,   -21,     1,     2,   -15,    -3,     7,     3,     6,     7,     2,    -9,    -3,    -2,    -6,     8,   -10,    -1,    -1,    -3,   -11,     8,     3,    -4,     6,    -2,    -9,   -21,   -23,   -20,    -7,    -3,    -6,     4,    12,     2,     5,     8,     1,    -3,     1,    -2,   -10,    -3,    -3,    -1,    -2,    -4,   -10,    12,     8,     4,    14,     2,   -10,   -16,   -20,   -15,    -3,    -2,     2,     2,    10,    -9,    -5,    -5,     4,     1,     1,    -5,    -4,     0,    -2,     0,     1,     2,    -3,     9,     9,     6,     3,    -1,    -8,   -12,   -15,    -9,    -1,     2,    -1,    -4,   -17,   -12,    -3,    -8,     0,     4,     6,     2,     1,    -4,    -6,    -2,     1,    -3,    -5,     6,    15,    -1,     3,    -1,    -8,   -12,   -17,    -5,    17,     3,     2,     3,    -7,    -6,    -9,    -4,     5,    10,     8,     7,    -1,    -2,   -11,     2,     2,    -2,    -5,     3,     3,    -2,     1,     4,    -6,    -8,   -18,     1,     9,    -4,    -9,    -1,     1,    -7,    -7,    -4,     4,     4,     8,     6,     0,    -1,    -2,    -1,     0,     1,    -7,     2,     3,    -3,     4,     0,    -1,   -10,    -7,     8,    11,   -16,   -11,     0,     2,    -2,    -2,    -9,    -3,     1,     6,     4,    -1,    -3,    -4,    -2,     0,     1,    -4,     6,     2,    -4,    -2,    -1,    -1,    -9,     0,     0,     6,    -7,    -3,     1,    -3,    -1,    -9,   -10,     0,     5,    10,     4,    -2,     2,   -16,     1,     1,    -4,    -2,     8,     1,    -7,    -6,    -6,    -4,    -5,    -3,     6,     0,     3,    13,     1,     1,     6,   -10,    -6,    -1,     6,     5,    -2,     3,     0,    -7,     1,     1,    -1,     6,     0,     2,    -4,    -6,    -5,     1,     4,     1,    -4,     6,     0,     2,    14,     0,     5,    -2,    -9,    -1,    -1,     6,     0,     0,    -3,    -7,     1,     0,    -1,     2,    -4,     3,   -10,    -8,    -8,    -2,     0,     6,    -5,     2,    -5,     6,     3,     2,    10,     4,    -2,    -4,     4,     6,    -1,    -2,     0,    -6,    -2,    -2,    -2,     8,     1,    -1,   -10,   -12,   -10,    -1,     1,    -1,    -3,     0,     3,     7,     1,     2,    10,    10,     7,     3,     0,    -8,    -4,     3,   -11,    -1,     0,    -3,    -2,    -6,    -5,    -7,    -3,   -14,   -12,    -5,     2,    -4,    -4,     3,     3,     7,     4,    10,     9,    -7,     0,    -6,   -14,    -7,    -5,     5,    -4,     0,    -2,     2,    -2,    -6,    -2,    -7,    -1,    -7,    -6,     2,     0,    -1,     0,     8,     3,     4,     3,    -6,    -8,    -4,     0,    -4,    -9,    -7,    -6,    -5,    -3,     1,    -1,    -2,     0,    -7,     0,    -4,   -10,    -6,     2,     0,    -5,    -7,    -1,     6,    -5,     3,    -3,    -5,   -14,     1,    -1,    -7,   -10,   -12,   -12,    -4,     0,     2,     0,     2,     1,    -4,    -5,     0,    -4,    -7,    -5,    -5,    -3,    -7,     0,   -10,    -6,     4,    -7,   -14,    -7,    -6,    -5,    -1,    -7,    -8,    -9,    -1,    -3,    -2,    -1,    -2,    -2,    -2,    -2,    -3,     1,    -1,    -3,    -2,    -7,    -4,    -2,    -2,    -5,    -2,    -1,    -3,    -5,   -11,    -6,    -3,    -2,    -2,    -1,     1,     1,    -2,    -2,     1,    -2,     2,    -3,    -3,    -6,    -4,    -2,    -4,     0,    -3,    -4,    -3,     1,     0,    -1,     1,     0,    -2,    -9,    -3,     0,     3,    -2,    -1,    -1,    -1,    -2,     2,     1,     2,    -2,     0,    -1,    -1,    -2,     1,    -3,     0,    -1,     0,     1,     0,     1,    -2,    -1,     1,    -5,    -3,    -1,     1,     0,     0,     0,    -1,    -2,    -1,     2,    -2,     0,     0,    -1,    -2,    -2,    -1,    -3,    -2,    -1,    -2,     0,    -2,    -1,    -2,    -2,     1,     2,    -2,     0,     1,    -1,     2,    -2,     1),
		    57 => (   -1,    -2,     2,    -1,    -2,     2,    -2,    -2,    -1,     1,    -1,    -1,     1,    -2,    -1,    -2,     2,     0,     0,    -1,     0,    -1,    -1,     0,     2,     1,     0,     2,     0,     0,     0,    -1,     1,    -2,     2,     1,    -2,    -1,    -1,   -10,   -11,    -9,    -6,   -21,   -25,   -26,    -6,     1,    -2,     0,    -2,     0,    -2,     0,    -2,     0,    -1,    -1,    -1,    -2,     1,     1,    -5,    -5,   -15,   -15,   -23,   -20,   -12,    -8,    -6,   -13,   -10,    -6,    -7,     0,   -13,   -11,   -10,    -9,    -8,    -4,     1,     1,     0,    -1,    -1,    -6,    -5,   -17,   -26,   -26,   -24,   -16,   -24,   -35,   -35,   -25,   -23,   -21,   -15,   -10,    -9,   -16,    -8,   -13,   -38,   -25,   -12,    -6,     0,    -2,     1,     1,    -2,   -10,   -11,   -19,   -26,   -36,   -39,   -47,   -50,    -8,    -2,    -4,    -7,   -12,   -27,   -37,   -30,   -20,   -15,   -14,   -23,   -31,   -31,   -18,    -4,     2,     2,     2,     1,   -13,   -19,    -8,   -15,   -10,    -3,     6,    -6,     6,    10,     9,     0,    -3,    -6,   -18,   -25,   -32,   -33,   -21,   -21,   -46,   -34,   -30,    -3,     1,     1,    -1,    -7,    -6,    -5,     6,     5,     4,     1,     5,    14,    13,     1,     2,   -11,    -5,     5,    -7,    -2,   -13,   -17,    -9,   -14,   -16,   -20,   -21,   -13,   -10,     1,     8,    -7,     2,    -2,    18,    11,    12,     9,    11,    14,    -1,     5,     8,     7,     1,     7,     9,    12,     6,    -4,    -3,    -3,    -6,   -15,   -32,   -20,   -13,    -9,     5,    -2,     9,     0,    15,     1,     4,     2,    -6,     8,     9,   -11,   -14,    -9,     6,     9,     6,     9,     7,     7,     6,    -4,    -1,   -15,   -18,   -19,    -9,    -2,     6,     7,     6,     9,     1,    -3,    -2,    -1,    -3,     2,     7,    -2,    -5,   -12,     1,     2,    12,    10,     3,     0,    10,     3,     8,   -14,    -3,    18,    25,    -2,    11,    -2,    -6,     6,   -13,     2,    -7,     2,     3,     0,     5,    -9,   -12,    -2,     1,     9,     9,    13,     8,     7,    -3,     8,    -3,    -2,    10,    16,    22,    -1,     0,     0,    -5,     8,     6,    -9,    -5,    -2,     8,     3,    -9,    -4,    10,    -3,    -1,     8,     4,    11,     7,    -7,     2,    11,     9,    -4,   -15,    -1,    14,    -1,     6,    10,     1,    10,    14,     1,    -9,     9,    -3,   -10,    -4,    -3,    -3,    -3,    11,     8,    10,     4,     1,    -1,     3,     1,     5,     2,     8,    14,    23,     0,     4,    14,     0,    10,    12,    -4,    -5,     4,     0,    -1,    -1,    -7,     1,    -7,     3,     2,     2,    -1,     2,    -5,    -2,    12,     4,    11,    12,    -2,    -6,     0,     6,     5,     2,     0,     9,    -9,     6,     5,    -3,     0,    -3,     1,    -6,    -4,     1,    -5,     7,     0,     5,    -4,    -5,     3,    -5,    -3,   -24,   -22,    -4,     2,     0,    -2,    -1,    -5,    -8,     0,     3,     2,     5,     7,     3,    -3,     1,     6,     9,    -5,     1,     5,     5,    -2,    -1,    -7,   -15,   -21,   -25,    -3,   -16,     1,     0,    -3,   -12,     3,     6,    -7,    -8,    -5,     4,     5,     1,     5,    13,     8,    20,     4,     2,     1,    -6,    -9,    -6,    -2,    -5,    -9,   -22,   -17,   -16,    -2,    -3,    -9,   -17,     5,     3,    -1,    -9,    -8,   -17,    -5,    -6,    10,    12,     9,     8,    -2,    -6,    -8,    -7,    -4,    -4,     0,    -1,    10,   -13,    -7,   -17,     4,     1,     5,   -29,     1,    -3,   -11,    -9,    -8,    -9,    -7,    -1,     2,     3,     5,    -5,   -16,     1,    -1,    -7,    12,    11,     3,    11,     3,   -20,     2,   -12,     2,     3,    -2,   -11,    -8,    -2,    -5,   -13,     0,    -7,    -9,    -2,     5,     8,    -2,   -17,    -1,     0,    -2,    -2,     4,    14,    -5,   -11,     8,   -22,   -19,    -6,    -1,    -1,    -6,    -6,   -22,   -17,   -13,    -9,   -17,    -6,   -16,   -15,    -7,     4,     2,    -9,    -2,     1,   -18,    -2,     2,     3,    -8,   -21,    -9,   -19,   -16,     2,    -2,     0,    -9,   -15,   -21,    -2,    -5,    -5,    -6,   -15,    -4,    -6,    -5,     4,    -5,    -3,     3,     0,   -14,    -7,    -8,    11,    -8,   -18,   -27,    -7,    -5,     0,    -4,    -4,   -12,   -14,    -1,     2,     0,    -6,     6,    -1,    -6,    -2,     3,    -7,    -1,     1,    11,    -1,    -3,     4,    10,    -1,   -12,   -48,   -25,    -2,    -8,     0,     1,    -2,    -9,   -17,     3,     4,     4,     3,    11,     6,     0,     5,    14,     8,    16,     2,     8,     8,     0,     0,     8,    -2,   -12,   -42,   -22,   -12,   -19,    -1,    -2,     1,     7,    -6,    16,    16,    16,    15,    14,     1,     7,    11,    12,    25,    22,     1,    14,    10,     2,     9,     8,     5,    -3,   -29,   -16,   -16,   -12,     2,     0,    -2,    -2,     6,     7,     9,     8,     9,     8,    11,    19,    18,    14,    11,     5,    -7,    22,     9,     6,     6,     0,    12,    13,    -4,    -4,   -13,    -9,     2,     0,     1,     2,    -9,    -7,   -12,     1,     9,     9,    14,    14,    15,    14,   -12,   -22,    -2,     9,     1,     4,    14,     7,    11,    14,     5,    -6,    -2,    -2,    -1,    -1,     1,    -1,    -1,     5,     5,    -3,    -6,    -1,     7,    11,     2,    -1,   -17,    -4,     4,    -6,     8,     5,     5,     4,    12,     6,    15,     1,     0,    -2,     1),
		    58 => (    1,    -1,    -1,     0,     1,    -2,    -1,     2,    -1,     1,    -2,    -2,    -1,    -2,     0,     1,     1,    -2,     2,    -1,     2,     0,     2,    -1,     0,     0,     0,     2,     1,     1,    -1,    -2,    -2,     2,     0,     1,    -1,     1,     2,    -4,    -7,    -4,    -5,    -3,    -7,    -7,    -8,    -3,     1,     2,    -1,     2,     0,     2,    -1,     1,    -2,    -2,    -1,    -1,    -1,    -2,    -4,    -6,   -15,   -15,   -21,   -11,    -1,    -1,    -8,    -8,   -13,     3,     2,    -7,    -7,    -7,    -7,    -3,    -2,    -2,     0,    -1,     0,    -1,    -4,    -6,    -4,    -8,   -16,   -30,     3,     7,     7,    -1,    -8,   -10,    -7,     8,    -9,   -12,     2,    -8,    -6,    -7,     7,    14,     0,    -5,    -8,     2,    -1,    -7,    -7,   -18,   -16,   -18,   -10,    10,    22,    19,    15,     8,    -2,    -1,     7,     7,     6,    16,    -3,   -10,   -13,   -16,    -8,   -13,   -17,     2,     9,    -3,     1,     2,   -13,   -15,   -13,   -18,    -2,    25,     9,    11,     6,    13,    14,     6,     1,     4,     7,    14,    -1,    15,    -1,     2,     6,    -5,    -6,    -4,   -13,    -5,     1,    -2,   -20,   -17,   -18,    -9,    -6,    12,    -5,     1,    10,     2,    -1,     4,    -2,     5,    -1,    -3,     4,     4,    10,     1,    -2,     7,    -5,    -8,    -4,    -3,     1,   -13,   -16,   -20,   -16,   -12,     0,     1,    -2,    -1,    -2,    10,     0,     3,   -10,     7,     3,    -2,    -3,     3,    -6,    -3,    -5,    19,    11,   -19,   -12,     6,     4,    -9,   -14,     2,    -2,    -1,    -2,    10,     4,     2,     3,     1,    -2,     2,    -1,    -2,    -3,    -1,     7,    17,    -7,    14,    11,    18,    19,   -11,    16,    18,     1,    -5,   -19,     4,    10,    -5,     1,     9,     5,     0,    -6,     0,    -2,     0,     5,    -3,    -4,     5,     2,    -2,    11,    11,    11,     8,     4,    -5,    16,   -20,    -2,    -2,   -22,   -15,    20,     6,    -7,     7,     7,     4,    10,     4,     4,    -3,    10,   -16,   -13,     1,    -3,     0,     3,    12,     5,    11,     8,   -17,     7,    -8,     2,    -3,   -10,     0,    19,    16,     4,    11,     3,     1,     4,     0,    -5,    -5,     3,   -14,   -13,   -10,     1,     0,     5,     7,     9,    10,    13,     4,    19,    -4,    -1,     1,   -15,     4,    19,    33,     1,     1,    11,     5,     0,    -7,   -10,   -10,    -1,    -7,     1,    -1,    -8,    -5,     7,     7,    17,     2,     8,    -7,    10,   -17,     2,    -2,    -9,    -1,     7,    18,     6,     3,     8,     1,    -1,    -3,    -2,    -4,    -2,     3,     0,   -13,    -6,    -5,     9,     4,    15,     1,   -10,   -11,     8,     3,     0,    -4,    -4,   -12,   -18,     2,    11,   -16,     9,   -20,   -14,    -4,    -8,    -9,     1,     2,    -5,   -14,     0,   -12,   -17,     5,    -1,    -5,   -14,    -2,    -9,    -6,     2,     2,    -7,     6,   -29,    -7,   -10,   -11,     5,   -12,    -4,    -4,   -14,     2,     5,    -8,    -6,     2,   -11,    -5,    -8,   -13,    -4,   -16,   -21,    -5,   -23,   -13,     2,    -3,    -4,     8,   -28,   -12,   -14,   -23,   -12,    -1,   -15,   -10,    -2,     8,    -1,    -4,   -11,   -19,   -10,    -1,   -10,   -15,    -8,    -5,    -8,    -8,   -26,   -13,     1,    -3,    -6,   -14,    -8,   -14,   -16,   -15,    -2,   -10,   -10,   -16,    -4,    -5,    -8,   -15,    -7,    -6,    -7,    -3,     1,    -4,    -4,    -2,    -3,   -25,   -12,   -19,    -3,    -3,    -9,   -25,     0,   -14,     0,     4,     2,    -2,    -5,    -7,     3,    -1,    -9,   -27,    -1,     2,     0,     5,    -2,    -5,     1,     0,     1,   -23,   -10,   -12,     1,     1,   -19,   -23,    -5,   -14,    -9,     4,    15,     4,     3,    -6,   -10,    -9,   -16,   -11,    -3,    11,     1,     5,     6,    -8,     4,    12,    15,   -30,   -22,   -15,     1,     0,    -7,   -19,   -15,     3,     7,     2,    13,    -5,    14,    -1,     7,     0,   -10,    -4,    12,     8,     2,     0,    10,    10,    10,    25,     6,   -37,   -23,     1,    -6,   -10,    -9,   -11,   -12,     3,    17,     2,    10,    17,     7,     6,     4,     9,     8,    20,    -1,    13,   -14,     6,     1,     2,    18,    16,    -6,   -28,   -17,     0,    -7,    -8,    -5,    -9,     7,    17,    10,    15,    13,    13,    18,    18,     8,    14,    23,    23,     4,     3,     6,    -5,     0,     0,    16,     9,    -9,    -2,   -17,    -1,    -2,     2,    -3,    -4,    16,    -1,     6,    -4,     7,     7,     2,     3,    15,    15,    15,    17,    15,    13,    15,    21,     5,    -6,    21,    11,    -5,    -2,   -18,     0,     2,     1,    -7,   -11,    -6,    -7,    -4,    -5,     6,    11,     5,     2,    14,     4,     6,    10,    22,    -2,    -1,    -3,     2,   -11,     3,     4,   -10,   -24,   -13,    -2,     2,     0,    -8,     1,   -30,   -24,    -2,    -2,   -10,   -18,    -9,   -10,    -6,    -5,     7,     8,    -3,    -6,     5,    -2,   -17,   -15,   -16,    -8,   -10,    -6,    -4,     0,     1,     1,     0,    -7,   -13,   -24,   -22,    -5,     4,     1,   -11,    -6,     5,     4,   -19,   -41,   -19,   -11,    -9,   -30,   -26,   -12,   -14,    -5,    -1,     1,     0,    -2,     0,     0,    -1,     1,    -6,    -5,    -6,    -4,    -8,    -7,    -2,    -2,   -10,   -16,   -19,   -15,    -8,   -13,    -6,    -7,     0,     0,    -5,     0,    -1,    -2,     1,    -1),
		    59 => (    2,    -1,     2,    -1,    -2,     2,    -1,    -2,     2,     0,     2,    -2,     1,     1,    -1,    -2,    -1,    -3,    -1,    -1,     2,    -1,    -2,     2,     2,     2,     1,    -2,     1,     2,     0,    -2,    -2,     2,     1,     0,    -2,    -1,     0,    -3,    -4,    -6,     2,    -3,    -1,    -4,     0,     2,     1,     2,     1,    -2,    -2,    -2,    -2,     2,    -1,    -2,     1,     2,    -2,     1,    -2,    -2,    -4,    -3,    -1,    -4,    -2,    -2,    -8,    -2,     2,    -2,     1,    -2,    -2,     1,    -1,     0,    -1,    -2,    -1,     2,    -1,    -1,     1,    -2,    -4,    -5,    -4,     0,    -6,   -10,    -3,    -8,    -3,   -11,    -7,    -8,    -2,     2,     4,     0,   -10,    -7,    -3,    -3,     1,    -3,     1,     2,     2,    -1,     1,     0,    -1,    -3,   -10,    -3,    -3,     0,    -5,     0,   -14,   -19,   -16,   -13,   -11,   -11,    -5,   -14,   -15,     0,    -2,     0,    -2,   -11,    -9,    -2,    -2,     0,     0,    -1,    -3,     1,    -2,    -6,   -20,    -8,    -9,     1,     3,     0,     3,     0,    -5,   -15,   -19,   -11,    -2,    -3,     0,    -1,     1,   -10,    -5,     1,    -1,     1,    -3,    -2,    -7,   -11,    -9,   -15,    -3,     7,     1,    12,    11,     9,    -1,    -5,     7,    -3,   -25,   -23,   -11,     0,     1,    -2,     0,     0,    -2,    -7,    -2,     0,    -3,     2,    -5,   -12,   -18,   -14,    -1,    -9,     3,    10,     1,     5,    -6,   -15,   -12,   -13,   -27,   -34,   -12,     2,    -1,     0,    -4,     0,    -2,    -6,    -5,    -3,    -5,     6,     2,   -13,    11,    -3,     9,     1,    -1,     2,    -3,     2,    -3,   -11,   -13,    -7,     3,    -8,   -18,    -3,    -3,    -5,    -6,    -2,    -1,     0,    -2,    -9,    -8,     3,    -1,    -8,     8,     8,     3,     6,    10,    -5,    -6,     3,     2,   -10,   -15,     7,     6,    -6,   -12,   -10,   -12,    -5,    -9,   -12,    -6,    -6,    -1,    -3,    -4,     4,    -3,   -13,    11,     6,     5,     2,     1,   -21,   -18,     3,    12,    -2,     7,     0,     0,    -6,   -11,   -12,   -14,    -9,    -8,   -10,    -2,    -9,    -2,   -14,    -6,     6,    -6,   -14,     5,    11,     9,     2,    -4,    -2,     8,    26,    -1,    -2,    -2,     9,    -4,    -1,   -18,   -20,   -13,   -12,    -4,    -9,     0,    -8,     2,    -5,    -6,     8,    -5,     5,     4,    -2,    -1,    10,     5,     2,     8,    17,    -7,   -14,    -3,     7,     0,    -1,    -7,   -11,   -18,   -14,    -8,    -7,    -8,    -9,     2,    -6,    -4,    -7,    -9,     1,    22,     3,   -10,     2,     4,    -5,     0,    -3,    -5,    -3,    -1,    -2,    -8,     5,    -8,   -11,   -10,   -10,    -5,    -5,    -7,     0,    -2,    -1,    -4,    -5,    -6,    -6,    14,     2,    -5,    -4,    11,     0,    -8,    -5,     4,     4,    -3,     0,     0,     0,    -7,   -13,   -14,   -15,    -6,   -10,    -1,    -1,    -3,    -1,    -4,    -5,     7,   -10,    -9,     2,    -3,    -7,     5,     2,    -5,   -15,    -6,     4,     4,     0,    -4,    -4,   -22,   -20,   -14,   -13,    -4,    -3,     0,    -6,    -2,     0,    -7,    -1,    -1,    -6,   -22,    -2,     4,    -8,     3,    24,     8,     3,     1,   -10,    -8,    -8,    -3,    -9,   -29,   -11,    -6,    -5,    -4,    -3,     1,   -10,    -1,    -1,    -9,     1,    -1,    -8,   -17,   -20,    -2,   -15,    -5,     6,    11,     7,     2,     1,   -12,   -12,    -8,    -7,   -19,   -12,    -4,    -7,   -11,     8,    -8,    -5,    -3,     0,    -8,    -1,     1,     0,    -5,   -13,   -16,   -15,   -16,    -7,     9,    -4,    -4,    -5,    -3,     0,   -11,    -4,    -8,   -14,     0,    -5,   -13,    -2,    -6,    -5,    -2,    -1,    -6,    -2,     0,    -4,    -2,     0,    -3,    -3,   -13,   -21,   -19,   -18,   -14,     8,     4,     1,    -8,    -8,   -12,   -14,    -7,     0,    -9,     9,    -6,    -5,    -1,    -3,     0,    -4,    -1,     0,    -1,   -10,    -1,   -10,   -11,   -18,   -24,   -14,    -1,     2,    -2,    -3,    -6,    -7,    -6,    -5,    -5,    -6,     2,     6,    -8,     0,     2,    -2,     1,    -4,    -2,     7,    -3,    -3,    -1,     2,     2,    -3,    -6,    -2,     2,    -8,    -2,     0,     0,   -13,    -5,    -9,    -5,    -2,     5,    10,   -11,    -2,    -1,    -2,    -3,     6,     0,     2,     4,     4,     5,     8,    -4,     3,     7,     3,     3,     5,    -2,     5,    -3,   -12,    -8,   -14,    -3,     0,     3,    -3,    -1,    -1,     2,     2,    -5,     3,    -2,    -2,     5,    -1,     4,    -3,     2,    -3,     0,    -1,    -1,     7,     1,     5,     7,    -5,    -5,    -7,    -2,     5,     3,     2,    -5,     0,     0,     0,    -1,    -1,    -3,     2,     0,    -7,     1,    -5,     6,    -6,   -17,   -13,    -4,     3,     6,     4,     5,     6,     5,     1,    -2,     4,     3,     4,    -1,     0,    -1,    -1,     4,    -1,    -2,     1,     1,    -4,    -3,     4,    -8,   -10,    -7,     3,   -13,   -10,     2,     9,     3,   -10,   -13,   -11,   -10,    -5,    -3,     4,     1,     2,     1,    -1,     2,     4,     0,     0,     0,     1,     3,     7,    -5,   -11,    10,     1,    10,     6,     3,    23,     9,   -10,     2,     1,    -2,     3,     3,     2,     0,    -2,    -2,    -1,     0,    -2,    -2,    -2,     4,     6,     3,    -7,    -3,     2,    -1,    -8,    -9,    18,    17,    -2,    -4,     8,     3,    -7,    -5,    -1,    -1,    -1,     2,     1),
		    60 => (    1,     0,     1,     2,     2,     0,     2,     2,     0,     0,     1,     2,     0,     0,    -2,     1,    -1,    -2,    -2,    -2,     2,     2,     0,    -2,     0,     0,    -1,     2,     0,    -1,     2,     1,     0,     1,    -1,    -5,    -5,    -6,   -11,    -5,     2,     3,   -14,    14,    17,    17,     1,    -2,    -3,    -3,     1,     0,     2,     1,     0,     0,     0,    -2,     2,    15,    18,    -5,    -8,     3,    -3,   -10,   -16,   -14,   -17,   -33,   -17,    -8,    -1,   -12,    -8,    -9,    -9,    -8,   -23,    -9,   -11,    -2,     1,     2,     2,    -1,     2,    16,     5,   -15,   -18,   -15,   -15,   -12,    -8,   -19,   -26,   -12,   -14,   -15,     6,     6,     0,   -12,   -12,   -18,   -25,   -13,    -9,   -10,   -19,     2,     0,     0,    -2,    -4,    -6,   -31,   -11,   -13,     1,    13,    -1,     2,   -15,     0,    -6,     5,    14,     6,    -1,     0,   -11,   -11,    -4,    -7,   -21,   -35,   -14,     1,    -1,    -2,    -8,    -5,    -7,   -16,     7,    -3,     3,    19,    12,    10,     2,     2,     8,     8,     8,     8,     8,     0,    -1,    -2,    -9,    -6,   -19,   -30,    -7,    -4,     1,     1,   -11,    -1,   -20,     5,    12,    12,    11,     8,    13,     6,     2,     1,     7,    -7,     3,    -3,   -10,     3,    -2,   -12,    -1,   -23,   -13,   -35,   -10,    -3,     0,    -5,   -10,   -11,   -12,    -1,    11,    11,    -5,     6,    -3,     2,     3,     4,   -11,   -13,    -5,    -3,    -4,   -11,    -3,   -10,    -2,    -1,   -12,    -7,   -18,     3,    23,   -14,    -1,   -15,   -14,     1,     1,   -11,     2,     4,    -6,   -11,     1,    -3,   -19,    -2,    -4,     9,    -2,    -5,    -6,     3,     0,     9,   -14,   -33,   -17,    -4,    -3,    -4,     8,     0,    -3,     4,   -11,    -6,    -2,     5,    -4,     4,     9,     3,     4,     9,     6,     8,     4,     5,     4,    -4,     0,     8,    -3,   -20,    -5,    -4,    -4,    -3,    11,     4,     2,    -7,    -3,    -7,     2,     7,    -2,    -3,    -1,     7,    23,    17,    15,    19,    -3,     7,     4,    -6,     4,     9,    -1,   -12,   -15,     0,    -2,    24,   -15,    -2,    -4,   -14,    -5,    -8,   -10,    -4,    -7,    -1,     6,    27,    10,    12,    30,    23,    20,    12,    10,     5,     5,     6,    15,   -14,   -15,    -1,    -2,     1,   -15,    -5,     8,   -15,   -13,   -15,   -12,    -3,    -6,     1,    14,    21,    14,    17,    12,    11,    12,     8,    -6,     1,    -1,     4,     7,    -7,   -12,    -8,     0,     2,     0,    -6,    10,    -2,     1,    -9,    -3,   -10,    -8,     4,     6,     2,    -1,     3,     0,    -5,    -2,    -4,    -5,     4,     2,    12,     4,     7,   -21,    -8,    -2,     0,    -3,   -20,    -7,    -4,    -9,    -3,    -1,    -6,    -6,     1,    -6,    -4,   -19,   -22,   -22,   -10,     5,    -4,     8,    18,    18,    10,    17,    14,   -18,    -2,    -2,     2,   -12,   -18,    -4,    -9,   -11,     5,    -1,   -13,   -12,    -9,   -14,   -13,   -30,   -17,   -12,    -3,    -7,    -1,    11,     7,     2,     8,    13,    16,   -19,   -17,    -2,     0,    -7,    -9,     7,    -5,   -13,     3,    -3,    -7,     0,    -6,   -11,   -16,   -17,    -2,   -14,   -12,    -4,     7,     7,    -4,    -6,   -11,    -2,    -5,   -27,    -6,     1,    -2,   -10,     1,     3,     2,    -8,     5,    -2,     3,     6,     9,     4,    10,    -7,    -6,   -10,    -2,    -2,     6,    -2,   -16,    -4,    -6,    -3,   -18,   -17,     5,    -1,    -1,    -8,    -6,     9,     8,     6,    -4,     3,    10,    11,     5,     2,    -6,   -13,    -4,    -4,     3,     3,     3,   -12,    -9,    -6,     6,   -15,   -16,   -13,   -10,     2,     4,    -3,    -5,     0,    13,     9,    15,    11,     3,     0,     2,    12,    -5,    -8,     0,    -1,     2,     2,    12,    -6,    -9,    -3,     6,    -1,   -27,    -4,    -3,     0,     4,   -12,    -9,    15,     9,     7,    12,     6,    18,     0,     5,    17,     5,     1,     6,     0,     4,    -1,     2,   -11,   -14,    -6,    -4,    -9,   -32,     3,     1,     2,    -2,   -12,    -7,     1,    -2,    13,    18,    14,    11,     7,     2,    10,     1,    -3,     7,     4,     0,     4,     3,    -5,   -10,    -2,     2,   -16,   -15,    31,     0,    -2,    -1,    -6,    -7,   -21,   -12,    -3,    17,    13,     2,    18,     8,    -2,    -6,     4,    11,     7,     5,    -5,    -4,   -12,   -12,    -5,    -1,   -11,    -7,    19,     4,     1,     2,    -6,   -14,    -5,   -13,   -11,    -2,    12,    10,     7,    -9,     9,    -3,     2,     5,     5,    13,    -3,   -13,   -21,   -14,   -18,    -6,   -12,   -17,   -16,    -2,     2,    -2,    -4,    -7,     4,     8,   -14,    -8,    -8,    -4,    -7,   -23,   -15,   -14,   -13,     7,    -3,    -1,    -8,   -19,   -11,   -20,   -17,   -13,   -11,    -5,    -1,     0,     1,     1,    -2,    -5,   -20,   -12,   -22,   -32,   -18,   -19,   -21,   -12,   -19,   -11,   -13,   -16,   -36,   -31,   -31,   -35,   -25,   -28,   -20,    -9,    -2,    -1,     2,     2,    -1,     0,    -1,     0,    -6,   -20,   -27,   -13,   -10,   -19,   -13,   -15,   -10,   -12,   -15,   -24,   -20,   -18,   -18,   -22,   -19,   -23,   -14,    -9,    -5,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -3,    -6,   -11,     1,    -1,     0,   -15,    -5,    -2,     0,     2,    -8,    -8,    -6,   -11,    -5,    -8,     1,     1,    -2,     2),
		    61 => (   -1,    -2,     1,     0,    -2,     2,    -2,     1,     0,    -1,    -2,     0,     1,     1,    -2,     0,    -2,    -2,    -1,     2,    -2,     0,    -1,    -2,     0,     2,    -1,    -1,     2,     0,     0,     0,     0,     1,     0,     0,     0,     1,    -1,    -1,    -4,    -4,     3,     1,    -4,    -3,     0,     2,     2,    -2,     0,     1,     2,     1,     1,     2,     0,     2,     1,     1,    -1,    -2,    -1,     2,    -1,    -2,    -1,     0,    -9,   -10,    -9,   -20,   -20,    -8,    -6,    -1,     5,    -6,    -5,    -2,    -5,    -5,     1,    -1,     1,     1,    20,    13,     2,    -4,     1,     8,     3,     2,    -3,    -2,   -16,   -39,   -30,   -23,   -16,   -14,    -9,     0,    -1,    -2,    23,     4,    -1,    -6,    -1,     2,     2,    -2,    17,    14,     6,    -5,    -9,    -6,   -15,    -7,   -13,   -15,   -25,   -27,    12,     6,     9,     7,     6,     5,     1,     6,     6,    -7,   -13,   -15,   -13,   -11,     2,    -2,    13,    20,    12,     3,    -4,    -7,   -30,   -18,   -28,   -26,   -26,   -15,     1,     6,    -4,    -7,   -17,    -9,    -4,     5,    11,    -1,   -10,   -17,   -15,   -14,    -1,    -1,   -10,     9,    17,    -9,    12,    18,   -11,   -27,   -31,   -30,   -15,    -6,    -1,    -6,    -4,     2,    -7,    -4,     6,     0,     1,    -3,   -13,   -13,    -8,    -7,    -2,   -14,   -18,    -3,   -11,    13,    14,    17,   -21,   -20,   -45,   -26,   -14,    -6,    -1,     1,     7,     6,     0,     9,    11,     2,    -9,    -6,   -15,   -11,    -9,    -6,     0,   -14,   -15,     5,   -11,     9,    12,     4,   -13,   -15,   -19,   -22,   -25,   -12,    -1,     7,     6,     6,     3,     6,     5,     2,    -6,   -11,   -21,    -8,   -18,    -3,     2,    -1,   -13,     3,    -6,    -9,    11,    16,     9,     4,    -4,   -25,    -7,   -19,    -1,    12,    19,     5,     7,     1,    -2,    -7,    -7,    -6,   -13,    -4,    -1,    -5,    -2,     6,   -15,    -5,    -7,   -13,    -1,    12,    -4,    -3,     8,    -2,    -8,   -16,    -1,     4,     7,     5,    -4,    -7,   -18,   -24,     1,    -2,   -11,     0,     0,    15,     1,     1,    -3,     7,    -1,    12,     8,   -17,   -23,    -8,     5,    -6,   -23,     1,     3,     6,     5,     0,    -8,   -21,    -8,    -4,     0,    -5,    -3,     0,     1,    12,     0,     1,    -6,    12,    -3,    15,    14,    -5,    -9,     2,    -2,    -9,    -7,     5,    10,     2,     5,     7,   -12,   -17,    -5,    12,    -3,    -7,   -10,     8,    -1,    11,    -2,     0,    -4,     8,     4,     6,    12,     3,     8,     9,    -5,   -11,    -9,     0,    10,    -1,     2,    11,   -20,   -34,   -18,    10,    -8,    -8,   -12,     0,     2,     2,    -1,     0,     8,     5,    17,    -8,    -9,   -25,     7,    -1,     2,    -6,    -7,     4,     4,    -6,     6,    -4,     1,   -15,   -11,    17,    10,    -2,    -6,    14,    16,     0,     1,     0,     1,    17,     8,   -19,    -1,    -3,     8,     1,    -4,     4,    -1,     4,    -7,    -7,    11,     8,   -22,   -24,    -8,     2,    -1,    -9,   -12,     7,     7,    -4,     0,     2,     8,    -4,    -1,     2,     0,   -14,     1,     0,   -17,     3,    -6,     6,    -2,    -2,    11,     2,   -13,   -25,   -14,     6,     0,     7,     8,     4,     0,    -3,    -2,     1,     1,   -15,     4,    -2,     3,    -4,    -6,    -8,   -12,     8,     2,     6,    -2,   -10,    -2,   -20,   -17,   -13,    -9,     3,    -6,     1,     4,     7,    -2,    -2,    -3,    -1,    -2,    -3,    -6,   -19,   -14,   -15,    -3,     0,    -3,     4,     2,     5,    -3,    -8,   -17,   -17,   -11,   -16,   -14,     2,     0,     7,     3,     8,     1,    10,    -2,    -1,     8,     4,     0,   -16,    -5,   -10,    -2,     7,     1,     5,    -3,     6,    -1,     1,   -12,    -9,    -5,   -15,   -11,    -1,    -9,     9,    12,    14,     3,     9,     0,     0,     8,    -1,     8,    -4,    -2,    -8,     0,    -7,     2,     1,    -5,     4,     8,    -4,    -1,   -15,    -1,    -5,     9,    -5,    -2,     6,    17,    15,     2,    -1,     9,    12,    10,     7,     4,    11,    -7,    -2,     1,    -5,     4,    -9,    -1,     1,     2,     2,    -9,   -20,     0,     7,    16,     5,    -1,     9,    15,     8,     1,    -1,     8,    11,     8,     7,    -2,     5,     2,   -12,   -11,    -3,    -8,    -8,    -1,    -1,    10,    16,     7,     2,    17,     8,     0,    -3,     3,    11,     2,    -2,     5,     1,     2,     2,     0,    -2,    -3,    -2,    10,    13,    17,    19,    -2,    -4,    -2,     4,     5,    20,     8,    12,     9,    -1,   -15,   -15,    -4,    -4,     6,    13,    20,    -2,     1,     1,     1,    -5,   -19,   -17,   -16,    -2,    -1,    17,    -7,    -5,    -5,     1,     1,    12,    -3,    -2,    -3,     4,    -1,     7,     1,    -7,    -6,     8,     6,     0,     2,     1,     2,    -4,   -10,    -8,    -6,   -26,    -1,    12,   -32,   -27,     0,    -3,     9,    -4,   -14,   -27,   -14,    -8,   -14,   -10,    -7,    -5,    -2,     1,     0,    -2,    -2,     0,    -1,     1,    -4,    -9,   -20,   -25,   -22,   -22,    -8,   -12,   -21,   -22,   -11,    -6,     6,   -13,    -1,    -4,    -2,    -4,    -1,     0,     2,    -2,    -2,    -1,    -1,     2,     2,     0,     2,     2,     0,    -2,    -1,    -3,   -11,    -9,     0,    -2,    -8,    -3,    -5,     1,     2,    -2,     1,    -1,    -1,     1,     0,     1,     1,     2),
		    62 => (   -1,     1,     0,     1,     2,    -1,     1,     1,    -1,     0,    -2,    -1,    -1,     1,     4,     2,     2,    -1,     2,     2,     0,     1,    -1,     0,    -2,     0,    -2,     0,     2,     1,    -1,    -2,     0,     0,    -2,     1,     1,     4,     2,    -1,     0,     0,    -1,    -7,     6,     3,     1,   -10,    -3,    -2,     0,     0,     0,     2,     0,     2,     1,     1,    -2,     0,    -3,    -2,     2,    -1,     2,    -2,     5,    18,    14,    22,     9,    -3,    -6,    -7,   -13,   -31,   -23,    -5,    -5,    -2,     0,     4,     0,     0,     0,    -1,    -2,    -9,    -8,     5,    13,    -2,    -3,    10,    -5,     2,    -4,     1,     0,     3,    10,     0,   -16,   -14,   -16,    -9,     9,     1,     0,    -1,     2,     0,     2,     2,    -6,     5,     6,     8,    22,    21,    -6,     2,    12,    12,     8,    19,    13,    11,     0,     2,     2,    -9,     3,     5,     3,   -14,   -15,    -5,    -9,    -2,     1,     2,     3,     1,    -2,    -9,    -7,    13,    -2,    -7,     4,     2,     7,     6,     0,     7,     7,    -1,     1,    -2,   -11,     7,    16,     2,    -8,    -8,   -10,    -5,     1,     1,     6,     4,    -4,   -15,     4,     5,    -3,     0,    -3,    -5,     0,    -3,     7,    -1,     0,    -8,     3,   -11,     1,     7,    21,     4,    -8,   -11,    -6,    -3,    -1,     0,    -2,    11,     0,    -5,   -14,    -1,     6,    -3,     6,    -1,     2,     5,    12,     9,    -1,    -6,    -6,   -13,     4,     0,     9,   -15,   -12,   -16,    -3,    -4,    -7,     6,     5,     1,    11,    -7,   -11,    -5,     3,     0,    10,    10,    -2,    -6,    -9,     2,     2,     1,    -3,    -1,     0,    -1,     2,     0,    -8,   -10,   -12,    -3,    -1,    -6,    19,    -5,     8,    11,   -13,     2,    -1,     1,    -1,    -9,     2,   -23,   -37,    -4,     5,     4,    -1,    -2,     0,    -1,    -1,     7,   -17,    -9,     5,    -6,    -2,    -3,    11,     4,    -3,    -1,    -5,    12,     4,    -9,    -8,   -10,   -20,   -28,   -14,   -11,     2,     0,    -7,    -1,   -10,     3,   -17,     8,    -7,    -4,     7,    -3,     0,     0,    -5,     8,     9,    -3,     0,    -3,    -3,   -21,   -16,   -27,   -31,   -32,    -7,    -4,     1,   -10,   -12,   -10,    -4,    -5,    -8,    13,     1,     1,    -6,    -1,     2,    -1,    -6,    -4,    -1,    -2,    -9,   -26,   -21,   -24,   -24,   -19,   -23,    -9,    -1,    -9,     7,    -2,   -11,   -10,    -2,     1,    -8,     8,    -1,     4,    11,    -5,     0,     2,     8,     0,    -6,   -14,   -24,   -35,   -39,   -38,   -20,   -16,    -7,    11,    -6,    -7,     5,    -1,    -5,   -14,   -11,    -4,   -10,     2,    -5,    -1,    11,     2,     0,    -3,    -4,    -1,    -1,   -16,   -20,   -27,   -29,   -19,    -4,    -2,     1,     3,    -9,    -9,    -1,    -3,   -13,    -9,   -11,    -2,     0,    -4,    -4,     1,     8,     8,    -2,    -6,    -1,    -2,   -17,   -13,    -5,   -11,    -3,     8,    11,     7,    -5,     4,    -3,    -8,    -2,    -9,   -13,    -9,   -17,     2,    -1,    -5,    -2,     7,     8,    17,    -2,     0,    -1,    -7,   -14,   -10,     0,   -10,    -6,     4,     3,     5,     1,     1,     3,   -17,    -3,   -10,   -20,   -11,   -17,    -5,     0,    -1,    -5,    19,     8,     7,     1,     0,     1,    -2,   -12,    -3,   -14,    -7,    -2,     1,     2,     6,     9,     5,    -2,    -6,    -9,   -16,   -23,   -14,     2,     0,   -13,   -13,   -10,     9,    -3,     7,     2,     2,    -5,     4,    11,    -3,    -3,    -4,    12,     8,     3,     3,    14,    -3,    -3,   -20,   -15,   -11,    -3,    -5,     1,     2,    -1,    -9,    -7,    25,    -9,    16,     1,    -2,     4,    11,    10,     1,    -1,     8,    16,    -3,     7,     7,    15,     8,   -10,    -7,   -11,   -16,    -4,    -1,     1,     0,   -11,   -15,     9,     9,    14,    18,     0,    -1,    11,    14,    14,    12,   -12,     6,    -2,    -2,     4,     7,    11,     6,    -1,     8,     1,    10,   -14,     2,     3,     5,     0,    -2,     8,    10,    13,     2,    -1,     6,    14,    12,     9,     7,    -7,    -5,    -5,     3,     4,     0,     7,    -2,    -1,     4,     8,    -7,     1,    12,     3,     8,     9,     8,    23,    27,     9,    -1,     1,    -1,    13,    12,     3,     0,    -2,     1,     4,    -6,     6,     2,     4,    -1,     8,     8,     2,   -19,    -4,     7,     8,    -3,     5,    -7,    -1,     4,   -10,    -5,    -2,    -1,    -2,     3,    -7,     5,    -1,     4,    12,    -1,    -2,     6,     0,    -6,     5,    13,     3,   -12,     9,     4,     0,    10,     7,    10,     8,     6,    -8,    -1,    -1,     0,    -8,    -4,    -9,   -15,   -24,   -35,   -23,   -10,     1,     3,     4,     5,    18,     1,    -8,     3,    12,    11,   -10,     7,    27,    16,    16,     6,     7,    -2,     0,    -2,    -4,    -3,    -4,    -8,    -6,   -12,   -23,   -23,    -5,    -1,    -4,     0,    13,    15,     7,    21,    -2,   -21,     2,     4,     3,     0,     8,     8,     6,     2,    -1,     0,    -2,     0,    -1,    -2,    -6,    -5,    -6,    -3,    -2,   -10,    -1,   -13,   -13,    -9,   -22,   -15,   -11,    -5,    -2,    -1,    -7,     1,    -2,    -2,     0,     2,     2,     2,     1,     2,     2,     2,    -2,     2,     2,     1,    -2,    -2,    -1,    -2,     0,     2,    -2,    -2,     2,    -2,    -6,    -5,    -1,    -2,     0,    -1,     0,     2),
		    63 => (    2,     2,     2,     0,     0,     2,    -2,     0,    -1,    -2,    -1,    -1,    -2,    -1,     0,    -3,     2,    -1,    -2,    -1,     1,    -1,     0,    -2,     1,    -2,     2,    -1,     2,     0,    -1,    -1,     1,    -2,     1,    -2,    -1,     1,    -2,    -5,    -4,    -6,    -7,    -6,    -4,   -11,    -6,    -1,     1,    -2,     2,     1,     0,    -1,     1,    -1,     1,     0,     2,    -1,     0,     0,     0,    -5,   -18,   -17,     9,     8,    -7,   -13,   -18,     0,    -6,    -5,    -3,    -3,   -13,   -10,    -8,    -9,    -4,     0,     0,     2,     2,     2,     0,    -4,    -1,     5,     5,    14,    10,    -1,    -6,    10,     9,     7,    17,     6,    -9,    -4,    -8,    -6,     3,     0,   -22,   -32,   -16,   -12,     2,     1,    -2,    -2,    -8,     9,   -17,     2,    16,     6,     3,    -6,    -5,    -5,     2,     8,    13,     0,     0,   -16,   -11,    -4,    -6,     4,     2,   -40,   -36,   -18,   -16,     2,    -2,     1,    -2,    -1,    -6,    -4,     8,     1,    -7,   -13,    -2,    10,    12,     2,     5,    -2,     4,     3,    -2,     4,     5,    19,     9,    12,    10,   -34,    -6,     1,     2,    -1,     6,     2,     7,    -3,     4,    11,   -15,    -1,     5,    13,     5,     5,    -7,    -7,    -5,     3,     5,     0,    15,    17,     0,    -3,     9,   -24,   -17,    -5,     2,     4,     1,     7,    22,     7,    16,     5,     1,    -1,     4,    11,     7,     1,     8,     7,   -13,    -4,     1,    11,     0,     3,   -14,    -3,     4,   -22,   -28,    -8,    -5,     0,     1,     3,     8,     3,    -4,    -7,     2,     2,     1,     5,    -1,    -7,    10,     6,     4,    -8,     7,    16,     7,    12,    -8,    -5,    -5,   -29,   -28,    -4,     1,   -10,    -2,    -5,     6,     6,    -1,    -5,     1,    -4,    -7,    -1,    -1,     4,     9,     5,    11,     8,     5,     5,    -5,    -7,    -5,    -7,   -33,   -35,   -33,   -11,     0,   -13,    -8,    -8,    -2,   -10,   -11,    -1,    -5,     1,    -5,     1,     8,     7,    -7,     0,     4,    16,     4,   -14,    -2,   -23,   -12,    -3,   -22,   -16,   -25,   -11,    -2,   -11,   -13,     2,    -5,    -5,    -4,     5,    -1,    -8,     0,     4,     1,    -6,    -7,    -6,    -1,    24,    10,     0,    -3,   -12,   -12,   -11,   -30,   -38,   -22,    -2,     0,    -7,   -16,     0,    -5,     2,    -3,    -8,    -5,    -1,    -1,     5,    11,     0,    -6,    -3,     6,    13,    11,    12,     8,    -4,    -3,    -5,   -40,   -20,   -10,     0,    -2,    -5,   -12,     0,   -13,    -9,    -7,     0,    -1,   -11,    -5,    -1,    10,    -2,    -3,    -8,    15,    13,     3,    10,     6,     2,    -9,    -5,    -3,   -25,   -19,    -7,    -4,     5,    -1,    -6,   -12,    -2,     1,    -2,    -4,    -7,     2,     5,     2,    -3,    -8,    -4,     4,    14,    11,    18,     7,    12,    -2,    -2,     7,   -26,   -18,    -3,     0,     4,     0,     0,    -5,    16,    15,     0,     0,    -4,    -9,    -1,    -7,    -2,   -10,    -6,     5,     7,     6,    12,     6,     3,     5,     4,    12,   -18,   -10,    -5,     0,     3,     1,     5,    -1,     5,    17,     9,    -4,     0,    -1,     1,     3,    -6,    -9,    -9,     9,    14,     9,     4,    12,    10,    -2,    -7,     0,   -25,   -27,    -9,    -1,    -1,    -1,    12,    -3,    -3,    14,    16,    -8,    -6,    -2,     1,     6,    -3,   -14,     2,    10,    10,    -3,    -7,    -2,    -2,    -4,    -5,   -27,   -25,   -12,    -3,    -7,     2,     4,    13,     1,    -3,    12,     6,     1,     4,     8,     4,     0,   -16,    -4,     8,     8,     0,    -6,     0,     4,     2,    -6,   -10,   -24,   -25,    -6,    -6,     1,   -10,    -2,     1,    12,    12,     8,    13,     6,     5,     8,    -1,   -18,   -19,    -9,    -1,   -15,   -16,    -5,    -3,    -2,    -7,    10,     2,   -15,   -23,   -23,   -11,    -1,    -6,    -7,    -4,     4,    15,     9,    11,    -2,     4,     5,     7,   -18,   -15,    -9,   -10,   -17,   -19,   -10,    -6,    -7,   -15,    13,    -2,    -4,   -17,    -5,    -2,    -1,    -2,     6,     1,    -3,     5,    10,     2,    -2,     0,     6,    17,     3,   -13,    -2,     1,     0,    -7,    -2,     3,    -3,     0,     5,    -1,   -12,   -19,    -8,     2,    -5,    -4,     8,     0,    -3,     5,     7,    -5,     4,    -3,    16,    18,    11,   -10,    -4,    10,     2,     2,     6,    -4,     0,    -1,    11,    -5,   -24,   -15,   -13,    -2,     0,     2,     3,     3,     0,     0,    -3,     2,     2,    10,    16,    19,     4,    13,     9,    13,     7,     5,    10,     1,    -2,     4,    -3,   -10,   -11,   -14,   -20,     0,     0,     0,    -5,    13,     1,    -3,     0,    12,    17,    17,    18,     2,     3,     4,     8,    10,    16,     5,    -6,    -9,     1,     3,    -3,     0,   -22,   -17,    -9,    -2,    -1,     0,     2,    -7,    -7,    12,    10,    11,    12,    15,     8,    -2,     4,     0,     7,    10,    12,    11,     7,     9,    11,     0,   -11,   -30,   -19,    -6,    -4,     1,    -2,     2,     0,    -7,   -16,    12,     8,     9,   -13,   -13,     3,     3,    -5,   -14,   -12,    -6,     5,     3,    -2,    -4,    -4,   -11,   -11,    -7,    -2,     1,     1,     0,    -2,     0,     1,    -1,     0,    -5,    -2,     1,    -4,    -8,   -10,   -11,    -6,   -10,   -11,    -8,     0,    -3,    -7,    -9,    -7,    -5,    -3,    -1,     1,    -1,    -2,    -2),
		    64 => (   -1,    -1,    -2,     0,     1,    -2,     2,     1,    -1,     0,    -2,    -2,    -4,    -5,    -2,    -2,     1,    -2,    -2,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     2,    -1,     2,    -1,     2,     1,    -1,    -9,    -7,    -5,    -4,   -10,    -8,    -3,    -9,    -4,    -6,    -4,     1,     1,    -1,    -2,    -1,    -1,    -3,     0,    -1,    -1,     0,     1,    -1,     0,     2,    -1,    -1,   -12,    -9,   -12,   -19,   -17,   -20,   -12,    -9,    -4,    -4,    -3,    -3,    -4,    -3,    -8,    -2,    -4,    -4,    -2,     0,    -1,     2,     0,    -2,     2,     1,    -5,    -7,    -2,    -6,   -17,   -26,   -14,    -1,    -6,   -15,   -11,     0,     0,    -3,    12,     4,    -6,    -2,    -8,     0,     6,    -1,     2,     0,    -2,     0,    -3,    -5,    -7,     0,     2,    -3,    -6,   -10,     0,    -3,    -7,    -9,    -7,    -9,    -6,    -8,     0,     6,    -6,    -5,     4,    15,     6,     5,    -8,    -4,     0,     2,    -1,    -3,    -3,   -10,    -2,    -9,     5,     0,     8,   -15,   -27,   -35,   -29,    -8,    12,     8,   -15,   -15,    -9,   -11,    -2,    11,     1,     7,    -8,    -2,     2,     2,    -2,   -11,    -9,    -3,     8,     3,     5,    11,   -11,   -27,   -31,   -47,   -33,    -6,     3,    10,    -4,   -21,    -7,     2,    10,    13,    -6,   -14,     3,    -6,    -2,   -11,     0,   -10,    -9,     0,    -1,     0,    11,    16,     6,   -16,   -39,   -54,   -17,     9,     7,     8,   -19,    -2,     6,    12,    26,     7,   -17,   -16,    -4,   -15,    -6,    -9,    -4,   -12,   -10,    -5,     5,     0,     4,    16,     7,   -10,   -47,   -35,   -10,     3,    13,    -1,   -16,   -11,     3,    10,     3,     8,   -20,    -3,   -12,   -13,     1,    -4,    -1,   -14,    -9,    -3,    -9,     7,    12,    11,     8,    -6,   -17,   -14,    -5,     0,     5,    -5,    -5,     0,    -1,     2,     0,    11,    -8,    -5,    -8,    -5,    -1,     2,     0,   -14,    -2,     0,    -3,     6,     8,    17,    11,     1,   -17,   -21,    -4,     9,     3,     1,     1,    -2,    -8,    -7,    -6,    -2,     6,     4,    -5,    -7,     2,    -4,    -3,    -9,     3,     5,     4,     2,    12,    16,     7,    -8,   -15,   -14,   -10,    -4,    -2,     1,    -8,    -4,     2,    -3,     2,    -6,    -3,     6,    -6,   -14,     2,    -4,     2,   -19,    -7,    -2,     7,    -4,     2,    11,     6,    -1,    -2,     3,    -3,     4,    -1,     1,    -1,     3,     9,    -2,     1,   -15,   -12,    -3,    -7,   -13,    -2,     0,    -5,   -12,   -14,    -9,     7,     5,    -3,    12,     5,     0,     0,     6,     2,     7,    -1,     2,     8,    14,    -3,     2,     2,   -19,   -19,    -1,    -8,     2,    -2,     4,   -14,    -3,     1,    -5,    -6,     4,    -9,    -6,    -1,    -2,     1,    -3,     4,    12,     3,     9,     8,     2,     3,     8,    -7,   -21,   -16,     3,    16,     2,     2,    -1,    10,     2,    12,    -1,    10,    -1,    11,    -7,    -5,    -9,   -10,     0,    -5,     8,     3,     0,    -3,     2,   -15,    -2,     3,     9,   -12,     6,    21,     2,     1,     0,    -7,     7,    -2,   -11,    -9,     6,    -2,     3,    -2,    -5,    -3,    -3,   -10,     3,    -3,    -1,    -1,    -8,   -22,     0,     3,    -2,    14,    18,     6,    -2,     2,    -1,    -4,     1,     1,    -8,    -7,     4,     3,     1,    -5,    -6,    -8,    -6,   -12,     4,     0,    -4,     0,   -11,   -10,     8,    -2,     4,     7,    19,    15,    -5,    -1,     0,    -3,    -2,    -2,   -11,    -8,     2,    -1,     0,    -9,   -15,   -16,    -5,    -7,     5,    -8,    -6,     3,    -4,    -6,    -2,    -3,     1,    -7,    -4,     1,    -4,     2,    -3,    -7,     3,    -5,    -9,    -3,     5,    -6,    -6,    -8,   -14,   -13,     0,    -2,     8,    -2,    -7,    11,    -4,   -14,    -5,    -1,    -6,    -8,   -10,     0,    -5,     2,     0,     0,    -7,    -9,    -9,    -9,     6,    -4,    -4,   -11,    -6,   -16,    -6,    -3,     1,     3,    -2,     2,     4,    -2,     3,     5,     1,    -2,   -16,     0,     0,     2,     2,    -8,   -10,     0,     0,    -3,     6,     3,    -5,    -9,   -23,   -14,    -2,    10,     2,    -2,    -3,    -1,     3,     1,     0,    -5,     9,    -1,   -17,    -8,    -1,     1,     1,     1,    -6,    -9,     1,     3,    -2,     4,    -8,   -14,   -16,   -10,    -3,     3,     3,    -6,   -12,    -3,    11,     1,     3,     6,    14,    -7,    -7,     5,     0,    -1,     1,    -2,    -2,    -5,    -7,     1,    -1,    -5,    -2,    -6,   -18,    -3,     5,     4,    -2,    -6,   -12,     5,     8,    -6,    12,     1,    -6,   -14,     5,     2,     0,     0,    -1,    -1,     1,    -7,    -6,    -6,    -9,     2,    -2,    -6,    -7,    -5,    -2,     5,     7,     0,     0,     4,     3,     3,     5,    10,    -7,   -17,     1,    -4,     2,    -1,     2,    -1,     0,    -3,    -1,    -6,    -4,     5,    -3,    -9,    -9,    -1,     6,   -14,    -7,    -7,     5,     5,     3,    10,     6,    -5,    -6,    -7,    -4,    -3,     2,     2,    -2,    -1,    -5,    -2,    -5,    -2,    -1,     2,     1,    -7,    -4,    -4,   -28,   -31,   -29,   -15,    -2,    -7,   -17,   -22,   -20,   -25,    -1,    -7,     0,    -2,     0,     2,     1,     0,    -1,     2,     0,    -4,    -9,   -10,    -6,    -4,   -10,   -10,    -9,   -10,    -4,   -11,   -17,   -12,   -10,   -11,   -13,   -14,     0,     1,    -1,     0,     2),
		    65 => (   -2,     2,     1,    -1,    -2,     0,     0,     2,    -3,    -2,     1,    -1,    -1,     0,     1,     1,     1,    -1,    -2,    -2,     2,    -3,    -2,     1,    -2,    -2,    -2,    -1,     0,     0,    -2,    -1,     0,    -1,    -1,     2,     2,    -1,    -3,    -1,    -3,    -3,    -4,    -5,    -5,    -4,    -5,     0,    -2,    -1,     1,     2,     1,    -2,    -1,    -2,     0,     1,    -2,     2,    -3,     0,     0,    -1,    -4,    -1,    -2,   -12,   -11,   -13,   -16,    -8,    -9,     9,     1,     5,    12,    -4,    -1,    -3,    -5,    -3,    -2,     0,     1,    -2,    -1,    -1,     2,    -2,    -5,    -4,    -7,   -10,     2,    -4,    -9,    -3,    -3,     4,    -8,     9,     7,     7,    15,    17,    10,   -12,    -9,     4,    16,     1,    -1,     2,    -6,    -3,    -4,    -5,   -14,    -7,   -12,    10,     9,     0,     1,   -14,    -8,    -4,   -16,    -4,     9,    -7,    -7,     4,    -1,    -6,    -2,    12,     9,    -9,    -1,     2,    -8,    -6,    -5,    -8,   -26,   -28,    -6,    10,     2,    -1,     5,    13,    -2,   -27,   -10,    -7,   -10,    -6,    11,     6,     6,    -6,    -6,     8,    12,    -4,    -2,    -2,    11,    -5,    -9,   -20,   -25,   -27,   -14,    -3,     7,    -4,    14,    13,    -1,    -8,    -9,     0,    -2,     4,    13,     5,    11,    -1,     1,    22,    23,     7,     2,    -2,    10,   -12,    -7,    -7,   -23,   -22,   -13,     8,     1,    -1,    11,     9,    -7,     7,    11,    12,    13,    14,    16,     4,    10,    -1,    -6,     9,    23,     1,    -1,    -5,   -10,   -10,    -6,   -24,   -20,   -10,    -2,    -3,    -7,    -6,    -1,    -6,     1,     7,    10,    13,    23,    17,    13,    -2,     4,     8,    -1,    -3,    12,     7,     1,    -1,   -16,   -17,   -16,   -15,    -9,    -8,   -13,     0,    -3,    -4,    -8,    -5,   -13,   -13,    -7,    13,     6,    -2,   -10,    -8,    -1,    -4,    -6,    10,     2,    12,     2,    -3,    -1,    -3,     3,    -9,    -3,   -18,    -7,     5,    -7,     0,     1,    -7,   -16,   -37,   -39,   -31,   -24,   -33,   -29,   -11,   -13,   -30,   -13,     1,    13,    15,    -2,    -1,     0,    -3,    17,     0,   -18,   -11,    -6,     0,     1,    -5,     0,    -6,    -9,   -24,   -31,   -43,   -40,   -36,   -40,   -25,   -20,   -25,   -16,    -9,     2,    13,     1,    -1,     1,     4,     8,    -7,   -15,    -6,    -5,    -3,     5,     2,     0,    12,     2,    -2,    -7,   -17,   -11,   -17,   -20,   -27,   -27,   -20,   -16,    -7,    -2,    -6,     0,    -2,     1,     7,     4,    -6,    -3,     1,    -6,    -9,    -4,    -5,    -2,     6,     7,     6,    -6,    -7,    -8,    -9,    -3,   -21,   -35,   -21,   -17,    -6,    -1,    -7,     0,    -4,    -3,    11,     3,    -9,    -4,     5,     2,     4,     0,     3,     4,    -1,    -5,     3,    -6,    -3,    -7,    -1,    10,    -3,    -8,    -6,    -6,    -4,    -2,    -2,     4,    -4,   -12,    -7,     5,     1,     8,    -8,    -4,     8,    -1,     0,     3,    -6,    -2,    -4,     4,    -5,    -1,    -6,     5,    13,    -6,    -3,     5,     1,    -3,    -8,     1,    -3,    -7,    -7,    -3,    -2,    -9,   -13,    -1,     1,     5,     7,     2,     6,     1,    -8,    -1,     2,   -13,     2,    -2,    -6,   -13,   -16,    -1,    -7,   -13,    -8,     0,    -2,   -10,     0,     2,   -10,   -12,    -4,   -10,    -3,     9,     8,     4,     9,    -5,    -4,    -4,    -3,    -5,     1,     5,    -7,   -10,   -20,    -3,    -9,    -2,   -11,     0,    -3,    -9,     4,     4,    -1,   -16,   -23,   -16,   -20,   -10,     7,    -3,    -3,   -13,   -11,     8,     3,     3,     0,    10,    -9,    -7,    -1,     3,    -2,   -11,    -6,     2,     0,    -7,   -11,    16,     0,     0,   -11,   -12,   -27,   -25,   -28,   -10,     2,    -7,   -16,     0,     7,     3,    -3,     9,    -9,    -8,     7,     7,    -6,    -2,    -3,     1,    -3,    -5,    -6,     3,     8,     3,     2,    -4,   -15,    -2,   -11,   -19,    -3,    -3,     3,    -7,     2,     2,     8,     7,    -4,    -1,     5,    -2,    -3,    -5,     2,     0,    -2,   -12,    -1,    12,     7,     1,     2,     0,     4,     5,    -1,    -2,     6,     2,     2,    -5,    -6,     3,    11,     2,    -7,     7,     5,    -4,    -2,    -8,     1,     2,     1,   -14,    13,     5,    -8,    -4,    -6,     4,    16,    12,    10,     2,    -8,     5,    -5,    -3,     4,    -2,    -1,     3,    -1,    -1,    15,    -1,    -4,    -2,    -2,    -1,     1,     6,    16,    14,     7,    10,     1,     2,    -9,     4,     8,     3,     1,    -2,     1,    -8,    -4,    -2,     2,     2,     0,     4,    16,    -3,   -10,     2,    -2,     2,     2,    -8,     3,    -4,    -4,    -1,     1,    -4,     1,     2,    -5,    -3,    -2,     1,     1,    -8,    -5,     6,    -4,    -9,     4,    20,     5,     8,   -11,    -6,    -1,    -2,    -2,    -2,    18,   -14,   -14,    -5,    -9,   -13,     1,    -8,    -6,     2,    10,    -3,    -3,   -22,     4,     4,     2,     6,    17,    26,    12,     8,     0,     1,     0,     0,     1,     0,    -1,    -2,    -4,    -4,    -5,    -7,   -13,    -3,     9,    11,     6,   -21,   -25,   -21,   -21,   -10,     5,    -8,     7,     6,    -2,    -2,     0,    -1,    -2,     2,     0,    -1,     0,     0,    -2,     1,    -2,    -2,    -4,     0,     1,     2,     4,    -5,    -1,    -1,    -1,    -3,    -1,     1,    -3,    -6,    -3,    -1,    -1,     2,     1),
		    66 => (    0,     1,     0,    -2,     2,     2,    -1,    -1,     1,    -2,    -1,     1,     8,    10,     1,    -2,    -1,     0,    -2,    -2,    -1,     2,     1,     2,     2,    -1,     0,     0,    -1,     2,    -1,    -2,     0,     0,     5,     4,     2,     1,    11,     1,     5,    12,    -5,    -5,    -3,     2,     7,    10,    12,     9,     9,     8,     0,     2,    -1,     0,     0,    -2,     1,    -3,     3,     8,     5,    -1,     3,     9,     8,     9,     6,     9,     7,    -4,     7,     8,    10,    17,    14,     8,    24,    16,    12,    10,     0,     1,     2,     1,   -14,     8,    -2,    14,    15,    15,    20,    20,    23,    24,    30,    20,    27,    19,     5,     2,     3,     2,    -8,   -10,    -7,    -1,    10,   -19,   -17,     1,     2,    -2,   -11,     1,     8,    13,    14,    19,    10,    21,    18,    10,    18,     3,    20,    17,     5,     8,     3,    11,    13,     7,    -3,    -5,    -6,   -13,    -5,    15,    -2,    -1,    -5,   -11,    18,     8,    11,    12,     8,     9,    16,     4,    -9,     8,    17,     9,     2,    12,     1,    -5,     3,   -11,    -2,     1,    14,     7,    13,     5,     1,     0,     0,     1,    13,     5,    14,     8,    -2,     6,    -3,    -8,     5,     4,     4,     2,     1,     0,   -16,     4,    -1,    -9,    -9,    -8,    -2,     5,    12,    17,     1,    -2,    -1,    -5,    14,     9,     5,     5,     1,    -5,    -8,    -3,   -11,   -15,     6,    -5,    -2,    -5,    -5,     2,    -5,    -3,    -3,    -3,     5,     1,    11,    12,    -2,    -6,    -7,   -26,    15,     5,     3,    -6,     0,     8,    -7,    -8,    -5,    -9,     0,   -12,   -21,    -9,    -5,    -2,     5,     5,    -5,    -9,    -9,   -21,    -2,   -16,     0,    -2,    -9,   -14,    12,    -3,    -9,    -6,     2,    -5,    -7,    -9,   -13,   -16,     0,     1,    -9,   -21,    -3,    -4,    -2,    10,    -2,    -2,   -14,   -26,   -16,   -14,    -2,    -2,   -10,    -8,     4,     1,    -9,   -10,    -2,    -6,    -4,   -13,   -16,    -7,     2,    -7,   -18,   -11,   -15,   -11,     2,     1,   -12,   -10,   -18,   -19,   -16,   -16,    -1,    -2,    -2,   -16,     4,     2,    -1,    -2,    -8,    -3,    -7,   -13,     1,    -1,    -2,   -11,    -9,    -8,   -10,    -5,    -5,     1,   -11,    -2,    -8,   -16,   -17,   -12,     2,    -2,    -8,   -15,    -2,     4,    11,     3,    -4,     4,    -1,     2,    -4,     6,    -8,    -5,   -13,    -9,   -12,    -9,     7,     5,    -7,     7,    10,    -1,   -23,   -12,    -1,     1,    -5,   -13,    -6,     5,    -1,    -6,    -6,    10,    13,     9,     9,     4,     6,     2,    -3,   -15,    -4,     6,     7,     8,    -5,     8,     6,    -7,   -24,     0,     0,    -1,    -2,   -13,   -18,     6,    -8,   -13,     4,     4,    13,    13,    14,     7,     3,    -9,    -2,    -9,     4,     5,     2,     6,     6,    -7,    -3,    13,   -19,    -4,     0,    -1,    -8,    -9,   -20,    -7,    -7,    -2,    -6,    -2,     3,     7,     0,    15,    10,    -6,    -7,   -16,     1,     8,    -1,     3,   -12,     2,     0,    11,    -8,   -23,     2,     0,   -12,    -9,    -5,     4,     3,     5,    -6,     7,     7,     3,    -4,    -8,    -5,    -5,    -6,    -8,    11,    12,    -5,    -4,     4,    -1,    -4,     9,   -13,   -19,    -2,     1,   -13,   -13,    -9,    11,     1,     4,    -3,    -9,    -5,    -2,    -5,    -8,     1,     5,     5,     8,     7,     8,     7,    -3,    -3,    -6,    -3,     8,   -12,   -27,     2,    -2,   -13,   -21,    -4,    -2,    -9,     2,    -1,     3,     9,   -14,    -1,    -2,     0,   -10,     1,     8,    21,    17,     2,    -6,     1,     3,     3,    13,     1,   -12,     2,     0,   -15,   -17,     2,     6,     6,    -2,     1,     1,    16,    16,     9,     4,     2,     5,     1,    11,     0,    17,    -2,    -1,    -3,    -6,   -14,     4,    -8,    -1,     0,    -1,   -14,   -21,    -1,    -1,     1,     7,     2,     4,    13,    14,    12,    -8,     3,     4,     3,     8,     9,     8,     8,    -1,    -2,   -15,   -19,    -5,    -5,     0,    -1,    -2,   -18,   -19,   -14,   -17,    -5,    11,    14,     0,     7,     1,    21,    10,     4,     2,    17,    10,     9,     6,     3,    -5,    -4,   -16,    -8,    -1,    -2,    -3,     0,     1,   -13,   -15,   -27,   -34,   -45,     0,     1,     8,     4,     3,     1,     0,     1,    11,    13,    19,    12,     1,     4,     4,   -14,   -12,   -30,    -8,    -3,    -2,    -1,     2,     2,   -16,   -20,   -23,   -21,    -3,    -6,     1,    -9,     3,    10,    -3,     5,    11,     1,    -9,     3,     0,     1,     7,   -16,   -20,   -20,   -13,   -16,     2,    -2,     1,    -1,    -3,    -7,    -8,   -11,   -21,   -29,   -38,   -26,   -34,   -17,   -17,   -10,     3,     5,     8,    17,   -26,    -4,   -14,   -12,   -11,    -9,    -5,    -2,     0,     1,     2,    -1,    -1,    -2,    -5,    -9,    -8,    -6,    -8,    -9,     3,     8,    -5,    -4,    -7,   -12,   -12,    -7,   -19,   -18,    -3,   -10,    -9,    -8,     2,    -1,     2,     1,     2,     0,     0,    -2,    -4,     2,    -3,    -1,    -3,    -2,    -4,    -2,     1,    -1,    -4,    -1,    -3,     0,    -3,    -2,     2,    -2,    -2,     1,     2,     1,     2,     0,     1,    -2,     2,     1,     1,     0,     0,     2,    -1,    -1,    -2,     1,     1,    -1,     0,    -1,    -2,     0,     1,    -2,    -3,    -1,     1,    -2,     0,     1,     0),
		    67 => (   -2,    -2,     2,    -2,     0,     1,     1,     2,    -2,    -2,     2,     1,     2,     0,    -1,     0,     2,     1,     2,     2,    -1,    -2,     2,     2,     1,     2,    -2,    -2,     1,    -2,     0,     0,     1,    -1,     2,    -1,     2,     1,    -1,    -3,    -2,    -4,    -4,    -9,    -9,    -6,    -1,     0,     0,    -2,    -1,    -1,     1,     2,     0,     2,    -2,    -1,     2,    -1,     0,    -1,    -2,    -1,    -4,     3,    -2,    -9,   -14,    -6,    -6,    -6,     2,    -1,    -2,    -2,    -3,    -3,    -1,     2,     0,    -1,     0,    -2,    -2,     2,    -2,     0,    -4,    -8,    -9,   -14,    -6,    -3,    -6,    -9,   -17,   -17,   -13,   -12,    -8,    -6,    -3,     0,    -2,     2,    -5,    -2,    -4,    -3,     2,     0,     2,     0,     0,    -2,    -6,    -2,   -10,   -11,   -15,   -18,   -26,     1,     2,     1,    -4,   -12,   -29,   -22,   -16,   -17,   -13,     1,    -8,   -10,   -11,    -7,    -3,    -2,    -1,    -2,     0,    -7,   -10,    -4,   -20,     1,    19,     4,    -4,     0,     6,    -2,     7,     2,     3,     0,    15,    -1,   -10,    -5,    -4,    -9,   -15,    -2,    -3,    -1,    -1,     1,     7,    -5,    -5,    -4,   -13,     5,     8,    13,     6,    -2,    -3,    -4,    -4,     6,     3,     0,     9,     4,   -18,    -8,     1,   -10,   -10,    -7,    -7,    -4,     2,     6,     8,     0,     4,     0,     5,     5,     7,     5,    -2,    -5,   -10,   -10,   -11,    -1,    10,    10,     8,    12,    18,     3,    -7,    -8,   -14,    -8,    -7,    -4,   -10,     3,    19,     1,     8,     5,     3,    12,    11,     1,    -2,    -5,    -3,    -9,     1,    11,     3,     3,     5,     6,    12,     7,    -1,   -18,   -11,    -2,    -5,    -4,     4,     4,     4,    10,     9,   -14,    -3,     1,     4,    -1,     3,    -8,    -5,     3,     1,    -3,     4,    10,    -3,    -3,     5,    -9,    -5,   -11,    -7,    -2,   -10,     4,     3,     1,    -3,     2,    13,    -3,    -3,     2,    -5,     5,     3,    -9,   -17,     3,    -1,     2,     2,    -2,     0,     3,    -3,   -12,    -3,    -9,    -9,    -1,    -7,     0,     3,     3,    -2,   -10,     0,     2,    -5,     8,     3,    -5,     2,     0,   -17,   -11,     0,    15,    -1,    -1,     0,    -1,   -10,    -7,    -9,   -20,   -11,   -12,    -9,     3,     2,     2,    -8,    -2,    -8,    -2,    -8,     7,    -2,   -11,    -6,   -18,   -19,   -13,    -8,    10,    -4,   -13,    -4,   -17,   -10,   -10,   -18,   -18,   -20,    -5,    -6,     1,    -1,     6,     7,    -3,    -2,    -2,    -7,     0,     1,    -7,   -10,   -17,   -35,   -22,   -12,    -3,    -6,    -1,    -5,   -16,   -14,   -14,   -17,   -22,   -19,    -3,   -12,    -6,     0,     8,     3,     8,    -1,     6,   -14,    -7,   -13,   -20,   -36,   -28,   -18,   -14,   -10,     0,   -10,     3,     8,     2,    -6,     4,   -12,   -14,    -5,    -3,    -9,    -4,     2,    -1,     0,     6,     5,    -3,    -9,   -25,   -15,   -14,   -20,     2,    -4,    -3,   -12,    -1,    -1,     9,    11,     3,     6,     6,    -3,     1,     2,     5,    -3,    -5,     1,     1,     0,    -7,    -4,     0,   -16,    -8,    14,    -5,    -4,    13,     4,    -1,    -2,    11,     4,     2,    10,    -6,    -2,   -10,    -6,    -3,    -2,   -15,    -7,    -2,     2,     0,    -7,    -6,    -9,   -18,    -9,    -6,    -4,     1,   -11,     1,    -3,     1,    -3,     4,     3,     9,     6,     1,   -17,   -19,   -15,   -13,    -5,   -24,   -13,   -17,     3,     1,     3,    -9,    -8,    -2,    -7,     1,    -6,     3,    -1,     1,   -10,     7,     3,    13,    -1,    14,    -7,     5,     8,     1,   -12,   -16,    -9,   -18,     2,   -12,    -1,     1,     1,    -1,    -2,   -17,    -6,    -6,     6,    -5,    -4,   -12,    -5,    -5,    12,    17,    -8,    -7,    -6,     5,     9,     9,    -6,    -2,     3,    -8,   -10,    -9,     0,     7,    -3,    -1,    -3,   -13,   -10,     0,     4,     5,    -3,   -25,    -7,    -3,     5,     4,    -7,   -13,    -5,    -2,     8,    -1,    -6,   -21,   -11,    -6,   -10,     2,    -3,     2,    -3,    -5,    -4,   -14,   -19,   -18,     4,    -5,    -8,   -14,    -3,     1,     7,     3,    11,   -14,    -6,    -9,    -5,     2,    -7,   -25,   -13,   -13,    -1,    -1,    -4,     1,    -2,    -1,    -3,   -12,   -16,   -15,    -9,   -12,    -6,   -13,    -8,     9,     2,     8,     2,     4,   -10,    -5,    -7,   -21,   -31,   -22,   -13,    -8,   -13,     1,     0,     2,    -3,    -8,   -17,   -18,   -16,   -24,   -20,   -28,   -19,   -17,    -9,    -4,    -5,     0,    -3,   -15,   -22,   -15,   -14,   -15,   -14,   -11,     4,    -7,   -11,    -2,    -2,    -2,     1,     0,    -7,   -18,   -21,   -21,   -30,   -29,   -21,   -14,    -4,     0,     3,    11,    -2,    -4,   -20,   -12,    -2,    -5,    -2,   -10,    -6,    -6,    -2,    -1,    -1,     0,   -11,     0,     2,    -8,   -12,   -16,   -17,   -26,   -16,     4,    -7,    -6,    -2,    14,     1,     4,    -1,     7,     9,     6,    -4,    -8,     0,    -1,    -2,    -1,     0,    -1,     0,    -1,    -6,    -6,    -2,     8,     4,     5,    -6,    -5,     7,    10,     5,     2,     0,     3,    28,    23,    14,     4,    -3,    -4,    -1,     0,     0,     0,    -2,    -1,     0,     1,     5,     1,    -1,    -4,     0,    10,    14,     8,     6,     6,     3,    11,    10,    17,    25,    16,     7,    -1,    -5,     2,     0,    -2,    -1,    -2),
		    68 => (    2,     2,     2,     0,    -1,    -2,     1,    -2,     1,    -1,    -2,     0,    -1,     1,     0,     2,     1,     1,    -1,     0,     1,     1,    -1,     0,     0,    -2,     3,     1,     2,    -1,    -1,    -2,     2,     2,     2,    -2,     1,     0,     2,    -1,     1,     0,    -1,    -2,   -10,    -9,     0,     0,    -1,    -2,    -2,     1,     1,    -1,     2,    -1,    -1,    -2,    -2,    -2,    -2,     0,     1,    -2,     3,    -3,    -6,    -2,     0,    -2,     1,    -1,    -5,    -1,     0,     0,    -2,    -6,    -2,    -5,    -1,    -2,     2,     2,    -2,    -1,     0,    -1,    -2,    -4,    -3,    -5,    -4,    -4,     0,     0,    -2,     1,    -8,    -6,    -2,    -1,     3,    -2,    -5,     1,     2,     2,    -2,     1,    -4,     2,     2,    -1,     1,    -4,    -3,    -3,    -7,    -7,     2,     0,    -2,     7,     7,    -5,     0,   -13,   -11,    -2,     4,     1,     3,    -4,    -5,     0,    -3,     1,     0,     0,    -2,    -2,     0,    -4,   -11,   -14,    -1,    -2,     0,     1,    -6,    -3,    -6,    -6,     2,    -3,    -8,    -3,    -4,    -5,    -2,    -4,    -6,    -3,    -2,     5,     0,    -4,    -2,     0,    -5,   -10,    -2,     2,    -2,     5,    -1,    -5,    -8,   -12,    -5,   -11,    -6,     0,    -1,     1,    -3,    -4,    -3,    -7,    -3,    -2,    -2,    -4,    -2,     0,     1,    -1,    -4,     0,     3,    12,     2,     3,     1,    -2,    -3,    -7,     2,     1,     3,     4,     4,     2,     1,     3,    -7,    -2,     2,     0,     3,     0,     1,    -2,    -1,    -5,    -2,     9,    15,    16,     6,    -2,    -9,    -7,    -2,     3,     2,     2,    -1,    -6,    -8,    -5,    -4,    -4,     1,     2,     3,    -3,    -2,     1,    -4,    -1,     1,    -6,    -8,     8,    12,    14,     6,    -5,   -13,    -8,     5,    -8,    -8,    -5,    -6,   -12,   -11,    -3,    -5,     5,     6,     7,     2,    -1,     1,     7,    -4,    -3,    -2,    -4,    -8,     5,     4,    11,     9,     6,    -6,     2,     5,    -1,     0,    -4,    -5,    -7,    -5,     0,    -4,     0,     3,    -1,    -5,    -5,    -1,    -7,    -3,    -4,     0,    -1,   -11,    -6,    -5,    -1,     9,    12,     8,    12,     8,     3,    -3,    -5,    -6,    -3,    -4,    -5,    -9,    -1,    -3,    -3,     2,    -3,    -5,    -4,     0,    -9,     1,     1,    -7,   -14,   -11,    -3,     1,    -5,     5,     2,     8,     1,     0,   -10,   -10,     0,     0,    -2,    -2,    -7,    -7,     5,     2,    -3,    -4,    -7,    -7,   -11,     1,    -3,   -10,   -16,    -6,    -9,   -10,   -10,   -10,    -8,    -5,     1,     1,    -6,     3,     3,     1,    -7,    -6,   -11,    -9,    -2,    -1,    -2,    -6,   -11,    -7,     3,    -4,    -3,     2,   -15,    -7,    -6,    -8,   -12,   -12,   -17,    -8,   -12,    -7,     0,    -3,    -9,   -10,    -1,     0,    -4,   -10,    -4,    -2,    -2,    -8,    -3,   -17,    -2,     1,     2,    -3,     3,     0,    -3,    -6,   -11,    -7,   -10,    -7,    -4,    -6,    -1,    -1,    -3,    -1,    -3,    -1,    -6,    -1,    -7,    -5,    -6,    -7,     3,    -6,    -7,     1,    -4,    -1,     4,     0,    -3,    -8,    -5,    -2,    -9,     0,     2,     0,    -5,   -10,   -11,     4,     5,    -5,    -4,    -1,     0,     0,    -5,    -5,     2,    -8,    -6,     2,     0,     0,     6,    -2,    -6,    -5,    -4,    -6,    -6,     7,     7,    -1,    -7,    -8,   -12,    -6,     3,     0,    -6,    -4,     2,     5,    -7,    -3,    -4,    -2,    -3,    -1,    -2,    -1,     1,    -5,    -4,    -5,    -4,    -7,    -6,     3,     0,     3,     1,   -10,    -8,    -8,     6,     2,    -3,    -9,    -4,     8,    -2,    -4,     1,    -1,    -7,     1,     1,    -3,    -1,    -6,    -2,    -2,    -4,   -14,    -1,     6,     6,    -1,     1,    -7,    -9,    -9,    -2,     7,     2,    -3,     1,     4,     5,     0,     1,    -5,    -6,    -2,    -1,    -5,    -4,    -5,    -3,    -2,    -5,    -9,    -1,     3,     8,     3,    -9,   -11,    -7,   -10,    -2,     4,     1,     0,    -1,     8,     2,    -2,    -1,    -7,     0,    -3,    -4,    -2,    -7,    -2,    -2,    -9,    -7,    -5,    -4,    -3,     3,     4,    -2,    -6,    -5,   -10,     1,     3,     2,     1,     2,     8,     0,    -3,    -3,    -3,    -1,    -8,    -3,    -3,    -5,    -3,    -6,    -5,    -3,    -5,    -7,    -2,    -2,    -3,    -2,    -5,    -4,    -6,     3,    -2,    -1,     0,     6,     2,    -2,    -9,    -3,    -1,     1,     2,     2,     0,    -4,    -4,    -8,    -7,    -5,    -3,    -6,    -1,    -8,    -4,     5,    -4,     0,     3,     1,    -2,     1,     4,     7,     3,    -4,     0,     0,   -11,     0,    -2,     2,    -3,     1,    -2,    -5,    -4,     2,    -4,    -1,     0,    -8,    -7,    -8,     2,     6,     6,    -6,   -10,    -6,     0,    -6,    -8,    -2,    -3,    -4,    -1,     2,     1,    -2,    -4,    -4,    -4,    -4,    -6,    -7,    -4,     0,     6,    -4,    -6,    -4,     0,     2,     0,    -2,    -5,    -4,    -8,    -6,     0,    -1,    -3,    -2,    -5,    -2,     0,    -1,    -1,    -1,     0,    -4,    -3,    -7,    -3,    -8,    -7,    -6,    -7,    -5,    -9,    -8,    -3,     0,     0,   -10,   -12,    -1,    -8,     0,     1,     1,     0,     0,    -1,     2,     2,     1,    -1,     1,    -1,    -2,    -1,    -4,    -3,    -1,     0,    -3,    -3,    -2,    -4,    -3,    -7,    -1,    -1,    -1,    -2,    -2,     0,     2,    -2,     1),
		    69 => (   -2,    -2,     2,     2,     2,     2,     0,     2,    -2,     2,     2,     2,    -1,     1,     0,     1,    -2,    -2,     2,    -2,     0,    -1,     1,    -1,     0,    -2,     0,     1,     0,     2,     2,    -2,     0,     0,    -2,    -4,    -5,    -5,    -4,    -6,    -8,   -11,    -6,   -13,   -12,   -12,    -6,     0,     2,    -2,    -6,     0,     2,    -2,    -2,    -2,    -2,    -1,    -2,    -9,   -10,    -2,    -2,   -11,   -14,    -6,    -7,   -10,     1,     0,   -28,   -16,   -15,    -9,   -16,   -12,   -21,   -24,   -17,   -14,    -9,    -4,     2,     1,     0,    -1,    -1,   -12,   -15,   -13,    -8,   -15,   -32,   -40,   -54,   -48,   -32,   -41,   -38,   -41,   -54,   -47,   -15,   -20,   -33,   -29,   -24,   -14,   -12,    -8,     2,     1,     2,    -2,    -7,   -11,   -17,   -22,   -31,   -22,   -24,   -27,   -17,    -5,     2,    -3,    -9,    -9,    -7,   -16,   -29,   -56,   -36,   -30,   -30,   -15,   -13,   -22,   -15,     1,    -1,     0,    -7,   -10,    -8,   -13,   -14,    -9,   -20,     3,     4,     1,     7,    16,     5,     6,    13,    13,    -2,    -8,   -16,    -7,   -33,   -14,   -20,   -21,   -15,    -4,    -1,     2,    -7,   -21,   -16,   -20,   -10,    -6,    -1,    10,    10,    -5,    -4,    15,     7,    15,    24,    15,     3,     5,    -4,    -2,    -4,     4,     1,    -7,   -16,   -19,     0,    -7,   -14,   -18,   -12,   -21,    -3,    -2,    -4,     4,     4,    -3,     9,    18,    17,    14,    29,    18,     0,     5,     9,    -1,     5,     5,     0,     2,   -18,   -14,   -13,   -16,   -13,   -14,   -16,    -2,     6,    -3,     0,     5,     2,     1,    12,    10,    16,    24,    19,    14,    12,    15,     1,     6,     4,     9,    10,     1,   -17,    -9,    -2,   -11,   -17,   -17,    11,     4,    10,     5,     6,    11,     2,    -3,     5,    14,    13,     8,     6,     5,     4,     3,    12,     0,    -1,    -4,    -5,   -18,   -22,   -14,    -1,    -8,   -24,   -11,    11,    11,     1,     2,    -1,    -2,     1,    -1,     8,     5,     3,   -10,     0,    -6,     0,    -1,     3,   -11,    -6,    -5,   -14,     9,   -23,    -9,    -1,   -37,     0,    -8,     3,    12,     5,    -4,   -11,    -3,    -3,    -8,     0,   -14,   -12,   -13,     0,     3,    -9,    -5,     8,    -5,   -16,   -10,   -13,    -1,   -19,    -8,     0,    -4,    -3,    -7,     9,     5,     4,    -5,   -12,   -12,    -4,     0,   -11,   -13,    -6,   -10,    -6,     3,    -8,   -12,     3,    -9,    -7,    -1,   -16,   -27,   -16,   -11,    -2,    -8,   -12,    -8,     4,    -4,     3,     2,     1,    -7,    -2,    -8,     1,    -4,    -6,   -12,     3,     0,    -4,    -6,    -8,     1,   -10,    -9,    -7,   -19,   -12,    -3,    -4,    -7,    -7,    -2,     6,    -3,    -1,     3,     0,    -1,     1,    -4,     6,   -12,    -8,     5,     1,     0,     5,     4,    -1,    -8,   -11,   -22,   -10,   -23,   -14,     0,     0,    -1,   -16,    -7,     3,     2,     6,     1,     8,     5,    -8,   -12,   -10,    -3,     6,     5,     9,     5,     8,    13,    15,     6,     3,   -16,    -9,   -22,    -5,   -15,     1,    -4,   -11,    -7,     0,     9,     9,    -2,     4,     1,    -3,   -13,   -14,    -4,    11,     7,     1,    10,    -3,     7,    12,     3,    -1,   -11,    -4,   -28,   -15,   -16,     0,    -1,   -16,     1,   -10,     3,    -9,    -4,     0,     4,    -5,    -9,    -2,    -6,     8,     2,     2,     4,    -6,     1,     3,    -5,   -23,   -26,    -8,   -34,   -20,   -11,     6,     1,   -19,    14,    -9,    -8,    -2,     0,   -14,    -7,    -8,   -12,   -18,    -2,    -8,    -5,     6,     4,   -15,     3,     1,   -11,    -8,    -9,   -11,   -27,   -17,    -8,     2,    -4,   -16,     7,    -2,    -9,   -12,    -5,   -15,    -6,     0,    -4,    -3,    -9,     0,    -9,     5,    -5,    -3,     2,    -2,   -10,     0,     9,    -5,   -18,   -13,    -5,     1,    -5,   -32,     2,   -12,     3,    -1,   -20,    -6,   -10,    -6,    -6,   -13,    -9,    -6,    -9,     2,     2,    -6,     2,    -8,   -13,     0,    17,    16,     7,    -9,     0,     2,    -1,   -27,     4,    -4,     5,     5,    -5,    -7,   -14,     3,    -3,   -10,    -7,    -1,    -5,    10,     9,    -2,    -9,   -14,    -2,     4,    13,    11,    -2,   -26,     1,     1,     0,   -20,     7,    -7,    -1,    -6,    -8,    -1,    -7,     0,   -11,     4,    -6,    10,     2,    12,    11,     1,    -9,    -5,     2,    16,    16,    12,   -18,   -19,    -1,     0,     1,    -3,     4,    -7,     1,     2,    15,     6,     0,    -6,    -2,     1,     6,    13,    10,     8,     6,     5,     0,    -4,    -2,     6,    12,    19,    -9,   -13,     1,    -2,     0,    -9,   -13,    -5,     6,    17,    22,    14,    10,     4,     8,     3,     6,   -11,    -7,    -9,     5,    22,    10,    11,     2,    -9,     3,     4,    -9,    -1,    -1,    -1,     0,    10,   -11,    -2,     9,    15,    20,    14,    13,     0,     5,    -3,    -9,     7,    -4,    -2,    14,    11,     6,    10,    -5,    -2,    -7,     0,     1,    -4,     1,    -1,    -2,     0,     9,     1,     5,    10,    18,    -4,     5,    -1,    -7,     6,    -5,    13,    12,     5,     1,     6,    -2,    18,     4,    -6,    11,     5,     0,     2,     0,     1,     1,    -1,     2,     0,    -9,     4,     2,     3,     0,     5,     7,     9,     5,     7,     2,     7,   -11,     0,     4,    -6,   -14,   -11,    -9,     1,    -1,     2,    -2),
		    70 => (    0,    -2,    -1,     1,     2,    -1,    -2,     1,    -1,     2,     0,    -1,     0,     0,    -2,    -2,     1,    -2,     1,     1,    -2,     2,     0,    -1,     2,     0,    -1,     0,     2,     2,     2,     0,     0,     0,     0,    -1,     2,    -2,    -1,     0,     2,     5,    -3,     1,    -2,     1,     1,     0,     0,    -1,     2,     2,     0,     0,     1,     1,    -1,     0,     1,    -1,    -1,    -2,    -3,     1,    -4,    -4,     0,    -4,    -6,   -10,    -4,     2,    -5,    -7,    -3,    -2,     0,    -3,    -1,    -3,    -1,     1,    -3,    -1,    -2,     2,    -2,    -2,    -1,     3,    -5,    -5,    -5,   -19,   -11,    -7,     1,     7,     4,   -10,    -2,    -2,     0,     1,    -4,   -11,   -10,    -5,     2,     1,    -1,    -2,     1,     2,     2,     1,    -4,   -17,    -5,    -1,    -6,    -2,    -4,    10,    14,    16,     8,     4,   -13,   -16,    -4,     2,   -13,   -14,    -7,    -4,    -4,    -8,    -5,     0,    -1,    -1,    -5,    -2,    -3,   -11,    -4,     1,     1,     0,     2,     5,    17,     5,     5,     8,    -3,   -15,   -11,     7,    -8,   -15,     1,     3,    -1,   -12,   -10,    -6,     2,    -3,    -2,    -3,     3,     4,     6,     6,     7,     2,     0,    14,     2,    -2,     2,     0,    10,     6,    -8,     0,    -5,    -3,    -2,    -3,    -3,   -18,    -9,    -4,     0,    -2,    -4,    -9,     2,     6,     9,     7,     3,     6,     1,     7,    -1,     2,    12,     7,    13,     4,     4,     5,     7,     5,    -9,    -4,    -4,    -4,   -10,    -8,     2,    -2,     9,    -8,     7,     1,     5,    -6,    -1,    10,     7,    -3,    -6,    10,     7,    -2,    -7,    -7,     9,     1,     3,     9,    -2,     1,    -8,    -6,   -15,    -6,     2,     0,    13,    -2,    -3,    -6,   -10,    -9,     7,     8,    10,    -2,    -3,     9,    -1,     1,    -5,    -1,    -4,    11,    -2,    -5,    -4,    -6,   -10,   -10,   -12,     2,    -1,     2,    12,     3,    -7,    -2,    -8,   -10,     6,     6,    -1,     0,     0,   -11,    -3,     7,     1,    -6,   -10,    -8,   -11,    -6,    -6,     6,    -2,    -4,    -9,     1,     1,    13,     0,    -6,    -9,    -2,    -4,    -6,    -1,    -2,     5,    -6,   -19,   -28,   -21,    -3,    -7,   -10,   -10,   -11,    -4,    -6,    -4,    -4,     5,    -6,    -4,    -6,     1,     0,    -2,    -4,    -9,   -11,    -5,   -11,    -5,    -2,    -8,    -1,   -23,   -28,   -33,   -15,     8,    -5,    -7,    -3,     2,     1,    -2,    -5,   -12,    -9,    -9,    -6,     0,     2,     3,     8,    -4,     0,     2,    -7,    -5,     3,     3,     0,   -17,   -28,   -12,    -6,     0,     5,    -3,    -6,     4,     8,    -3,    -3,   -10,    -8,   -12,    -3,     0,     1,    -2,     7,     5,    -1,    -6,    -5,    -9,     6,    14,     0,   -16,   -12,    -9,   -11,   -14,    -2,     3,    -1,     2,     7,     2,    -4,    -7,    -1,   -11,    -2,     0,     0,    -3,     4,     7,     2,   -15,    -6,     2,    11,    18,     1,    -8,   -14,    -4,   -11,   -24,    -2,    -2,    -3,     9,     5,     9,    -7,    -9,     8,    -9,   -10,    -1,     0,    -2,     5,     5,    -8,   -11,    -6,    -2,     4,     9,     9,   -11,    -7,    -9,    -6,   -30,    -1,    -4,    -4,     7,    -4,     6,    -6,   -13,    -5,   -20,    -5,     0,    -2,    -6,     3,     3,    -6,   -10,    -3,    -1,     5,     9,     3,    -3,   -15,   -21,   -38,   -16,    -1,    -9,    -3,     4,    -5,     0,     1,    -5,    -8,   -15,     1,     1,    -1,    -5,    -1,    -2,    -9,   -11,    -8,    -7,     5,    10,     3,    -5,   -13,   -28,   -30,   -20,   -11,    11,     0,     8,    -4,    -1,     0,    -7,    -8,   -10,    -3,    -2,     3,    -5,    -2,    -2,    -4,   -12,    -8,    -4,    13,     5,    -4,     2,    -6,   -13,    -9,    -5,    -3,     1,    -1,     5,    -1,    -7,     2,     2,   -19,    -4,     0,     2,     2,    -1,    -6,     5,     9,   -14,    -8,    -7,     1,     6,    11,    -9,    -3,    11,     0,    -5,    -3,     2,    -6,     1,     4,    -8,     6,     2,   -15,     6,     2,    -1,     2,     0,    -2,    -3,    -1,   -18,    -4,    -9,    -6,     2,     7,    10,     9,     7,     8,    -8,    -6,    -3,     2,     7,     1,     1,     3,     3,    -2,     5,     7,     0,     0,    -1,    -3,    -6,    -3,    -8,    -4,    -4,     0,    -6,     7,    -1,     6,     7,    -2,     4,    -4,     1,     6,     8,     4,     2,     5,    -2,     1,     5,     4,     0,     1,    -2,    -7,     1,    -3,   -12,   -16,    -6,     6,    -2,    -5,    -2,     9,     6,    12,    17,    17,     4,    -9,    -8,    -4,    -2,    -6,     2,   -10,    -4,     1,     0,    -2,    -4,     1,     6,    -3,    -8,    -7,   -11,    -5,    -4,    -6,    -4,    -4,    -6,     0,    -1,     3,    -1,    -8,    -4,     1,     1,    -4,    -3,    -1,     1,     0,     1,     2,     2,    -1,    -3,     0,    -5,    -1,    -2,    -2,    -2,    -4,    -3,    -4,    -1,   -18,   -13,   -15,    -8,   -10,   -12,    -8,    -7,    -2,    -2,     2,     1,    -1,     1,    -2,     2,    -1,     0,    -7,   -10,    -1,    -2,     0,    -4,    -4,    -3,    -9,   -12,   -10,    -9,   -15,   -15,    -3,   -13,   -10,    -2,    -2,    -2,    -2,     0,     2,     0,     2,    -2,    -1,     2,     1,    -1,     1,    -2,    -2,    -2,    -3,     1,    -5,    -3,    -2,    -2,    -2,    -2,     0,    -2,    -5,    -4,    -2,    -1,     1,    -1,    -1),
		    71 => (   -1,    -2,    -2,    -2,    -1,    -1,     1,     0,     1,    -2,    -1,     1,     1,    -1,     2,     1,     1,     1,     2,     0,    -2,     0,    -1,    -2,    -2,     2,    -2,     2,    -1,    -1,     1,     2,     1,     1,     1,     2,    -2,     1,    -1,     1,    -1,    -1,     7,     2,     5,     0,    -3,    -2,    -2,     2,    -1,    -2,    -1,     1,    -2,     1,    -2,     2,    -1,    -1,    -2,     1,     1,     2,    -8,    -9,    -5,    -4,   -11,    -6,    -9,     0,    11,    -1,    -3,    -3,    -7,   -18,   -13,    -9,    -3,    -4,     0,    -1,     1,    -2,    13,     1,     1,    -4,    -4,    -2,    -8,   -12,   -13,   -17,    -1,     2,   -17,    -5,     8,     9,     9,     8,     9,    10,    -4,    -1,    -3,    -1,    -1,     2,     1,    -2,    11,    11,     3,     5,     1,    -1,     4,     0,     4,    -2,    -1,     5,    -9,   -13,    -2,     3,     6,    10,    -6,     8,    -4,     2,    -2,    -8,   -11,    -4,     2,     1,     6,     2,     3,     5,    -1,    -2,    -8,    -5,    -5,     1,     9,     0,     7,     8,     3,   -11,    -1,     6,     5,     5,     3,     2,    -3,    -9,    -2,    -5,    -1,     0,    -8,    -7,    -3,     4,     2,    -2,   -21,   -31,   -14,     1,    -3,    -6,    -4,    -2,     1,   -13,     8,    -2,     2,     8,     5,     2,    -1,     0,    -5,    -3,     1,    -2,    -9,    -9,   -11,     4,     4,   -10,   -20,    -9,     0,    -8,    -2,    -9,    -2,   -10,    -7,    -5,     5,     3,     6,    12,     4,    -3,    -5,     1,   -10,    -2,    -1,    -4,   -13,    -9,   -13,    -4,    14,     3,   -16,    -7,     2,    -3,    10,     9,     1,    -3,    -6,    -8,   -12,   -15,     1,     6,     8,    -5,    -8,    -1,   -11,     0,    -1,     0,    -7,   -11,    -8,    -1,     2,     8,     6,     1,   -10,    -5,    -5,     6,     2,    -1,    -9,    -8,   -14,   -20,    -8,    -3,     3,     9,    -4,    12,    10,    -4,    -1,    -4,    -8,    -5,    -6,    -6,   -10,    -6,     7,    -5,   -12,    -4,     2,    10,     3,   -10,    -3,     1,   -10,    -5,   -14,   -16,     7,     8,    -6,    10,     8,     9,    -1,     0,    -3,    -3,    -6,    -6,   -10,   -10,   -13,   -16,   -13,    -1,     3,     0,    -4,   -10,    -8,     1,   -12,   -10,    -5,    -7,     6,     8,    -5,     9,     6,    15,     2,     2,    -4,    -5,     0,    -2,     0,     0,   -10,    -5,    -2,     2,     9,     8,    -2,    -4,     2,    11,   -14,   -13,    -5,    -5,    -6,    -3,     0,    13,    16,    19,    -1,     1,    -1,     0,    -1,     5,     4,     2,     9,     9,    -4,    -3,    -3,   -14,    -1,    -2,     2,     3,   -19,   -18,   -11,   -10,   -11,   -17,   -11,    16,    13,    -1,     2,    -2,     1,     3,    -3,     6,     6,    -3,    19,    17,     6,   -10,   -16,   -13,     2,    -2,     9,    -1,    -8,   -15,    -6,    -9,    -7,    -3,    -1,    -1,     1,     0,     0,    -2,     1,    -4,    -6,    -5,   -10,     5,     8,    17,     1,    -6,    -4,    -1,    -2,    -1,     5,    -2,    -4,   -11,   -11,   -13,   -10,    -9,   -12,    -1,    -1,    -4,     1,     1,     1,    -6,    -1,     4,    -9,    -1,     7,     4,     3,   -10,    -1,    -3,     2,   -12,     0,    -5,   -10,   -20,   -13,   -19,   -12,   -10,    -1,   -13,    -7,    -2,     2,    -1,    -1,    -6,     0,     4,    -5,   -13,    -4,    -9,   -12,   -22,     3,     9,     2,    -1,     0,   -10,   -19,   -16,    -7,   -12,   -10,    -5,    -3,    -7,    -9,   -13,     5,    -1,    -4,    -1,   -11,    -9,   -14,   -17,   -18,   -29,   -22,   -25,   -11,    -3,    10,     2,     1,    -6,   -17,    -9,    -8,    -7,    -7,    -7,   -10,    -5,    -9,    -4,     0,    -2,     2,    -7,    -8,   -21,    -8,   -15,    -6,   -15,   -18,   -24,   -16,   -12,    11,     9,     1,    -2,    -9,    -4,   -10,    -7,    -1,     2,    -4,    -4,    -6,     0,    -1,     1,    -3,     4,     7,    -3,     3,    -5,    -7,     6,     6,     0,     3,   -13,    12,     9,     9,     6,    17,     2,     9,    -8,   -10,    -2,     4,    -6,    -4,    -1,     4,     0,    -6,     9,    12,     7,    11,     9,    -1,    -5,     2,    -4,   -10,    -9,     5,     6,    12,     1,    13,     4,    12,     3,   -16,    -9,    -5,    -2,    -9,     0,     4,     4,   -17,    -8,    16,    21,    13,     7,     2,    -7,   -12,    -7,     0,    -5,    -3,    20,     8,    -6,     3,     1,     5,     2,    -9,    -9,    -7,    -1,     1,     0,     2,     2,    -3,    -7,     3,     1,     8,   -10,   -15,    -6,   -16,   -13,     2,    -1,     0,     4,     2,     1,     2,    -3,     1,    -7,     0,    -4,    -5,   -11,    13,    -1,     1,     1,     0,    -4,     1,    -1,    -3,    -3,    -9,    10,     8,     2,    -4,   -17,   -15,     4,    -3,     6,   -10,   -26,   -12,    -9,   -13,    -9,   -13,    16,    17,     2,    -1,     1,    -2,    -3,    -1,    -2,    -5,    -3,    -3,    -6,    -7,   -14,   -11,   -22,   -10,   -17,   -12,   -25,   -17,   -12,   -18,    -5,    -4,    -4,     0,    -2,    -4,     0,     0,     0,     0,    -1,    -2,    -3,    -1,    -5,    -1,    -5,     0,     0,   -17,   -12,     6,     4,    10,   -17,    -5,    -4,     0,    -4,     0,     1,     2,     0,     2,     2,    -1,    -1,     0,     0,     2,     2,    -2,     0,    -2,     2,    -5,    -4,    -2,    -3,    -6,    -6,    -4,    -1,     2,     2,    -2,     2,    -1,     1,     1,     0,    -2,     2),
		    72 => (   -2,    -1,     0,    -2,    -1,     2,    -1,     1,     1,     0,     1,     1,    -6,    -5,     3,     2,     2,     2,    -2,     2,    -1,     2,     0,     2,    -1,     1,    -1,     0,    -1,     0,     0,     0,     0,     1,    -3,     0,   -11,    -7,   -11,   -14,   -10,   -14,    -6,    -9,    -3,    -7,    -9,   -20,   -14,    -4,    -4,    -4,     2,     0,     1,     1,    -2,     0,    -3,    -3,    -8,    -1,    -1,   -13,    -5,    12,    10,    -1,    -3,   -20,   -16,   -27,   -18,    -5,     0,    -4,   -23,    -6,    -8,    -3,     5,     2,    -1,     2,     0,     1,    -4,   -10,    -5,     2,     1,     0,     4,     4,     7,     0,   -11,   -25,   -19,   -21,   -21,   -17,   -19,   -16,   -19,   -14,    -9,    -4,     1,     1,     2,     1,     1,    -2,    -7,    -1,     1,    -5,     6,     6,     2,    -4,     8,     2,    -8,   -22,   -19,   -16,   -18,   -11,   -18,   -17,   -11,   -13,    -9,    -7,     1,    -2,    -8,    -3,    -2,     2,    -5,     0,     5,    -7,    11,    10,    11,     1,     6,    -6,     5,     0,    -8,    -1,   -22,   -22,   -16,   -10,    -6,   -11,   -14,    -5,    -8,    -3,    -2,    -4,    -2,     1,    -2,     2,     5,    12,     8,     2,     7,     9,     0,    -3,    -2,     6,    -2,   -10,   -11,   -12,   -12,    -6,    -5,   -11,   -11,    -9,   -14,    -5,    -4,    -4,     0,    -1,    -1,    -5,    -2,    -2,    -9,    -5,     1,     3,   -11,    -1,    -3,    -3,    -7,    -8,   -11,    -3,   -12,   -14,   -12,   -16,   -18,   -20,   -14,    -9,    -8,    -5,    -8,    15,    -3,     0,   -14,    -4,     3,    -4,     1,    -5,     5,    -5,    -6,     7,     7,     1,    -4,    -4,    -9,   -11,   -21,   -22,   -18,   -17,   -19,    -8,   -11,    -5,    -2,    -7,    -4,     5,   -16,    -3,     1,    -6,     0,    -1,     4,     1,     3,     1,    21,     6,    -3,    -9,   -12,   -10,   -13,   -13,   -26,    -7,    17,   -15,    -5,    -6,     0,    -5,    -4,    -2,   -19,     7,    -1,     0,     0,    -8,    -9,    -4,     2,    -3,     5,    13,    10,    -7,   -11,    -7,    -8,   -13,   -13,     3,    10,    -7,   -11,    -9,     0,    -1,   -14,    -6,    -7,    -6,    -6,    -4,    -6,     0,     3,    14,    -8,   -12,    -3,     4,     1,    -3,    -2,   -10,   -13,   -18,   -10,     1,    -2,   -10,   -19,    -2,    -2,    -2,   -17,    -2,    -1,     4,   -11,   -19,    -2,    -6,   -10,    -6,    -1,    -1,    -5,    -2,     5,    -3,    -2,   -13,   -10,    -3,     3,   -17,    -5,    -6,    -9,     2,    -2,    -3,   -13,    -1,    -3,    -4,   -15,   -20,    -5,    -8,   -14,    -8,    -5,     1,    -6,     5,     1,     2,    -6,    -7,     4,    12,    16,     3,    -4,    -3,    10,    10,     1,    -1,    -3,    -4,   -11,    -1,   -17,   -12,    -5,   -11,    -4,    -5,     0,     4,     3,     4,     6,    -1,    -7,     0,     5,    13,     7,    -2,    -4,     1,    20,    10,    -1,    -4,    11,    -9,    -2,    -1,    -3,   -10,    -6,    -2,     3,     0,     9,    14,     5,     6,     0,    -3,    -3,     1,     7,     2,    -7,   -10,     0,     3,     6,    12,     1,     0,    12,    -3,     7,    -9,     1,    -3,   -16,    -4,     3,     9,     1,     7,     6,     5,    11,     6,     1,     5,    -1,     5,     5,     5,     4,     7,    -3,    12,    -2,    -1,    17,     3,     9,    -5,     9,     1,    -4,     2,     6,     8,    -1,     2,     9,     8,     9,     7,     9,    13,     8,    10,    -4,     2,    -1,    -5,   -13,    11,    -1,     1,     7,     6,     5,     4,    13,    -1,    -7,     2,     7,     8,    -5,     3,    -4,     6,     4,     1,     8,     5,     2,     8,     6,     9,    15,     8,   -10,     8,     0,    -9,     1,    14,    -2,     9,     6,     3,    -1,    10,     3,    -2,    -8,    -6,    -3,     7,    -1,    -1,    -4,    -6,    -7,     0,     9,    15,     9,     5,     9,    18,    -1,    -4,     3,    10,     1,    -3,     2,    -5,     5,    -2,     0,    -1,    -2,     1,     2,     0,   -12,   -18,   -15,   -15,   -13,    -4,    -7,    -4,    -4,   -13,     7,    -1,     2,    -1,    -2,     6,     4,     3,    15,     0,    -1,    -2,     9,    -8,     3,    -6,    -7,    -7,   -23,   -35,    -5,    -7,   -12,   -14,   -15,   -21,   -21,   -10,    -9,     0,     2,     2,    -1,    -1,    -1,     5,     3,    -7,    -7,    -8,   -11,    -4,    -5,   -10,    -8,   -22,   -34,   -31,    -9,    -6,   -12,   -19,   -23,   -17,   -17,   -14,   -22,     0,     2,    -2,     2,    -2,    -3,    -5,    -6,   -10,    -1,    -1,   -15,   -16,   -29,   -25,   -33,   -26,   -31,   -30,   -21,   -22,   -20,   -22,   -19,   -27,   -21,   -12,   -21,     2,     0,     2,    -7,    -2,   -24,    -6,   -15,    -4,     2,   -11,     2,    -7,   -45,   -32,   -28,   -23,   -27,   -29,   -25,   -24,   -23,   -24,   -19,   -19,     3,     8,     7,     0,    -1,     0,    -1,     1,    -6,    -4,    -1,    -3,   -18,   -24,   -26,   -16,   -25,   -24,   -17,   -20,   -21,   -16,   -12,   -20,   -21,   -18,    -5,    -5,     0,     4,     5,     1,     0,    -2,    -2,     1,     0,    -8,   -13,   -12,   -18,   -23,   -17,    -6,    -7,    -8,   -12,    -4,   -10,    -8,    -4,   -14,    -7,    -5,    -9,    -2,    -2,     0,     1,    -1,    -2,     1,     1,    -2,     0,    -2,    -2,    -1,     2,    -3,    -6,    -1,    -3,    -9,    -5,    -1,    -4,    -4,    -7,    -4,    -5,    -6,    -5,    -2,     2,     2,     0,     0),
		    73 => (    2,     0,    -2,     1,    -2,     2,    -1,    -2,    -2,     0,     1,     2,    -3,    -2,    -4,     0,    -1,     2,    -2,    -2,     1,     1,     0,     1,     1,    -2,    -1,     0,    -1,     2,     2,    -1,     0,     0,    -2,     0,     0,     0,    -3,    -3,    -2,    -3,    -7,    -5,    -3,    -3,    -1,     1,     0,     1,     1,     0,    -1,    -1,     2,     0,    -1,     0,    -2,    -1,    -1,     1,     1,    -3,    -4,    -7,   -20,   -19,   -19,    -4,    -4,    -1,    -3,    -3,     1,     0,    -6,    -1,     0,    -4,    -2,     0,    -1,     0,    -2,     0,     0,     0,     0,    -4,    -2,    -1,     3,     1,    -3,   -11,    -7,   -10,   -14,   -16,   -15,    -6,    -5,    -2,    -4,    -5,    -8,   -10,     0,     0,    -2,     0,    -1,     0,     2,     1,     0,    -2,    -4,   -14,   -11,   -26,     3,     9,    -2,    -2,     8,     2,     0,    -2,    -1,     0,    -2,     8,    16,   -11,   -11,    -9,    -1,     0,    -1,     0,     2,    -2,     1,    -8,    -6,    -8,   -19,   -20,    -8,     9,     7,    -9,    -4,    -5,     0,    -6,    -5,    -8,     1,    -9,    -4,    -7,    -7,   -23,    -7,    -2,     0,     1,     5,     4,     0,    -7,     3,    -4,    -3,     6,    13,     3,    -2,     5,    -3,     3,     4,   -10,    -4,   -12,     1,     0,    -7,    -1,    -6,   -11,   -16,    -5,     2,     2,     2,    -1,     2,   -23,   -18,    -8,     2,     1,    -1,   -10,     3,    16,     1,    -7,    -8,    -3,     0,    -3,    -4,    -7,    -4,   -12,   -17,   -10,   -13,    -2,     0,    -1,    -2,    -4,     0,   -16,   -11,     1,     2,     2,    -5,    -4,     8,     7,    -2,    -4,     2,    -5,    -4,    -2,    -2,    -3,     0,    -6,   -30,    -9,   -20,     2,    -2,    -3,     2,    -4,    -9,    -9,    -4,     5,    -2,     3,     6,    12,     8,    -3,    -3,    -7,     4,     7,    -5,     1,     3,    -2,     4,     2,   -24,    -9,   -12,   -10,     1,    -6,    -1,    -3,    -5,    -9,    -4,    -9,     5,     1,     4,    12,     7,   -11,   -14,    -5,    -7,    -5,    -8,     3,    10,    -8,     3,    -1,   -23,   -19,   -17,    -8,    -2,    -8,     0,     5,    12,     8,     3,     0,    11,     2,   -11,   -13,   -44,   -17,    -7,    -9,    -7,    -2,    -6,     2,     7,    13,    -1,     6,   -19,   -13,    -8,     2,    -1,    -5,    20,     4,    14,     9,     1,   -16,   -13,   -22,   -22,   -30,   -23,    -3,     1,    -4,    -4,    -9,    -6,    -2,     4,     9,     8,     7,   -12,     3,    -6,     0,    -1,    -8,    -9,   -12,   -14,   -11,    -9,   -34,   -30,   -23,   -12,    -7,     2,    12,    12,    -7,     1,    -2,    -4,     1,    -2,    -4,    -4,    -2,   -14,    -9,   -11,    -4,     0,     3,     6,    -5,   -10,   -26,   -25,   -30,    -4,     8,     4,    -5,     0,     7,    -1,     3,    -2,     6,     0,    -9,   -12,    -6,    -7,     1,    -8,   -18,   -11,    -4,    -2,     1,     0,    -3,   -13,   -28,   -36,    13,    12,     2,     3,     5,    11,    10,     9,     2,    -2,    -2,     2,    -2,   -14,    -9,   -17,    -7,    -8,   -11,    11,    -3,    -1,     2,     5,    -4,    -6,   -10,    -4,    -4,     6,     9,     9,    10,     9,     7,     8,    -2,    -1,    -6,    -2,    -7,   -17,   -11,   -11,     2,    -5,    -7,    -3,    -4,     2,     2,     5,     4,   -12,   -13,    -6,    -9,    -3,     4,    14,     5,    14,    13,     3,   -13,    -9,     1,    -3,    -1,   -17,   -12,    -8,    -6,   -19,    -7,    -2,    -1,    -5,    -3,     1,     5,   -12,   -22,   -24,    -7,   -12,    -1,     5,    10,    13,     2,     1,    -6,    -6,   -11,     4,    -2,     2,    -6,    -6,   -16,   -19,    -3,    -2,    -2,    -2,    -6,     1,    -1,   -18,   -17,   -20,   -18,   -24,   -17,   -21,    -8,   -16,    -6,   -11,    -6,     8,     5,    10,     1,    -8,     3,    -8,   -17,   -19,    -1,    -9,    -3,     1,    -6,     4,    13,    -5,    -2,   -19,   -31,   -32,   -48,   -64,   -47,   -38,   -13,    -2,    -6,    -2,     9,    12,     7,     3,    -5,    -8,   -22,   -18,   -12,    -3,     2,    -3,    -2,     9,    20,    12,     0,    -2,   -12,    -2,   -10,   -10,   -15,   -10,    -8,     0,     4,    -1,     0,     6,     0,     6,    -2,    -6,   -15,   -11,    -4,    -6,     2,    -2,     1,     3,    11,    21,    20,    14,     9,     8,     5,    11,     5,    -4,     3,     3,     3,     5,    -2,    -3,    -1,    -6,    -4,   -11,    -7,   -12,    -7,    -1,     0,     2,     2,     2,    -5,    14,    14,    13,    11,     2,    -4,     5,     0,     8,    14,     0,     7,   -14,     3,    -1,   -10,     7,     2,    -4,    -3,   -13,    -8,    -1,     2,    -2,    -1,     3,     9,    18,    -3,     9,     8,     1,     1,     7,     8,     5,     6,    -1,    -3,    -5,     4,   -26,    -7,     5,     6,     9,    10,   -16,    -4,    -6,     0,     2,    -1,     3,   -10,     0,    27,    17,    15,     6,     8,     1,    -4,     2,    -4,   -10,    -4,    -4,   -10,   -26,    -5,    -8,   -17,    -6,   -20,   -12,    -7,    -9,     2,     1,     2,     0,    -8,   -16,     0,     2,    -3,    -3,   -13,     0,     2,    -5,     2,     0,   -13,    -2,     6,     5,    -6,    -3,    -5,     2,    -2,    -2,    -1,     1,     0,     2,    -2,    -2,     0,    -2,    -6,    -2,    -1,    -2,   -15,   -13,   -10,    -7,    -9,    -9,    -9,     1,    -1,    -5,   -11,    -9,    -2,    -8,     0,    -2,    -1,     0,    -1),
		    74 => (   -1,     0,    -2,     0,     0,     2,    -1,     1,     2,     2,     1,     2,    -2,    -8,    -2,    -1,    -2,    -1,    -2,     2,    -2,    -2,    -1,     1,    -1,     2,    -1,    -1,     0,     0,     3,    -2,     2,     2,   -10,    -9,    -3,    -8,   -15,    -9,   -18,   -11,     5,   -27,   -25,   -17,    -5,    -1,   -12,    -2,     0,    -4,    -2,     1,     1,    -2,    -1,    -2,    -4,   -10,   -15,   -10,    -5,   -14,    -9,    -9,   -24,   -31,   -24,    -5,     3,    -8,   -14,   -11,   -16,   -21,   -21,   -13,   -14,   -17,    -4,   -10,     2,    -2,    -2,     0,    -7,   -19,   -32,   -11,   -12,    -1,   -22,   -25,   -15,   -21,   -36,   -12,     4,    -2,    -9,   -14,   -19,    -6,    -5,   -10,    -6,   -18,   -21,    -9,    -1,     1,     0,     0,    -4,   -28,    -3,     1,     1,     4,    -1,   -14,   -11,   -10,    -3,     7,     9,     4,     2,     6,    10,     0,    -5,     2,    21,     1,    -2,    -4,   -19,    -6,    -1,     1,    -7,   -13,     2,     6,     4,    17,     9,     7,     7,    -3,     6,    10,    16,     4,    -1,    12,     4,    14,    -3,     9,     9,    16,    16,     9,   -18,     0,    -2,     1,    -6,    -4,    11,     7,     3,    17,    14,    16,     9,     6,     3,    16,    20,    26,    16,     3,    -7,     0,     6,     1,    -2,    15,    20,     6,     4,   -11,     0,   -10,    -9,     5,    11,     5,    11,    18,     8,    37,    24,    33,    18,    20,    18,    17,    10,    12,     4,    13,     6,    -5,    -4,     2,     8,    -8,    21,   -15,   -11,   -12,    13,     6,     6,     1,    14,     7,    -1,    31,    18,    20,     3,    -4,    -2,     5,    -6,    -6,    -6,    -2,     3,     2,   -14,    -5,     0,     5,    10,   -16,     1,    -5,    10,    -8,     1,    -8,   -11,    -5,    -5,    -1,     6,   -13,    -5,     2,    -4,     2,   -10,     5,    -2,    -3,    -3,    -4,   -17,     0,    -3,   -10,   -10,    -8,     2,    -6,     6,    -5,    -5,   -12,   -20,    -9,   -10,     3,    -5,   -16,     0,   -13,   -11,    -6,    -5,    -1,   -13,     0,   -16,    -9,    -4,   -10,   -22,    -6,    -2,   -13,     2,   -11,     6,    -8,   -11,    -9,     7,   -15,     2,    -7,   -14,    -4,    -2,    -4,    -8,    -3,     2,     9,   -11,   -10,   -27,   -11,    -7,   -16,   -26,    -6,   -11,   -21,    -2,     2,     2,    -9,   -15,    -4,    -2,   -10,    -2,     2,    -8,     4,    16,     8,   -15,     0,     3,     6,    -4,    -7,     0,     8,    -4,   -10,     2,    13,   -10,   -17,    -1,    -5,   -14,   -13,   -15,    -2,     1,    15,     8,    -6,     5,    14,    18,    -2,     5,     2,     0,     7,     9,    -2,     1,    -8,    -9,    -4,     2,     7,    -5,    -2,    -2,     8,   -25,   -17,     0,     0,     0,    23,    13,     8,    13,     9,     6,    -4,    -5,    -2,     3,     3,    -4,    -2,   -11,   -13,    -3,    -2,    -1,    10,   -14,    -2,    -2,     2,    11,     2,    13,    -1,     8,    11,    13,     7,     2,     2,    12,     8,     3,    -1,     6,    12,    -3,    -6,     1,     1,    12,     7,    -5,    -1,    -9,   -14,     1,     0,   -16,     4,    -6,    -6,    -6,    -5,     1,    -1,     7,     7,     1,     0,     3,    -2,     4,     5,     3,     6,    12,     8,     9,    -2,     5,     2,    -8,    -6,     1,    -1,   -10,   -13,     0,     1,    -7,    12,     2,    -2,   -13,    -5,     1,    -9,    -2,    -9,    10,    -2,    -4,     3,     1,     9,     4,    17,     5,   -20,    -4,    -7,   -11,    -2,    -4,     1,     2,     9,     5,     2,   -11,    -5,   -13,    -9,     5,    -6,     1,    -6,    -8,   -16,    -5,    13,    21,    13,     8,    14,     9,    -5,    -9,   -13,     1,   -10,   -14,    28,    -7,    -5,    -8,   -14,    -5,   -12,   -15,   -15,    -1,     1,     5,     7,     3,   -16,     0,     6,     7,     5,     9,     1,     3,    -1,    -4,   -10,     2,    -3,    -7,     7,    -9,   -13,   -15,   -16,    -9,     7,     1,     1,     0,    -2,     1,     6,     9,    -2,    10,    10,    15,     9,     4,    -3,   -15,   -17,    -7,    -2,    -4,    -1,   -11,     9,     6,    -6,   -10,    -8,     2,     4,     0,     5,   -11,    -5,    -3,     6,     7,     6,    -2,    13,    28,    21,    22,     7,    -5,   -24,   -16,     1,    -4,    -4,    -4,   -13,   -29,   -15,     0,     5,    12,    -5,    15,     2,    -3,     0,   -11,    -6,    11,    10,    -1,    21,    24,    27,    17,    14,     1,    -1,    -5,    -3,     2,     2,    -1,   -19,   -25,   -46,     8,    13,    20,    12,    22,    17,     7,     0,    -4,    -7,     4,    -2,    10,    23,    22,    10,    -9,    10,     0,    14,    -5,     0,     0,     1,     1,    -7,   -24,    -4,    19,    21,     6,    15,     2,    17,    -5,    -1,    -1,   -16,    -7,    -9,    12,    21,     0,    -7,    -4,    -1,   -13,    12,   -12,    -1,     0,     0,    -7,    -1,    20,    28,     9,    -8,    -5,     2,    10,     9,   -10,     6,   -13,     4,     2,    -3,    -3,    -2,    -3,    -5,    -5,     2,    -5,   -13,   -10,     2,     1,    -2,     0,   -18,    31,    26,    15,    -5,   -11,   -18,   -31,    -6,    -9,   -10,    -6,   -23,   -24,   -16,    -4,    -1,   -18,   -37,   -32,    -8,     2,    -2,     2,     2,     0,    -2,     1,    -1,    -4,    -1,   -11,   -12,    -8,    -9,   -13,   -15,   -12,    -4,    -9,    -4,   -20,   -29,   -23,   -14,   -15,    -7,   -10,     1,     2,     0,     0,     0),
		    75 => (   -2,     2,    -2,    -1,     0,    -1,    -2,     1,    -1,    -2,     0,     0,     2,     1,     1,    -2,     2,     0,     2,     0,     2,     1,     0,    -1,     2,     1,    -2,    -2,    -1,     0,    -2,    -1,    -2,     2,     0,     0,     2,     1,    -2,    -3,    -4,    -8,    -6,    -4,    -3,    -8,    -5,     0,    -1,    -3,     1,     1,    -2,     2,    -1,     1,     1,    -1,    -2,    -2,     0,     1,    -6,    -4,   -12,   -13,   -15,   -15,    -8,   -10,   -23,    -4,     3,     3,    -2,     7,    13,     1,     0,     4,    -6,    -1,     2,     0,     1,     0,    -3,     3,     7,   -10,   -12,   -12,    -7,    -4,    -4,    -6,     2,     4,     7,     9,     7,    -1,    -8,    -6,     3,     8,     2,     7,     3,     2,     3,     2,     2,    -2,     0,     6,     0,    -1,     6,    10,     3,    10,     0,   -12,    -7,    -1,     4,    10,    11,     1,    -1,    -8,    -2,     1,     5,     7,     5,     8,    -5,    -7,    -2,    -1,     1,     1,    -7,     0,    10,     5,     6,     1,    -2,    -9,   -11,    -2,     0,    -3,    -1,     0,    -1,    12,     9,     0,     8,     8,     7,     6,    -6,    -6,     1,    -2,   -11,    -7,     4,     6,    13,     4,     1,    -1,     0,    -6,    -7,    -3,    -1,     0,    -2,    -6,     3,    13,    14,     9,     7,     4,     7,     7,     5,     3,    -2,     1,     1,    -9,     2,    16,     2,     3,    -6,    -3,    -4,    -2,    -4,    -6,    -1,    -6,    -1,    -2,    -4,     1,     6,    -3,     8,     7,    15,     8,     6,     7,    -2,    -7,    -8,   -14,     3,     1,     1,     2,    -5,     1,     0,     7,     4,     5,    -1,    -8,    -8,   -12,     2,     3,    -4,     1,    12,    15,     7,    11,     7,     4,    -1,    -4,   -18,   -12,     1,     3,     1,     1,    -5,    -4,     6,     8,    12,     9,    -4,    -5,   -10,   -10,    -4,     0,     5,    12,    15,    14,    12,     2,    10,     3,     1,    -1,    -3,   -18,     0,     0,    -1,     5,    -5,     2,    -1,    12,    16,     2,     7,     0,   -11,    -4,     1,     7,    13,    20,    19,    15,    14,     7,     1,    -7,     2,    -3,    -2,   -12,     4,     0,     3,     5,     6,    -2,    -5,    11,     9,     1,     7,    -7,   -10,   -16,    12,    11,    19,     7,     9,     9,    12,    11,     2,    -8,     1,     1,     0,   -14,     4,     6,     7,     7,    12,     8,    -7,     0,     3,     1,     2,    -4,   -10,    -1,     6,    12,     7,     0,    -3,     8,     5,     5,    12,    -9,    -2,     0,    -2,   -15,     0,     5,     5,    10,     7,    11,    14,     6,     5,    -4,     0,   -10,    -6,    -5,     0,    10,     9,    10,     0,    -6,    -7,    -1,     9,    -8,     2,     0,    -3,   -20,    -2,     3,     7,     9,     8,     6,    15,     2,     3,     1,     0,    -8,    -4,     4,    14,    11,    10,     8,     6,    -5,    -9,    -9,    -6,     1,     2,    -3,    -5,    -2,     4,     7,    -1,     3,     8,    12,    14,    -1,    -1,     1,     7,     2,    -1,     6,     8,    12,     6,     6,     3,     0,     2,   -10,    -6,   -13,    -1,    -4,    -9,    -1,     5,    18,     5,     3,     7,     8,     7,    -9,     1,     3,     2,     6,    -6,     2,     0,     2,    10,    18,     8,     1,    -5,   -10,    -8,   -16,    -2,    -1,    -7,     4,     6,    17,    11,    10,    13,    11,    -4,    -5,    -8,     0,     8,    -6,     1,    -2,    -2,    -1,     7,     5,     9,     2,    -2,   -11,   -17,   -18,     0,     1,   -11,     2,     3,    15,    11,     9,    14,    11,    -1,   -10,   -17,     4,     6,     0,    -1,    -5,    -6,    -8,    -2,     0,    -1,     4,     5,    -8,   -21,   -12,     3,    -3,     8,     1,     3,     7,     8,    15,    11,    -1,    -6,    -6,    -9,     5,     0,     2,    -5,     2,    -3,     1,     2,    -1,    -1,     7,     3,    -8,   -23,   -10,     2,    -1,     5,     5,     4,     3,     8,    10,    13,     0,    -5,    -8,     2,     1,    -5,    -4,    -3,     1,     7,     7,    -3,     4,     4,     8,    -9,    -2,   -16,    -1,     0,     0,     2,     1,     3,     7,     9,    12,    12,     9,     0,     5,     3,     2,     0,    -3,    -1,    -1,     3,     8,     9,     1,     3,     2,   -10,    -1,   -10,    -2,    -2,    -1,   -11,    -1,     4,     2,     8,     6,    13,     7,     3,    12,     6,     2,     1,     1,    -4,    -6,    -5,     2,     3,    -6,    -4,    -5,   -13,     1,     9,    -2,     0,     0,     3,     0,    -6,    -1,     5,    10,     6,     4,     0,     6,     5,     5,     4,    -4,   -15,   -10,    -6,    -5,    -3,   -10,    -6,   -10,    -3,     4,     7,     1,    -2,    -2,    -3,     0,    -8,    -4,     7,     3,     3,     6,     7,     5,     2,    -4,     2,     0,    -9,    -7,    -3,    -8,    -9,    -7,    -5,    -4,     3,   -16,    -6,     1,     2,    -1,     2,     8,   -15,   -12,    -1,     4,    -5,    -9,     9,     5,     5,     2,     0,     4,     6,    10,     7,    -2,     6,     3,    11,     3,     1,     0,    -1,     0,    -1,    -2,     0,    -8,   -12,   -16,   -18,    -3,    -1,    -4,    -3,     9,    -2,     3,     8,     5,     5,     2,    -4,    -2,    -8,    -6,     2,    -9,     0,     0,     2,    -1,    -1,    -2,    -2,    -2,    -4,    -3,    -1,     0,    -2,     0,     2,     0,    -4,    -2,    -4,    -2,    -1,     1,    -2,    -6,    -3,   -13,    -9,    -4,    -1,     2,     2,    -1),
		    76 => (    1,    -1,     2,    -1,     0,    -1,    -2,     1,     1,     2,    -1,     1,     1,     1,    -1,    -2,     1,     1,     1,    -1,     2,    -1,     1,     0,    -2,     1,    -2,     0,    -1,    -2,    -1,    -1,    -1,     2,     3,     4,     8,     4,     3,     5,     4,     3,    -2,    -3,    -6,     1,    -1,    -1,    13,     6,     2,     4,     2,     1,     0,     1,     1,    -1,     3,     2,    11,     4,     0,     8,    10,     1,    -3,     0,     0,     2,    -6,    -3,    -3,     4,     0,     3,     5,    17,    20,    16,    15,     7,    -2,    -1,     1,     0,    -5,    -5,    -1,     0,     1,    -2,    -2,    -1,    -4,    -2,   -15,   -15,   -15,    -8,   -10,   -12,     4,    15,    16,    10,     4,    15,    15,     1,   -12,    -2,     2,     2,    -4,     1,     5,     3,    -5,    -7,    -8,    -1,    -4,    -7,   -14,   -18,   -20,   -15,    -7,    -8,    -6,     2,     2,    12,     1,    14,     5,    -4,     8,     9,    -2,    -1,    -6,    -7,     5,     2,    -3,    -4,    -3,    -2,    -9,   -12,   -13,   -12,    -9,    -4,    -6,    -2,     0,     1,    -4,     4,     8,    12,    14,    13,    16,     9,    -2,    -1,     1,    -2,     2,     3,    -4,    -2,    -7,    -2,    -8,    -8,    -5,    -8,   -16,   -17,   -14,    -3,    -3,     4,     0,    -4,     2,    11,    14,     8,     6,    14,     2,    -1,     1,    -1,     7,     3,    -8,    -2,    -1,     5,   -11,   -12,   -11,   -19,   -13,   -19,    -6,     1,     3,    -5,    -5,     2,    -6,    -6,     4,     8,     6,    15,     0,     0,    -1,    -3,     8,     1,   -13,    -6,    -4,    -2,   -15,   -16,   -19,   -18,   -15,   -11,     3,     2,     5,     1,     0,    -4,    -5,    -3,   -14,    -7,    12,    -8,     1,    -2,     0,    -6,    11,    -1,   -12,    -2,     3,    -2,   -14,   -16,   -18,   -18,   -10,     4,     5,     3,    -1,     2,    -3,    -5,    -5,   -10,   -12,    -8,    -6,    -4,    -1,    -2,     0,    -4,     8,    -3,    -8,    -2,    -2,   -12,   -26,   -20,   -14,    -3,    -1,     5,    -5,    -6,   -13,   -17,    -3,    -4,    -9,   -10,    -8,    -7,    -6,    -8,     1,    -2,     3,    -6,     3,     2,   -13,   -12,   -11,   -25,   -15,   -14,    -6,     1,     6,     0,    -6,   -20,   -25,   -16,   -16,    -9,    -7,    -9,   -13,    -2,    -3,    -4,    -3,    -1,    -3,   -10,     2,    -4,   -10,   -13,   -15,   -15,   -17,     1,    -5,     5,    -2,    -4,    -6,   -14,   -22,   -16,   -13,    -8,    -4,    -5,    -1,    -3,    -8,    -3,     2,     2,    -1,    -6,    -2,    -2,    -8,    -9,    -1,    -5,    -5,    -3,     4,     6,    -4,     2,     1,     0,    -4,    -5,    -3,   -16,    -9,    -2,    -1,     0,    -9,    -3,     0,     0,     1,    -5,    -6,    -7,    -5,     1,     8,    -6,     2,    -4,     6,     1,     2,    -7,     4,     0,    -2,     1,     1,   -10,   -18,   -15,    -2,     1,    -4,    -5,     0,     0,    -5,    -3,    -7,    -9,     5,     4,    -4,     2,    -5,     4,     9,    -1,    -3,    -4,    -1,     4,     1,    -6,   -11,   -12,   -16,    -7,    -4,    -3,    -3,    -7,     1,     1,    -4,    -6,     2,    -8,    -3,    -2,     2,     1,     0,     1,     5,     3,     1,     3,    -2,    -6,     3,     1,   -10,   -15,    -9,    -4,    -6,     1,    -5,    -3,    -2,    -2,    -6,   -10,    -3,   -11,    -8,     1,     3,    -2,    12,    -6,    -4,   -11,    -7,    -5,    -7,   -10,     9,     6,     1,    -9,    -3,    -5,    -7,    -5,    -6,   -12,     2,    -2,    -2,    -2,     8,    -4,    -9,    -5,     0,     2,     0,    -4,   -10,    -7,     0,     4,     0,     0,    11,    16,    11,     0,    -4,    -7,    -4,    -1,   -12,    -2,     0,    -2,     1,    -6,     5,    -5,    -7,     1,    -9,     4,    -3,   -10,    -3,   -13,     0,     7,     3,     5,    13,    10,     9,     1,   -10,    -7,    -2,     0,    -1,    -5,    -2,    -1,    -3,    -7,     7,     0,    10,     5,    -3,    -2,     0,    -4,    -4,     0,    13,     2,    -4,    -6,     0,     2,     0,    -5,    -8,    -8,     1,    -1,    -2,     0,     2,    -2,    -7,    -6,     3,    -1,     0,     1,     8,    -8,     5,    10,     9,     6,     4,     1,    -2,    -7,    -7,    -9,   -12,   -11,    -8,    -3,    -1,    -2,     1,    -2,     0,     0,    -3,     1,    -3,    -5,   -17,    -5,     8,    -3,     1,     9,    14,     6,    -9,   -10,    -5,   -11,    -9,   -10,   -10,    -2,    -2,    -7,    -5,    -7,     1,     2,    -2,    -2,     1,    -6,    -8,    -3,   -10,     6,     5,     2,     5,     8,     8,     2,    -2,    -5,    -2,   -15,   -12,    -9,    -1,    -3,    -1,     1,    -5,    -6,    -2,     1,     1,     2,    -1,    -1,    -3,    -5,    -2,    -3,    -7,    -6,    -3,    -5,    -3,    -6,    -2,    -2,     3,     0,    -1,    -7,    -2,    -4,    -3,     2,     0,    -3,     1,    -1,    -2,     2,    -2,    -2,     0,    -9,   -10,   -11,    -6,    -4,    -2,     0,     0,    -2,    -2,     1,    -3,    -1,    -2,    -3,    -8,    -3,    -2,    -4,     0,    -1,     1,    -2,     2,    -2,     0,    -1,    -2,    -4,    -4,    -3,    -2,     0,    -5,    -4,    -2,     0,    -1,     0,    -2,     1,     0,     1,    -5,    -2,    -4,     0,     0,     2,    -2,     2,    -2,     1,     2,     2,     1,     2,    -2,     2,     2,     2,     1,     1,    -1,    -1,    -3,     0,    -1,    -3,     1,    -1,    -2,    -4,     1,    -1,     0,    -2,     0,    -2),
		    77 => (    0,    -1,    -1,     1,     1,     0,    -2,     2,     0,     0,    -1,     2,    -1,     2,     1,     1,     1,     0,     0,    -2,    -2,    -2,     2,     1,     0,     0,     2,     0,     1,     1,    -1,     0,     0,    -1,     0,     2,     1,    -1,    -3,     0,    -1,    -2,    -3,    -9,   -11,    -7,     2,     2,     2,     0,     0,     0,     1,     0,     0,     2,     1,     2,     0,    -2,     0,     2,    -1,    -3,    -1,     0,    -6,    -4,    -1,    -1,    -2,    -2,     0,     1,    -3,     0,     0,    -1,     0,    -2,    -1,     0,    -1,     2,    -1,     0,    -2,    -2,    -2,    -1,    -1,     1,    -6,    -6,    -6,    -7,    -4,    -6,     1,    -7,    -9,   -17,    -5,    -9,    -5,    -5,    -9,    -2,    -4,    -2,    -2,     2,     1,     0,     1,    -1,    -7,    -3,    -6,   -17,   -14,   -12,   -16,   -24,   -28,   -21,   -15,   -28,   -20,   -23,   -22,   -13,   -14,    -5,   -19,   -11,    -7,    -5,    -2,    -2,    -2,     2,    -3,   -10,    -2,    13,    11,     8,    18,    17,     0,     7,     3,     6,    -4,     0,    -2,    -9,    -1,    -6,   -10,   -21,   -21,   -15,   -20,   -17,    -5,    -2,     2,     0,    -1,    -6,    -4,     7,     9,    13,    14,     0,     3,     8,    12,    13,    16,     4,    13,    10,     7,     8,     9,     2,     6,    -1,    -3,    -6,     0,    -5,     0,     2,    -3,    -2,    -6,    -5,    -6,    10,    -3,     2,    -2,     9,    15,    15,     6,     9,     6,    14,     2,     5,     7,    -1,     1,    -2,     2,    -3,    -4,    -3,    -7,     4,     0,    -4,    -4,   -11,   -10,    -8,   -14,   -12,   -14,    -1,     2,    -4,     2,     3,    -2,     6,    -3,     0,    -9,    -5,   -11,   -10,   -10,    -4,    -7,    -8,     0,    -1,    -3,     3,     1,    -8,   -14,   -11,   -23,    -7,   -14,    -9,    -7,   -11,    -6,   -10,     1,   -11,     0,    -2,    -9,    -6,    -7,    -9,    -8,    -3,    -8,     5,    -1,    -4,    -9,    -8,     0,   -10,     0,    -6,   -11,    -6,   -13,    -7,   -20,   -24,   -25,    -7,    -5,     2,    -4,    -6,    -1,   -17,    -4,   -14,    -9,    -5,   -10,     4,    -1,    -2,    -8,    -1,    -7,    -8,    -8,   -15,   -20,   -17,   -26,   -17,   -28,   -17,   -13,    -5,     0,    -4,    -6,    -7,    -5,    -5,     7,     9,    -7,   -16,    -8,     7,     0,     1,    -4,     2,     0,    -7,   -11,   -21,   -17,   -24,   -16,   -20,   -16,   -10,    -9,    -3,    -1,   -12,   -15,    -6,    -7,     2,     3,    -3,    -1,    -1,    -5,     7,     2,    -1,     4,     0,    -3,    -8,    -5,     1,    -9,    -2,    -7,    -4,    -4,     0,    -1,     2,     5,    -6,     1,    -3,     8,     9,    -3,   -10,    -8,    -1,    -9,    -8,    -2,    -1,     0,    -3,     6,     0,     4,     9,     0,     1,     3,     5,     8,     5,     5,     5,     5,     1,     5,    17,     0,     2,     4,   -17,   -10,    -6,    -6,     2,     0,     0,    -4,     1,     8,     7,     6,    10,     9,    -3,     4,    -1,    -4,     1,     0,     4,    11,     7,    -2,    -3,    -8,     2,    -6,   -20,   -20,   -13,    -2,    -5,     2,    -2,    -5,    -6,     2,     1,    -2,   -12,     0,    -1,    -1,    -8,    -1,     2,     2,     9,     4,     0,    -1,    -3,     2,    -4,   -12,   -16,   -18,   -11,    -8,    -7,    -1,    -1,    -6,    -5,    -9,    -4,     7,    -9,    -4,    -2,    -4,     6,     0,    -5,     4,    -3,    -8,    -8,    -1,    -1,     6,    -2,     2,    -3,     3,     5,    10,   -13,     1,     1,    -2,    -6,     0,    -6,    -7,    -3,     0,   -11,    -7,     7,     3,    -5,    -3,    -3,   -20,   -13,    -2,     1,    -7,    -9,   -11,    -9,    -3,     7,    13,   -12,    -1,     1,     2,    -3,     5,    -8,    -2,   -15,   -16,    -4,    -7,     1,    -7,    -6,    -3,   -10,   -27,   -11,    -1,    -3,   -21,   -27,   -13,   -15,    -7,     9,    -6,    -4,     2,     3,     3,    -2,    -7,    -3,    -5,   -10,    -8,    -5,     0,     6,    -7,    -6,    -5,   -11,   -16,    -8,   -21,   -20,    -8,   -11,   -13,    -6,   -15,   -17,    -4,    -2,    -1,     1,    -1,     0,    -5,     5,     0,     2,    -4,     1,     1,    -1,     8,     4,    -6,    -3,    -8,    -3,   -12,    -9,   -17,   -11,    -5,    -4,    -8,    -8,    -3,     1,     1,    -1,    -3,    -3,    10,     0,    -4,     3,     5,    -1,     0,     1,    -1,     5,   -12,    -1,     6,    -1,    -6,   -15,   -20,   -13,    -3,     0,   -12,    -4,    -6,     1,     1,    -1,    -4,   -17,    -1,   -11,     2,    -1,     0,    -6,    -4,    -2,     0,     8,    -5,    -5,   -14,   -15,    -9,    -9,   -18,    -8,    -9,     0,    -1,    -1,    -7,    -1,     0,    -1,    -4,   -11,    -5,    -8,    -1,     8,     5,     2,   -11,     1,     5,     7,    -2,     9,   -15,   -15,    -3,    -3,   -15,   -16,   -12,     3,    -2,    -8,    -4,     2,     2,    -2,     3,     4,     5,     2,   -12,     3,     6,   -13,    -2,     6,     8,    -6,    -3,   -11,   -18,    -9,    -5,    -6,   -10,    -7,    -4,     0,     1,    -3,    -1,     1,     0,     1,     1,    -9,    -3,    -7,    -1,    11,    11,     7,     1,     1,     8,     8,    10,     0,    -1,     1,     1,     2,     1,     0,     1,     0,     1,    -2,     2,    -2,     0,     0,    -1,     2,     3,     0,     1,    -1,     4,    -1,    -5,    -1,     3,     3,     2,     0,     0,     0,     3,     2,    -1,     0,     1,     4,     2,     2,     0,    -1),
		    78 => (   -2,    -2,     0,     2,     1,     2,    -1,    -1,     1,     0,    -1,     2,     1,    -1,     2,     1,    -1,     2,     1,     1,    -2,     0,     2,    -2,    -2,     1,     1,     2,     1,     2,    -2,    -1,    -2,    -2,     0,     0,     2,     1,     0,    -2,     1,     1,    -1,    -7,   -12,    -9,    -1,     1,     0,     0,     1,     2,    -1,    -2,    -2,     0,     2,    -2,     0,     2,     2,     0,    -1,     1,    -4,    -6,   -14,   -10,    -3,    -2,    -3,     0,     0,    -4,    -5,    -3,    -3,    -6,    -9,    -4,    -5,    -4,    -1,     1,     0,     0,    -4,    -1,    -1,    -8,    -5,   -12,     7,     4,    -3,    -4,    -1,    -4,    -8,    -4,    -2,    -6,    -1,    -3,    -4,    -3,     1,     2,     0,    -3,    -7,     2,     0,     1,     1,     0,    -8,   -12,    -1,     0,    -3,   -12,   -11,   -15,    -4,    -4,    -1,   -10,    -4,     9,     9,    -5,    -4,    -6,    -8,    -6,    -1,    -5,     2,    -3,     2,    -2,    -1,    -1,    -7,   -10,     3,     2,    -7,   -13,   -10,    -8,    -9,    -2,    -4,     0,     1,     2,     6,     3,     1,     0,    -4,    -2,    -1,    -3,    -2,    -7,     0,     2,    -6,   -12,    -2,   -10,     0,     2,    -1,    -1,    -7,    -7,     2,     2,    -1,     5,    -2,    -1,     1,     0,     2,     0,     2,    -1,     0,    -1,    -2,     1,     1,   -10,    -5,    -1,    -6,    -4,     3,     0,     2,     2,     5,     0,     1,    -7,    -1,     9,     2,    -2,     7,    -6,    -2,    -1,    -3,    -5,    -4,    -4,    -3,    -2,    -4,    -5,    -5,     0,    -6,    -4,     5,     0,    -1,    -1,     2,    -1,    -4,    -4,    -1,     9,     5,   -10,     2,    -3,    -9,    -4,    -2,     1,    -1,     3,    -1,     1,     0,    -4,   -10,     0,    -2,   -13,     3,    -3,     3,    -1,    -1,    -9,    -6,    -3,    -2,     7,     3,    -9,     3,     0,    -2,     0,    -1,    -4,    -8,    -1,    -5,   -12,     1,    -3,    -9,     2,    -2,   -11,   -11,     1,    -1,    -8,     2,     0,    -3,    -8,   -11,     3,    -6,     3,     1,     0,    -2,    -6,    -6,   -10,    -7,    -3,     7,    -9,     1,     1,    -5,     0,    -6,   -11,   -10,     3,    -3,    -9,    -3,    -6,    -9,   -12,    -4,     6,    -1,     0,     5,     3,    -3,   -11,    -7,     5,     0,     0,    10,   -10,    -2,     1,    -6,    -6,    -8,    -6,    -7,     0,     0,    -6,    -6,    -6,    -5,   -10,   -10,     6,     5,     2,     5,     2,    -1,     2,     4,    -6,    -4,    -5,    -4,   -15,    -1,     0,    -9,    -6,   -10,    -9,    -7,    -2,    -4,     1,   -13,    -9,   -13,   -14,    -6,    -1,    -3,     1,     8,     3,     1,     3,    -4,    -5,    -7,    -8,    -8,     0,     1,    -1,     1,    -5,    -1,    -5,   -12,    -5,    -3,     0,    -1,    -4,    -2,   -18,    -5,    -6,   -12,    -7,    -4,     1,     0,    -3,    -8,    -8,    -7,    -2,   -23,    -3,     0,     2,     0,    -4,     0,    -1,    -6,    -7,    -5,     2,    -1,    -7,    -1,   -13,    -1,     1,    -5,    -1,    -3,    -5,    -4,    -3,    -5,    -6,    -3,    -2,   -20,    -8,     0,    -1,    -1,    -3,     1,    -3,    -4,    -1,    -3,    -6,    -4,    -4,    -7,    -3,     4,     0,    -4,     1,    -4,    -5,    -5,    -3,    -6,    -4,    -3,     0,   -11,    -8,     2,     0,    -1,    -3,    -1,    -4,    -5,    -3,    -5,   -11,   -11,    -8,   -13,     2,     6,     4,    -3,    -8,    -2,    -1,    -1,    -3,    -5,    -3,     0,    -2,     0,    -8,     0,     1,     0,    -5,     0,    -4,    -3,     0,    -6,    -9,    -2,   -10,    -1,     5,     2,    -1,     2,    -8,     0,    -2,    -4,    -8,    -1,    -3,     2,    -1,     0,    -4,     1,    -2,    -7,    -7,     1,    -3,    -2,    -7,   -11,     0,    -3,    -5,     4,     4,     0,     6,     7,    -3,    -1,    -4,    -6,    -3,    -3,    -1,    -1,     0,   -12,   -10,     0,     1,    -2,    -1,     1,    -7,    -5,    -4,    -5,     4,    -1,    -4,    -2,    -4,    -8,     0,    -2,     5,     1,    -3,   -11,    -7,    -6,    -3,     1,    -2,    -9,     2,    -9,    -4,    -3,     0,    -5,    -9,    -7,   -12,    -1,     8,     0,    -9,     2,    -4,    -8,   -11,     0,    10,     2,     2,    -6,    -2,    -5,    -4,    -4,     0,   -11,     0,    -4,    -4,    -1,    -4,    -1,    -8,    -3,    -5,    -3,     5,     4,     2,     2,    -4,    -8,    -8,     6,     6,     0,    -1,    -3,    -9,    -8,    -4,    -4,    -2,    -7,     1,     0,     1,    -3,    -1,    -4,    -7,    -6,    -4,    -7,     0,     5,     5,    13,     4,     1,     0,    12,     0,    -3,   -12,    -5,    -4,    -6,    -2,    -3,    -1,   -13,     1,     1,    -2,    -2,    -3,     0,    -3,    -8,    -5,    -7,    -4,    -5,    -6,     1,    -1,     2,     2,     6,   -12,   -12,   -10,    -9,    -4,    -1,    -3,    -8,    -2,    -2,     1,    -1,     2,    -7,    -5,    -2,     0,    -4,    -8,    -7,    -7,    -7,   -17,    -2,     3,     1,     7,   -12,   -17,   -12,    -7,    -1,    -3,     0,     1,     0,    -5,    -4,     1,     0,     1,     2,    -2,     2,    -6,    -5,    -4,     0,    -6,   -10,   -12,   -10,   -13,   -18,    -9,    -4,     0,    -1,    -4,   -14,    -8,    -7,    -2,     0,     2,     0,     1,     2,    -2,    -1,    -1,    -2,    -1,    -4,     0,    -3,    -2,    -3,     0,     2,    -6,    -1,    -1,    -7,    -8,     0,     1,    -3,    -2,    -1,    -2,     0,    -1,     2,     2),
		    79 => (    0,     0,     2,     0,    -1,     2,    -2,     1,     1,    -2,    -1,     1,     2,     1,     1,     1,     1,    -2,     0,     0,     1,     0,     1,    -1,     0,     2,     1,    -1,     1,     1,     0,     0,     2,     1,     2,     2,     2,     2,     0,    -4,    -4,    -4,     1,     1,     1,    -1,    -1,     1,    -2,     0,     1,     2,    -2,     0,     2,    -2,     0,    -1,     1,    -1,     2,     0,    -2,     0,    -1,    -3,    -2,    -3,    -1,    -2,    -5,    -2,    -2,    -2,    -2,    -2,     0,     1,     2,     2,     0,     0,     0,     1,     0,    -1,    -2,     1,     2,    -2,    -2,    -3,    -4,    -3,    -6,   -11,    -2,    -7,    -9,    -7,    -9,    -1,     4,     8,    -5,    -3,    -5,    -3,    -1,     0,     2,     0,     0,     2,     1,     1,     0,    -2,   -10,    -3,    -3,    -8,    -8,     9,     6,     7,     0,    -7,    -8,   -13,   -16,   -14,   -17,    -8,    -6,     2,     1,    -9,    -5,    -2,    -2,     1,     0,    -2,     0,     0,    -2,    -4,   -16,   -20,   -13,    13,     0,     2,    -4,     6,    18,    -6,    -2,    -3,     6,    -9,    -9,    -4,    -6,    -8,   -10,    -1,     0,    -7,    -3,     0,    -2,   -11,    -1,   -16,    -6,    -9,    -5,    -7,     5,     5,     9,     5,     3,     4,    -5,   -12,   -14,    -3,    -7,    -4,    -2,    -4,    -6,    -4,     2,    -2,    -4,     1,    -2,   -16,   -15,   -30,    11,   -18,     4,    11,     6,     5,     4,    -6,    -5,   -15,   -28,   -13,    -8,    -7,    -6,    -6,    -4,    -4,    -5,    -5,    -4,   -13,    -5,    -3,    -5,   -10,   -20,   -22,    14,    -4,    10,    12,    10,    -7,   -18,    -3,   -13,    -4,   -10,     6,    -3,    -8,    -4,    -8,    -9,    -6,   -16,     0,     0,    -9,    -5,    -2,   -12,   -12,   -28,    -5,    12,     0,     7,     1,   -14,   -13,   -10,     1,    -3,     5,   -11,     4,    -2,   -10,     2,    -6,    -4,   -11,    -7,    -3,     1,    -3,     1,     2,    -6,    -5,   -12,     8,    13,     9,    -6,     3,   -10,     5,    19,    12,     0,     9,    13,     7,    -9,   -20,    -9,   -13,    -5,    -8,    -1,    -8,    -2,    -5,     0,    -2,    -5,    -7,    -3,     0,     8,     2,     1,     1,    10,    13,    17,     6,    11,    14,     4,     0,    -8,    -9,   -13,   -11,    -2,   -10,     0,    -7,     2,    -1,    -4,     1,    -3,    -7,   -12,    -6,    -3,    -4,    -3,     3,     0,     9,     0,     1,     4,     5,     0,     2,    -5,    -6,    -1,   -19,   -18,    -7,   -10,    -3,     1,    -3,    -3,   -11,    -7,    -6,   -12,    -3,    -5,     3,   -11,    -4,    -2,     6,    -1,    12,    10,     0,   -20,    -8,   -10,   -13,    -3,    -7,    -9,    -6,    -9,     0,    -1,    -3,    -6,    -8,    -6,    -6,   -12,    -5,   -16,    -2,   -11,    -7,    -1,     6,    -7,    -3,     4,     2,    -8,   -14,    -9,    -2,     7,    -3,    -1,    -8,    -4,    -2,     2,     2,    -2,    -7,    -1,    -5,    -3,   -25,   -21,     1,     5,     9,     9,    -2,    -2,   -10,     5,     5,   -17,   -14,   -17,     2,     6,    -4,     2,    -5,    -4,    -6,    -1,    -2,    -5,    -3,    -1,    -5,    -5,   -13,   -29,   -25,   -15,     0,    -3,   -16,   -10,    -9,    -1,    -9,    -8,   -22,   -14,    -4,     4,    -1,     3,    -6,     1,    -3,     0,    -1,    -7,     1,     1,     5,     4,    -6,   -10,   -19,   -24,   -37,   -20,   -12,    -5,    -7,    -5,    -7,    -9,   -20,   -12,    -4,   -10,   -10,     6,    -2,    -4,    -3,     8,     2,    -6,    -4,    -4,    -9,    -6,    -7,   -10,   -11,   -16,   -31,   -13,    -7,    -5,   -12,    -5,    -3,   -11,   -17,   -24,   -10,   -11,   -16,    -8,    -1,    -2,    -5,     2,    -4,    -1,     0,    -3,   -13,   -16,    10,    -9,   -12,   -14,   -20,    -6,    -6,    -3,    -6,    -8,   -13,    -6,     0,   -18,     3,    -1,    -3,    -5,    -4,    -5,     3,     0,    -4,    -3,    -2,    -3,     3,   -11,     3,     4,    -5,     1,    -7,    -4,    -4,    -7,   -11,    -7,   -10,    -1,    -5,   -16,     0,     6,    -1,    10,     3,    -2,     1,     0,     2,    -6,    -4,     5,     8,   -15,     0,     8,    16,     4,    -2,    -3,    -3,   -14,   -10,   -13,    -2,    -1,     0,    -4,    -8,    -2,    10,     6,     7,    -8,     0,     1,    -2,   -14,    -8,     0,    -4,   -16,   -10,     8,    11,     1,     8,     1,    -1,    -2,    -7,    -1,    -3,     5,     2,    -1,    -6,    -5,     4,    13,   -11,    -2,    -2,     2,     2,    -1,    -6,    -1,    -9,    -9,   -13,     0,     8,     7,    12,     5,     5,     7,     5,    -1,    -3,     5,    -1,     4,   -11,     4,     3,    10,    -3,    -2,     1,    -1,     0,    -1,   -13,     0,     0,    -3,     0,     4,    -1,     5,    -2,    -9,    -6,     0,    -3,     3,     0,   -10,   -13,     7,     0,     1,     3,    -1,    -2,    -2,    -1,     0,    -1,     4,    -5,     0,     0,     7,    11,    -1,     3,    -7,    -9,    -9,   -10,    -4,     1,     2,    10,   -11,   -14,     8,     2,     7,     6,    -1,    -1,     1,    -1,     1,     2,    -1,     6,     2,    -1,    -4,     2,   -19,    -1,    10,     4,    -2,    -1,    15,    -5,   -15,   -12,    -7,    -9,    -2,     1,    -3,     4,     4,    -1,    -2,    -1,     0,     2,     2,    -2,    -4,    -3,     2,     2,    -4,    -6,    -2,     7,     1,    -4,     0,     7,    13,    -8,     1,     0,     1,    -3,    -2,     1,    -2,     2,     1,    -1),
		    80 => (    0,     2,    -2,     2,    -1,     1,     1,    -2,    -2,    -2,     0,     1,    -2,     2,     1,     2,    -2,    -2,     2,     2,     0,     2,    -1,     0,    -1,    -2,    -2,     1,    -1,     2,     2,    -1,     3,     2,    -1,     2,    -1,    -2,    -2,     2,     1,     3,    -4,    -2,     1,     1,    -3,    -1,     0,     1,     0,     0,     0,    -1,    -2,     0,    -2,     0,    -2,    15,    14,     0,     2,     3,    -2,    -4,    -1,   -11,    -9,   -15,   -17,   -15,    -9,   -11,    -9,   -11,    -8,    -9,   -10,    -6,    -9,    -4,    -1,    -1,    -2,    -1,     2,    18,    11,     6,    -3,    -4,    -8,    -7,    -7,    -4,    -6,     7,     2,    -5,     2,    -3,    -4,    -1,     2,   -17,   -12,   -10,     0,    -3,    -8,    -2,     0,     1,    -2,    -1,    -4,    -5,    -8,    -8,    -8,    -5,    -5,    -7,   -11,    -5,    -3,     2,    -7,     1,     9,     3,     9,     5,    17,    -5,    -1,    -6,   -10,    -1,     0,     1,    -3,     3,     2,     1,     3,   -14,   -17,   -15,   -16,   -23,   -13,     0,    -2,    -3,    -5,     5,     5,     4,    12,     7,    18,    -3,    -1,    -7,    -9,    -4,    -2,     1,    -4,    -3,     3,    12,     2,     2,   -13,   -23,   -19,   -20,    -3,    10,     0,     3,   -14,    -5,     0,     2,    -2,    14,    10,    -9,   -17,   -20,   -11,     0,    -2,    -1,    -2,    -4,     7,    14,     3,    -5,    -8,    -5,    -7,     3,     0,     1,    -9,    -2,    -4,    -3,    -1,     7,     4,    -8,     6,     5,    -3,    -4,   -15,     4,     6,    -5,     6,    -5,     1,     9,     6,    -6,    -7,   -11,   -16,   -15,    -6,    -5,     9,    -7,     4,    -2,     4,     3,     2,     9,     8,     5,   -10,   -14,   -15,    -3,    -1,    -1,     7,    -2,    -6,     8,    -5,    -8,    -4,   -20,    -6,   -13,    -5,    -3,     9,     5,    -9,    -2,     4,     0,     5,    -2,     4,    10,     9,     3,   -11,     1,     1,    -1,     4,    -1,   -10,    -4,   -16,    -6,    -8,     3,    -7,    -3,     8,    -1,     2,     6,     1,    -9,   -15,    -6,    13,     8,    11,    10,     9,     4,   -18,    -2,    -2,     7,    -6,    -5,   -12,   -12,    -9,     8,     2,    -2,    -5,     2,     2,    -6,    -3,    -8,   -19,   -23,   -22,     0,     4,     5,     0,    -1,    -3,    -1,   -10,    -1,     2,     6,    -2,    -3,    -5,    -9,    -8,    -1,    -2,    -3,     7,     8,     7,     8,     4,    -4,   -33,   -30,    -7,     6,   -10,    -3,     4,    16,    -2,    -4,    -9,     0,     2,     5,     4,    -8,    -6,    -5,     0,     3,     3,     6,     1,     7,     5,     6,     1,    -9,   -40,   -15,     8,    -1,    -9,   -11,     1,    31,     9,     7,    -8,    -2,     0,    -1,     0,   -21,    -5,    -3,     4,    10,     0,     3,    -9,     0,    -3,    -4,   -33,   -28,   -30,   -13,    -7,    -6,    -6,     3,     2,    14,     4,    -4,   -15,     0,     0,     1,    -5,   -23,     3,    -7,     1,    12,     4,     4,   -13,    -5,     7,    -1,   -23,   -16,    -5,    -1,    -8,    -5,   -16,     2,     3,     9,    15,   -10,   -16,    -4,     2,     2,     0,   -16,     4,    -1,    -1,    11,     7,    -6,    -6,     1,   -10,   -16,    -6,    -2,     1,    -4,     3,    -9,    -4,    -9,    -4,     1,     8,   -13,    -7,     1,     0,    -3,    -7,    -8,     3,    10,     4,    11,    -5,     3,     0,    -7,   -22,   -15,    -9,    -2,    -7,     0,    -1,     4,     4,   -11,    -8,     3,     7,   -14,    -8,     1,    -2,     1,    -5,    -1,     5,     1,     3,    10,    14,     6,   -11,   -22,   -17,    -7,     1,     2,    -2,     0,     4,    -8,    -1,    -3,     4,     2,     2,    -7,    -4,    -3,     2,     3,   -13,    -4,    16,    -1,     1,     7,     3,     7,   -10,   -20,    -8,   -11,     0,     3,    -8,     2,    -6,    -4,   -12,    -3,     4,     0,     6,    -9,    -2,     2,     1,     4,   -19,     5,    13,     3,     7,    -2,     5,     4,    -2,     4,    -4,    -5,    -3,   -14,    -3,    -4,    -3,   -13,   -15,    -5,     2,    -2,     2,    -8,     2,     3,     1,     2,   -18,     5,     3,     2,     7,    11,     3,     5,     0,     0,    -7,    -4,     1,     6,     0,    -2,   -10,   -13,   -18,   -18,   -11,    -3,     9,    -5,     2,     3,     1,    -2,   -21,     0,     0,     9,    12,     5,     4,     3,     5,    -6,    -7,     2,     8,     1,   -18,   -14,    -6,    -7,   -21,   -12,    -2,    -2,     8,     1,     0,     3,     2,     0,    -3,   -15,   -17,     2,     2,     0,     2,     7,     8,     7,     1,     6,     6,   -11,   -17,   -11,   -15,   -14,   -20,    -9,     3,     0,   -12,     0,    -1,    -2,     0,    -1,    -4,    -3,    14,    19,    -1,    -4,     1,    10,    17,    11,    15,   -16,   -14,   -14,   -29,   -24,   -14,   -15,    -7,     2,    -2,    -1,     6,     2,    -1,    -2,     2,    -2,     0,     0,   -10,   -19,   -17,   -18,   -15,   -10,   -13,   -15,   -20,   -15,    -6,   -17,   -18,   -16,   -19,   -14,    -1,    -4,    -3,    -3,    -1,     0,    -2,     1,     2,     1,    -1,    -2,    -2,   -14,   -19,    -5,     0,    -5,    -8,    -9,    -5,    -7,    -6,   -10,   -11,   -18,   -19,    -4,   -12,    -5,    -5,    -3,     0,     1,    -2,     1,    -2,    -2,     2,     2,     0,     1,     2,    -2,    -1,     0,     1,     2,     2,    -1,     0,     0,    -1,     1,     0,    -3,    -2,    -3,    -3,    -2,     0,     0,     2,    -2),
		    81 => (   -2,     1,     2,     2,    -1,    -1,     0,    -2,    -2,     1,    -1,     2,     0,    -1,     2,    -1,     1,     0,     1,     0,     2,    -1,     2,     0,    -2,     2,    -2,     2,    -1,     1,     2,     0,     0,    -2,     0,    -1,     1,     2,     0,    -1,     0,    -4,     3,     3,    -1,    -3,     0,    -2,    -1,     0,    -1,     1,     1,    -1,     1,    -1,    -2,     1,    -2,     2,    -1,     2,     0,    -2,    -3,    -3,    -3,    -2,     0,     0,    13,    16,    33,    24,    12,    -8,     2,   -11,    -8,    -6,    -1,     2,     2,    -1,    -1,     0,     6,     5,    -3,    -8,   -17,    -6,    11,     4,    -7,   -13,   -11,    -3,     5,    18,    20,     4,     1,    -9,     1,    11,    -3,     0,    -8,     0,     1,    -1,     2,     2,     6,     6,    12,     5,    -4,    -5,    17,    13,     8,    -2,    -1,    -7,    -2,     5,     6,     3,    -4,    -4,     9,    11,     5,     8,    -1,    -6,    -6,    -8,     0,    -2,    -1,    -2,    14,    26,    11,    10,     7,     3,     2,   -13,   -13,     3,     8,     2,    -4,     2,     1,     5,     9,     9,     8,     3,     1,    -3,    -7,    -7,     2,     1,   -17,     1,     2,     6,    11,     4,    -8,   -10,     5,    -3,     0,    -2,    -1,    -3,   -10,     7,     4,    12,     7,    -2,     3,    -1,    -1,    -2,    -4,    -2,    -2,     2,   -19,   -16,   -16,    -1,     6,     8,   -13,     2,     9,    -7,    -2,   -11,    -2,     7,    -2,     3,     7,    13,     2,    -1,     4,    -4,    -4,     0,    -8,    -4,    -1,    -2,   -21,   -13,   -15,    -3,     3,     1,    -3,     6,     3,     2,     6,   -10,   -11,     2,     8,     1,     8,   -11,    -6,    -5,     3,    -7,    -1,    -1,    -8,    -1,     1,    -1,   -21,    -8,   -10,   -11,     0,     6,     9,     1,     2,    15,    12,    -7,   -14,    -4,    -7,    -7,    -8,    -6,    -5,    -6,    -8,     0,    -3,     2,     1,    -3,     0,    -1,   -16,    -3,   -18,    -9,   -16,     2,     7,    10,     4,    17,     4,    -4,    -7,    -4,   -10,    -8,    -3,   -15,    -9,   -11,    -1,    -1,    -3,    -2,     3,     0,     0,     3,    -4,    -2,   -15,    -8,   -14,     0,    -7,     5,     1,     9,     4,    -3,    -2,   -10,     1,   -11,   -10,   -13,    -8,    -7,     2,     0,    -2,    -2,    -1,     3,    -1,    -1,    -2,    -6,   -10,   -11,     5,     9,     2,     1,    -5,     1,    -1,    -8,   -11,    -3,    -3,   -12,    -4,   -14,   -20,    -9,    -5,    -5,    -2,    -3,     1,     4,     0,    -1,    -3,    -2,   -14,     6,     9,     9,    13,    -5,    -7,    -1,    -3,   -11,    -5,     7,    -3,    -8,    -9,   -29,   -13,   -11,    -9,    -8,    -7,    -1,    -1,    -1,    -1,     0,     2,    -1,   -12,    11,     9,    -2,    -4,   -17,   -22,   -12,    -8,    -7,     3,     4,    -1,    -7,   -12,   -19,   -17,   -20,   -13,    -8,    -5,    -8,     1,     2,    -2,     1,    -1,     4,    -2,   -10,    -6,    -6,   -11,   -14,   -18,   -19,   -22,    -2,     9,     2,    -3,    -8,   -11,   -25,   -14,   -15,   -12,   -13,   -29,    -4,    -1,    -3,     1,    -1,     3,    -6,    -5,    -6,    -9,    -9,   -19,   -10,   -12,   -20,   -18,    -2,    13,     9,    -3,   -11,    -9,   -20,   -17,   -21,    -7,   -14,   -10,    -4,    -3,    -4,    -1,    -1,    -1,   -11,    -3,    -5,    -8,   -15,   -15,   -14,   -16,   -35,   -19,   -16,     6,    -6,    -5,    -6,     1,    -7,   -10,    -7,     0,    -8,   -15,   -16,    -1,    -6,    -3,     1,     2,    -3,    -3,   -12,   -24,   -14,   -24,   -16,   -17,   -44,   -38,   -21,     0,    -8,    -3,     3,    -4,    -3,     9,     6,    13,    -6,   -29,    -6,    -6,    -5,    -1,     0,    -3,    -5,    -8,   -22,   -13,    -3,    -1,    -9,   -12,   -21,   -14,   -11,    -7,     5,    10,     1,    -9,    -1,     4,     0,    -1,     6,    -2,    -1,   -10,    -3,     1,    -2,    -6,     8,    -1,   -17,    -7,     3,     3,     7,    14,     2,    -4,     1,     5,     5,    14,     8,    20,    15,    12,    -1,     5,     6,     3,     2,    -7,     2,     5,     2,    -8,     9,    11,     4,    11,    10,    12,    12,     7,     7,    -1,     5,     5,    11,     3,    12,    19,     6,     7,    -1,    -9,    -5,     4,     8,    -9,     2,     5,     1,   -24,   -14,     7,    17,     6,     1,     3,     5,     5,     4,     3,     4,    -2,     4,    -4,     4,     2,    10,    11,     6,   -18,   -12,     3,    -2,    -1,     0,     2,     1,    -2,    -7,     4,    -4,     6,    -3,    -1,    -5,    -7,     1,     1,     7,    -9,   -14,   -19,   -15,    -5,     3,     9,    10,    -4,   -10,   -10,   -13,     6,     1,     0,     0,    -2,     0,    -4,    -7,   -10,    -2,     3,     6,    -3,    -2,   -18,   -12,   -23,   -19,   -17,   -10,    -7,    -2,     2,     4,    -6,    -8,   -11,    -2,     0,     2,     0,    -1,     2,    -3,    -1,    -1,    -5,    -2,    -1,   -11,    -5,    -7,   -10,   -12,    -8,   -15,   -11,   -13,   -15,   -13,   -16,   -13,   -10,    -4,     0,     1,     1,    -2,    -2,     2,    -1,     1,    -4,    -4,    -5,    -4,    -3,   -11,     0,    -2,    -5,    -8,    -6,   -10,    -3,   -11,    -6,    -9,    -7,    -5,    -4,     1,    -2,    -1,     2,    -1,     1,    -1,    -1,    -2,     0,     2,     1,    -1,     0,    -1,    -4,    -4,     0,    -3,    -2,    -3,    -3,    -2,    -2,     0,     0,     0,    -1,     0,     1,     1,    -1,     2),
		    82 => (    1,     1,    -2,    -2,     0,    -1,     1,    -2,     2,     0,     0,     1,    -2,     0,     3,     2,    -1,     0,    -2,     1,    -1,    -2,     2,    -1,    -2,     1,     0,     0,     0,     2,     2,    -1,    -2,     2,     1,    -6,    -9,    -4,    -9,    -8,    -9,   -17,    -7,     1,     8,     1,   -10,   -19,   -12,    -7,    -9,    -3,    -1,    -1,    -1,     1,     1,     2,     0,   -13,   -14,     2,    -1,    -2,     0,    15,    13,     6,     3,     4,     2,     6,     0,    -1,    -7,   -12,    -7,    -6,    -4,     0,     2,     3,     0,     0,     0,    -1,    -1,   -15,   -19,    -2,    -1,     5,    -5,     6,     3,     2,    -4,     5,    11,     6,     6,     1,    -6,    -8,    -5,     2,   -10,   -24,     2,     3,     1,     0,     0,     1,    -4,     4,     4,    -6,     2,    -2,   -13,     6,    12,     2,     2,     7,     9,     3,     6,     3,    13,     2,    -1,    -4,   -11,    -5,    -8,    -3,    -5,     0,     0,    -2,     4,    -1,    -1,     3,     4,   -12,    -1,     3,    -8,    -6,     3,     0,     0,    -2,     9,    -4,     2,    -6,    -4,    -4,    -7,    -4,   -16,    -1,    -6,    -5,    -1,     1,     1,    -6,    -6,     1,     1,     9,    -8,    -7,     3,    -5,   -11,    10,    -1,     3,    12,     2,     3,   -10,    -5,    -1,    -6,    -9,   -20,     8,    -4,    -3,    -2,     1,    -2,    -5,    -6,    -3,     6,     0,    -8,    -7,     7,     2,     0,    -8,     1,     5,    -1,     2,   -13,    -3,     6,     9,    -2,   -20,    -7,     2,   -10,    -4,    -4,     4,    -4,    -8,    -5,   -12,    -7,     1,     5,     4,    10,     6,   -11,    -7,   -14,    -1,     0,     3,     4,    10,     1,     2,     1,    -9,   -16,   -20,    -7,    -3,     0,    -4,    -2,    -7,    -4,   -17,   -14,   -18,   -22,    -6,     1,   -11,   -17,    -1,    -2,   -10,    -3,     4,     7,    -7,    -3,    11,     0,    -9,    -9,   -11,    -7,    -6,    -2,     1,    -2,   -11,   -12,   -16,   -18,   -35,   -49,   -44,   -36,   -29,    -9,   -11,    -2,   -12,     1,    -5,     5,     1,    -1,    -4,    -1,    -4,   -15,   -12,    -6,    -2,    -1,    -7,    -7,   -13,   -13,   -16,   -25,   -30,   -39,   -34,   -28,   -16,   -12,   -16,    -4,   -11,    -8,   -18,   -17,     1,     0,     1,     6,    -5,   -15,    -2,    -6,    -4,     2,    -8,   -17,   -12,   -21,   -15,   -14,   -18,    -5,    -4,    -3,     3,    -2,    -3,     2,    -7,   -13,   -15,   -11,    -6,    -3,     5,    11,   -12,   -12,    14,     2,    -3,    -2,    -7,     1,    -4,   -10,    -7,     2,    19,     8,    -2,    -5,     4,    18,    12,     5,     3,     0,     0,    -7,    -8,    -1,     7,    14,    -1,    -3,     6,    -1,     0,     0,    -7,   -10,    13,     8,    -2,    13,    19,    16,    11,    16,    12,    10,    16,    14,    -2,     8,   -13,    -7,    -3,     6,    -1,     3,     3,    -3,     9,     8,     7,     0,    -5,     2,    29,    13,    16,     9,     9,     8,     8,    14,     5,     7,     4,    -7,     5,    -2,     2,    -6,     0,    -7,    -5,    -3,     8,    -2,    12,    22,    14,     0,     1,     3,    12,    -4,    15,    23,    11,     5,     7,     9,     1,    -8,     5,     5,     4,     3,     4,    -1,     1,    -7,    -9,    -5,    -3,   -10,    17,    22,     9,     2,    -4,     1,    -6,     7,     5,    15,    -4,     7,    -6,    -8,     4,     0,    -3,    11,     7,     7,     1,    -1,    -7,    -2,   -17,   -12,   -14,   -18,     2,     5,    15,     1,    -2,    -9,     3,    -1,    11,    12,     0,     0,    -5,    -8,    -4,     0,     3,    -3,    -1,     8,     2,     7,    10,     5,    -5,    -8,    -7,     3,    11,     6,    14,     1,    -8,    -8,    -4,     7,     7,     8,     7,     4,     2,    -7,     2,     1,    -3,    -7,    -2,     2,     0,     9,    10,     2,     8,     9,     4,    13,    12,    10,     7,    -2,   -10,     1,    -1,     5,    16,     5,     1,    -2,    -9,    -5,   -10,   -13,   -12,   -12,    -2,     0,    -9,    -7,    -2,    -3,     0,    -4,     3,    15,    -2,     4,    -1,    -3,     6,     0,     4,     7,     5,     4,     4,     6,    -8,    -9,    -2,    -3,   -12,    -8,    -8,    -9,    -3,    -8,    -1,     6,    10,     4,     9,     5,    -8,    -5,    -1,    -2,    -2,    -1,     3,     7,    -8,    -7,    -3,    -2,    -7,    -2,     2,    -4,   -11,   -14,    -5,    -9,   -10,   -14,    -2,     1,     2,    -3,    -5,    -6,   -14,   -16,    -2,    -2,    -2,     4,    13,    12,     2,   -13,    -3,    -8,   -15,    -4,    -9,    -1,   -18,   -10,   -17,    -6,    -9,   -11,   -19,    -9,     0,     8,   -12,   -11,    -8,   -11,     2,     1,     2,    -7,    -5,    -5,    -2,    -4,   -10,   -12,   -20,   -23,   -17,   -14,   -22,   -17,   -14,   -14,    -6,    -9,   -19,   -24,   -14,   -22,   -13,     4,     6,     7,     1,     0,     1,    -3,     0,    -5,    -4,    -3,    -7,   -13,   -18,    -6,    -4,    -6,   -16,   -13,    -8,   -12,   -15,    -9,   -20,   -15,    -9,   -12,    -4,    -5,     4,     9,     0,     1,     2,    -1,     1,    -4,    -7,    -6,    -4,    -5,    -2,    -2,    -1,     0,    -1,    -7,    -3,   -16,   -12,   -10,    -7,    -4,    -3,    -2,    -5,     2,     0,    -1,     0,     2,     2,     0,    -1,    -2,     0,     0,    -2,     1,     2,    -5,    -2,    -2,    -4,    -1,    -1,    -1,     0,    -3,    -3,    -6,    -7,    -5,    -2,     0,     0,    -1,    -2),
		    83 => (    2,     0,     1,     1,    -1,    -1,    -2,    -2,    -2,     0,    -1,    -2,    -1,     0,    -4,    -3,    -1,    -1,     1,     0,     2,     0,     2,     2,     1,    -2,     2,     2,     0,     1,     0,    -1,     1,    -2,     1,    -2,    -2,    -1,    -4,    -3,    -4,   -11,    -8,    -8,    -4,   -12,    -6,    -6,    -4,    -3,    -3,    -1,     2,     1,    -2,    -2,    -1,     1,    -1,     0,    -5,    -5,    -6,    -6,   -12,   -16,     6,    -1,    -5,   -10,   -13,   -13,    -9,    -1,     2,   -11,   -15,   -20,   -18,   -15,    -3,     2,    -2,     1,    -1,     2,    -3,    -3,    -3,     6,    11,    28,    27,    10,    12,    11,     9,     4,    -2,    14,    18,    12,    10,    23,    41,     4,   -26,   -27,   -14,    -7,     1,     1,     2,    -1,   -16,     1,     6,     8,     3,    17,    22,     0,    12,     6,     7,    -2,     5,     0,     8,    12,    10,    10,     4,   -14,   -14,   -53,   -41,   -15,   -11,     1,     1,     2,    -2,    -1,    -2,     9,    20,    24,     3,     6,     9,    -4,    -8,     1,    -5,    -1,    11,    -6,    -2,     7,     2,    -3,    -4,     3,     4,   -20,    -9,     1,     1,     3,     5,    -1,    -3,    17,    26,    22,    11,    11,     5,     1,    -7,     4,    -1,     7,     6,     2,     3,    -2,     1,    -3,    -1,     2,     8,   -23,   -11,    -4,    -1,     1,     1,     5,    -2,     4,    25,    32,    16,     1,     2,    15,     2,    -9,     3,    -1,     6,    -4,    -8,     4,    -4,    -4,    -7,    -3,     7,   -21,   -13,    -6,    -7,    -3,   -10,    -1,     4,    18,     3,     8,     2,    -4,    -3,   -12,   -14,    -8,    -4,    13,     6,     8,   -10,     7,     2,    -9,     6,     1,    -6,   -14,   -13,    -1,     0,    -5,   -24,    -5,    26,    25,    11,    11,    13,    -6,     5,    -8,    -7,    -4,    -6,    -6,     1,    14,     7,    -2,     5,    -5,    15,    12,   -28,   -12,    -9,     1,    -2,    -1,   -27,     2,     5,    13,    15,    19,     0,    -5,   -13,   -15,    -8,   -13,    -4,    -7,    -1,     8,    10,     4,   -11,    -9,     5,    18,   -13,   -13,   -11,     0,    -2,   -10,   -12,    14,    22,    20,    13,     5,     9,    -5,    -2,   -12,   -12,    -4,    -1,   -11,     2,     2,     6,   -10,   -13,    -7,     1,    -5,   -34,   -24,   -11,    -2,    -2,    -3,   -13,     5,    14,    21,    14,     8,     2,    -9,     4,    -5,    -7,    -7,    -8,     2,     2,    -1,     2,     5,    -7,   -15,    -6,     1,   -21,   -15,    -5,    -2,     2,    -3,   -11,     1,    22,    15,    10,     7,    17,    -1,     7,    -5,    -7,    -3,    -5,     9,   -23,    -6,    11,     9,    -8,    -9,   -11,     7,    -4,   -24,    -6,    -2,    -1,     6,    -2,     5,    10,    16,    16,    -2,     7,     0,    -5,    -3,     0,    -6,     4,   -11,   -11,    -3,     6,     7,     5,     3,    -4,     6,    -4,   -33,   -14,     2,    -3,     7,    -6,     3,     7,    20,    12,   -11,    -6,   -13,    -1,    -9,    -4,    -9,    -7,    -4,   -11,   -12,    -4,    13,     1,     4,     7,    15,    16,   -33,     6,    -7,     2,     1,     3,    21,    20,    17,     3,     7,   -15,     1,     1,   -12,   -20,    -3,     2,    -5,   -12,    -9,    10,    16,     3,    -6,     7,     2,    11,   -37,   -16,    -9,     0,     4,    -4,    10,    13,     3,    -5,     2,    -6,    -4,    -9,    -9,     0,     0,   -12,    -8,     3,     4,     8,    15,    -2,     1,    -8,    -6,    -8,   -30,    -9,    -4,    -5,     3,    -2,     7,    17,    12,     0,    -1,    -5,   -12,     0,    -4,   -10,     9,     0,     9,    -1,     6,    15,    -8,     5,    -6,    -4,   -19,    -5,   -30,    -2,    -8,    -2,    -5,     5,     3,     7,    11,    -6,    -8,   -10,   -18,    -9,   -11,    -2,     3,    11,    10,     1,     9,     8,    -4,     5,    -2,    -5,    -7,     5,   -15,   -12,    -9,    -1,     4,   -12,     3,     6,     8,     0,    -3,   -11,     0,    -9,    -8,    -4,     0,    10,     7,    19,    13,    -3,    -3,     8,     7,     8,     9,    -1,   -21,    -9,    -1,    -3,    -3,     5,    -1,     2,   -11,     8,    14,     0,    -4,    -7,     0,     4,     9,    14,    15,    11,     5,     7,    14,    -1,     7,    12,    -3,   -17,   -21,   -11,    -2,    -2,     0,    11,     8,   -11,     6,    14,    16,    -3,     3,     8,     4,    -5,     3,     9,     5,    -7,     6,    -4,    11,     2,    10,    21,     4,   -13,   -14,    -9,    -2,     2,     2,     5,     1,    -6,    -3,     6,    14,     5,     4,     3,     7,    -1,    -5,    -4,     7,     5,    -1,    -5,    -9,     1,    22,    21,    10,    18,     7,   -11,     2,     1,     0,    12,    20,    18,     0,    14,    13,     9,    16,     5,    -5,    -4,     2,     5,    -5,    -1,     2,    -9,     5,    28,    18,    10,    12,   -18,   -11,    -3,    -1,     2,     0,     3,    -6,     0,    17,    13,    -2,     5,     6,    -8,    -3,     6,    17,     1,    -2,    -2,     3,     8,     9,    -8,   -22,   -25,   -24,   -19,    -6,    -4,    -2,     0,     2,     0,    -3,   -24,    11,     6,     2,     7,    -6,    -5,   -11,   -11,    -6,    -9,     1,    22,    23,    21,     4,    -5,    -9,   -26,   -13,    -1,    -1,     1,     2,     0,    -2,     2,     1,    -4,    -7,    -7,    -3,    -5,   -15,   -13,   -11,    -9,   -15,   -13,    -8,    -1,    -3,    -1,   -11,   -14,    -4,    -5,    -3,     2,     1,     2,     1),
		    84 => (    0,    -1,     2,     1,     1,     0,     1,     1,     2,     0,     0,     0,    -8,    -4,    -3,    -4,     0,     1,     1,    -2,     2,     0,     1,     0,    -1,     1,     0,    -1,     1,    -2,     1,    -1,    -1,    -5,    -8,   -11,    -6,   -10,   -10,    -9,   -12,   -13,    -3,   -12,   -11,    -2,    -6,    -6,   -11,    -7,    -5,    -9,     0,     1,     2,    -2,     2,     1,    -5,    -9,   -12,   -15,   -14,   -14,   -23,   -20,   -28,   -30,     3,     6,    -1,   -15,   -14,   -18,   -26,   -14,   -29,   -13,   -14,    -9,    -5,    -7,     2,     1,     2,    -1,    -2,   -27,   -17,   -19,   -11,   -16,   -12,   -24,   -21,   -22,   -14,   -30,    -3,    -2,   -15,    -9,    -8,    -1,    11,     0,   -13,   -16,    -9,    -6,    -3,     0,     1,     2,   -12,   -26,    -2,     0,     5,     0,   -13,     1,    -4,   -18,    -2,    -4,    -8,   -11,    -5,    -1,    -3,     2,     0,    -8,     3,     4,     6,    -5,   -17,    -3,    -2,    -2,   -13,    -2,     1,    -4,    -1,    -3,     7,    -4,     9,     0,    11,    -9,    -5,   -12,    -8,     7,    -2,     2,   -11,    -5,     2,    -1,    -6,     6,    -7,    -1,    -1,     2,    -7,   -11,     5,    13,     8,   -12,    -4,   -13,    -1,     4,    -1,    -8,   -20,   -21,   -16,   -12,   -17,    -9,   -20,    -1,    -1,    -2,    -5,    -2,     0,    -9,     2,   -24,    -9,     0,     6,    10,   -10,   -13,   -18,    -8,    -4,    -1,   -14,   -11,   -14,   -18,   -16,    -5,    -9,   -11,   -10,    -8,    -8,    -6,     3,    12,    11,   -15,    -8,   -20,    14,     4,    11,     4,   -17,   -19,   -21,    -9,   -17,   -12,    -9,    -2,   -24,   -14,   -14,    -3,    -6,    -3,   -10,   -11,    -7,    -2,    10,    11,     0,    -5,     0,   -16,    12,     3,    -9,    -1,   -13,    -8,   -10,   -11,   -16,    -5,     0,    -6,   -14,    -6,    -9,    -4,     1,     6,     5,    11,     6,     8,    12,    -9,   -15,    -5,     3,   -10,     8,     2,    -7,     7,    -5,   -12,    -6,    -1,    -1,     1,     9,    -3,    -7,    10,     8,    16,    -4,     1,     7,     5,     4,    -1,    -2,     2,    -8,    -3,    -2,   -12,    -2,     0,     1,    14,     0,     1,     4,    16,    12,     7,    15,    -4,     1,    10,    16,     3,    -6,    -3,     0,     2,     7,     6,    -3,    -3,   -17,   -15,    -1,    -1,     7,     8,    -2,    11,     9,     6,    10,    12,    12,    11,    14,     6,    -4,    -1,     1,    -3,    -8,    -1,    -3,     6,    11,     6,    17,    10,     8,   -17,     2,    -3,    -1,    14,     6,    13,     5,     9,     1,     7,     7,    18,    16,     9,     0,    -5,     8,     5,   -10,     2,     3,    12,     8,    11,     9,    23,    21,   -10,     2,     3,   -22,     6,    21,    15,     7,     6,    13,     9,     7,     6,    11,     0,    -4,    -6,     9,    15,    -8,    13,    -6,    15,     7,    -6,    -1,    13,    13,    -2,    -1,     4,    22,    10,     0,    12,     4,    -5,     3,     6,     7,     6,     4,     3,    -3,     9,    14,     3,     0,    11,    -1,    -1,    14,     8,    -6,     9,    26,    -3,     0,     1,    -5,    14,     5,    11,    14,    10,     7,     3,    -1,    -4,     5,     0,    -3,    15,     5,     7,    15,    19,     6,     3,     0,     0,    -2,     8,    16,    -6,    -2,    -4,     6,    -5,    18,    13,     6,     8,     1,     2,     1,     0,     1,     5,     5,     5,     8,     2,     1,     9,    -7,     0,     3,     3,     3,     2,    10,    -1,   -14,     0,    13,     6,    14,     0,    -3,    -3,     4,     9,     1,     7,     2,    10,    11,     2,     2,     3,     6,    -5,    -4,     1,    -3,    -7,    -4,   -15,    -5,    -5,     1,   -10,    -7,    18,    -1,    14,     2,   -12,     6,     2,    -7,     2,     1,    -4,     9,     1,    -5,    -6,    -8,   -16,   -11,    -9,   -16,   -18,    -5,   -11,    -6,    -5,    -1,    -2,   -13,    12,     7,     0,     1,     1,     3,   -10,   -23,   -13,   -17,    -8,    -4,   -10,    -5,   -13,   -15,   -13,   -23,   -18,   -13,   -16,    -5,   -26,    -5,     0,    -1,    -4,   -20,     6,     8,     3,   -11,   -18,    -6,   -11,   -16,    -9,   -14,   -10,   -16,    -7,     0,    -6,   -10,   -16,    -6,   -13,    -7,   -11,     3,   -15,   -17,    -1,    -3,     0,     0,   -15,   -23,    -4,     0,   -18,   -20,   -18,    -3,    -5,   -12,   -14,    -8,    -4,    -9,   -11,    -9,    -4,   -12,     3,     2,     8,    -8,    -6,    -3,    -4,    -2,    -1,    -1,   -20,    -9,   -23,     0,     6,     1,   -14,     7,    -7,    -5,    -6,    -7,    -5,    -6,     1,    -7,    -3,    -7,     3,    -5,   -12,   -17,     1,    -1,     2,    -1,     1,     0,    -3,   -18,    -1,     5,     8,     7,     5,    -9,    -3,   -16,     6,     8,    -8,    -1,    -9,   -20,   -13,    -2,     6,    -3,   -10,   -28,    -4,    -7,     1,     0,    -2,    -6,    -3,     4,   -14,     3,     0,    -6,   -13,    -5,    -5,   -17,   -14,    -7,   -21,    -3,    -7,   -10,   -16,    -4,    -1,     7,    -2,   -18,    -8,    -6,    -1,     1,     2,     0,   -15,    -7,    -4,   -15,   -17,    -7,    -8,   -25,   -18,   -13,   -26,   -23,   -17,   -23,    -9,    -5,   -25,   -34,   -33,   -29,    -8,    -7,    -2,    -2,    -1,     2,     0,     2,    -2,    -1,    -3,    -3,    -3,    -5,    -6,   -20,   -22,   -12,   -16,   -21,    -7,   -11,   -22,   -14,   -16,   -19,   -14,   -13,    -4,     2,    -1,     1,    -2),
		    85 => (    1,     0,     2,    -2,     0,     0,     1,    -3,    -1,    -2,    -2,    -2,    -2,    -3,     0,     1,     1,    -2,     1,     0,    -1,    -2,     0,     1,     3,    -1,    -2,    -2,    -1,     2,     0,    -2,    -2,    -1,    -2,     2,     1,     2,    -4,    -9,    -9,   -10,    -8,    -7,   -11,   -10,   -12,   -15,    -9,    -8,    -4,    -2,    -2,     1,    -1,    -1,     1,     2,    -4,    -5,    -3,    -3,    -7,    -5,   -24,   -19,   -28,   -25,   -20,   -20,   -20,    -3,    -2,     4,     5,    -5,     6,     3,    -2,     6,    -9,    -5,     2,     1,     1,     2,    -7,     8,    12,    -8,   -27,   -21,    -4,     2,     8,   -14,   -17,    -3,    -9,    14,    10,     5,    19,    15,    17,    32,    25,    18,    -8,     8,     6,     0,    -1,    -1,    -9,     9,   -27,   -24,   -13,    -8,   -26,    -7,     9,    -7,    -6,   -12,     4,    12,    12,    20,    37,    17,    18,    22,    38,    18,   -12,     3,    -9,    -7,     1,     2,   -12,    12,   -30,   -10,    -9,    -8,     0,     9,    11,     2,    -8,   -13,     5,     5,    13,    18,    22,    23,    29,     6,    18,     6,    -7,    -9,   -13,   -14,     1,     1,    -3,   -28,    -4,    14,    14,     6,    12,     6,     6,     0,     0,   -12,    -1,     1,     3,    -1,    16,    26,    16,     0,    14,    12,    19,    19,     3,     4,    -1,    -4,    -2,   -31,   -17,    -7,     7,     3,     1,     0,     0,    11,    -9,    -5,    -6,   -19,    -5,    -7,    11,    20,     7,     9,    30,    25,    22,     6,    10,    18,    -8,    -9,   -13,   -33,   -10,   -12,     5,     8,    -2,    -1,   -11,     5,     7,    -1,    -7,   -14,   -19,    -3,    -6,    19,    13,    14,    25,    22,    14,     2,     8,    11,     2,     0,   -13,   -18,    -9,    -7,    -4,     5,     3,    -7,     3,     2,    -2,    -1,   -11,   -19,   -19,   -15,    -3,    16,     2,     4,    13,    18,    18,     9,     1,    -1,    -1,    -3,    -9,   -28,     5,     0,   -12,   -13,     0,     7,   -11,     9,     8,    -7,   -11,    -8,   -22,   -18,     5,     3,     3,    14,    12,    20,    23,     4,    -7,    -7,    -1,    -2,     1,   -20,     5,   -10,     1,   -10,     3,    -4,    -6,    -1,     3,    -6,   -15,    -8,     9,     4,    -1,     2,   -11,    -4,    10,    17,    21,    14,    -8,    -6,     1,     0,    -4,   -15,    18,    -3,    -3,     7,     6,     9,    19,     2,    14,    -4,    -4,   -12,    -3,    -5,    -3,   -11,   -12,   -10,     0,     4,     6,    17,    25,    -8,     2,    -1,    -2,   -18,     2,     3,    -3,    12,     0,     0,     6,     8,    11,    -4,    -9,    -2,    -4,    -9,   -14,     4,    -4,    10,   -11,   -16,   -16,   -11,    18,    -8,     0,     1,    -6,   -19,    10,     5,    16,    -2,     0,     9,     9,     9,    -5,     2,     3,    -2,    -1,    -6,     3,    -1,    10,    -3,     8,     0,    -3,   -19,   -19,    -8,     4,    -1,   -12,    -4,    14,    19,     2,     8,    -4,     4,     8,    -2,    -3,     1,    -4,   -18,    -6,     3,    -3,    -3,    -5,    -3,     1,     6,     5,    -9,   -15,    -4,     0,    -3,   -14,    -5,     5,    16,    21,     8,     2,     4,    -6,    -7,   -10,     1,    -5,   -10,   -16,     1,    10,     2,    -7,     8,    12,    -1,   -12,   -25,   -22,    -6,     1,    -4,   -17,    -3,    12,    21,     8,    27,    15,     1,    -2,    -5,   -19,    -4,     3,   -10,    -5,    -8,     3,     2,     8,     2,    10,     1,    -8,   -25,   -38,   -23,    -5,    -3,   -17,    -1,     3,     6,    23,    18,    17,     8,   -12,    -4,   -16,   -18,     6,     3,    -4,   -13,    -5,    -4,    10,    -2,    -2,     2,   -11,   -25,   -22,   -19,     2,    -6,    10,    14,     1,    13,    20,     9,     0,     2,     3,     3,    -8,   -13,     3,     8,     4,     4,    -6,     0,   -10,     6,    -1,     7,     9,    -5,   -25,   -15,    -1,    -5,    16,    12,    15,    28,    12,     1,     5,    12,     2,     6,    -5,     5,     1,    13,     4,     3,     3,     4,    -5,     0,    -1,     9,   -11,     5,   -31,     1,    -1,    -3,   -14,    -2,     9,    18,    27,     6,    -5,     2,    -4,    -7,     3,     1,    -2,    -7,     0,    -1,     5,    -1,     2,     5,     5,     2,    -7,     4,     4,     0,     1,    -1,   -25,   -13,    -3,     2,    -3,    11,     0,     4,    -2,     6,    -5,    -5,    10,     5,     6,    10,    -2,    11,     5,    -2,    -8,     2,     2,     8,    19,    -1,    -1,    -1,     8,    -4,     3,     1,     6,     4,    -4,    -4,    14,     7,     8,    12,     8,     8,     6,     4,   -21,    -8,     2,    -5,   -11,    -2,    12,    10,    23,    -2,     0,    -2,   -14,    -9,   -17,    -2,     0,     0,     8,    10,     4,     5,     9,    13,    11,     8,    12,     5,     5,     0,    -4,    -4,    -5,   -14,     4,   -23,   -10,    -1,    -1,    -2,    -3,    11,   -25,   -23,     0,    -5,     1,    -5,    -2,    -2,    -1,     4,    -8,    13,    14,    12,     4,    13,    12,    12,    23,    21,    16,    -6,    -1,    -2,    -1,     2,     1,    -9,   -14,   -17,   -22,   -31,   -15,    -6,    -4,     6,    13,    31,    16,    22,     6,     2,    -6,     6,     1,     1,     0,   -17,    -7,    -1,     0,     1,    -2,    -2,    -2,    -1,     2,     4,    -3,    -4,    -5,    -5,     2,    -1,     3,    -2,   -25,   -12,    -4,    -2,    -8,    -6,   -16,   -20,   -14,   -12,    -2,     1,    -2,     2),
		    86 => (    0,     1,    -2,     2,     2,     0,     1,    -1,     0,     0,     1,     1,     9,     6,    -1,     0,     1,    -1,    -1,     0,     1,    -1,     0,    -2,     2,    -1,    -2,     0,    -2,    -1,    -2,    -2,     1,     0,     8,     9,     9,    10,    10,     4,    12,     8,   -13,     1,    -2,     7,     6,     9,    12,     4,     3,    -1,    -2,     2,     1,    -1,     0,    -2,     4,    -1,     6,     2,     9,     6,    11,    13,     8,     6,    11,     6,     5,     1,     8,     8,    12,    13,    21,    18,    13,     6,     2,     6,    -2,    -2,    -2,    -1,    -8,    -1,     2,     9,    17,    19,    18,    17,    20,    16,    10,    15,    10,    -4,     1,    13,    12,     0,     4,    17,    19,    18,    13,    -5,    -1,    -1,     0,     2,   -17,    -8,     8,    17,    21,    14,     5,    12,    19,    10,    15,    -2,     4,    -6,     8,    10,     3,     6,    15,    -7,     1,     8,     7,     8,    -3,     5,    -1,     0,   -11,   -10,     9,    11,     8,    10,    13,    15,    17,     6,     9,    -1,     3,    -1,    10,     5,    -9,    -7,     2,    -4,     8,     9,     9,    15,     6,     3,    -2,     0,     0,    -4,     9,     3,    13,     4,     2,    15,    19,     5,    -5,    -6,    -5,    -4,     2,    -3,     5,     3,     3,    13,     4,     6,     6,     6,    -1,    -5,     0,     2,    -1,    -7,     4,     5,     2,    14,     9,    17,     8,     2,     0,    -7,    -1,    -7,     0,     4,    16,     3,    11,     5,    -3,    -8,     5,    -1,    -6,   -12,    -1,    -1,    -8,   -12,    11,     4,    -3,     5,     8,     8,     8,     0,     4,    -7,     4,    -5,    -9,    16,    -8,     4,     9,    16,   -12,   -15,   -17,   -23,   -15,   -20,     1,    -2,   -12,   -13,     4,    -2,    -5,     1,     6,    -1,     1,     5,     3,    -3,     0,    -6,   -10,   -17,   -10,     6,     7,    -5,   -15,   -12,    -4,   -20,    -7,   -17,     1,     0,    -9,   -15,     3,    -7,    -6,    -6,    -4,     1,     2,    -6,     4,     1,     2,   -12,   -15,   -17,   -10,     6,     0,    -8,   -17,   -16,   -16,    -6,    -8,   -25,     0,    -1,    -9,   -19,    -2,    -1,    -1,    -9,   -15,    -6,    -3,     5,     6,    -4,   -10,    -8,    -6,    -5,     6,     6,     0,    -7,   -11,    -7,   -10,    -6,   -19,    -7,    -1,     0,    -2,   -12,    -3,     2,    -4,   -11,   -24,    -2,    -1,     2,     0,    -3,    -5,    -1,     7,    19,    16,     4,    -6,     3,    -9,    14,     5,    -6,   -19,    -7,    -1,     0,    -3,   -12,    -3,    -6,    -8,   -24,   -30,   -11,    -4,    -3,    -6,     3,    -6,     3,    10,    -5,    -2,     5,    -5,     5,    -1,    19,    -9,   -10,   -16,    -1,    -2,     0,    -3,   -14,   -12,    -5,   -15,   -14,   -18,   -10,    -1,     0,     0,    -3,     1,     5,     1,    -6,   -12,    -6,    -6,     0,     6,    14,    -2,    -2,    -2,     0,     2,    -2,    -4,   -13,   -18,   -11,   -10,    -4,   -27,   -22,   -10,     0,    -3,    -4,    -7,     6,     4,   -10,    -8,     2,    -3,     1,     2,    -1,     0,     6,   -13,   -20,     2,    -3,    -6,   -23,    -4,     6,   -10,    -3,   -19,    -9,    -4,    -2,    -7,   -12,    -6,     1,     4,    -1,     4,    -2,    -2,     3,     2,     2,     4,     4,   -13,   -17,     0,     0,    -6,   -20,     4,    -6,     0,     3,    -2,     2,     5,     8,    -7,   -15,    -9,    -4,     2,    -2,     6,     1,    -2,    -5,    -1,    10,    12,     8,    -9,   -22,     0,    -2,    -4,   -24,    -4,    -8,    -2,     2,     2,    11,    16,    13,     7,    -4,    -2,     3,     4,    10,    10,     4,     8,     8,    -4,     6,     9,    13,    -9,   -10,     2,    -7,   -20,   -18,     0,    -6,     7,     9,    12,     2,    22,    20,    15,     3,     6,    -1,     0,    -3,    -1,     4,     4,     1,    -1,    -2,     1,     0,    -7,    -4,     2,    -6,    -5,   -15,    -6,    -7,    -8,    19,    16,    17,    26,    21,    21,    12,    16,    17,    -1,    -9,    -2,   -11,     2,    -1,    -4,    -6,   -14,    -3,   -15,    -1,     2,     0,   -14,    -7,    -7,   -14,    -8,    12,    37,    22,    17,     8,    12,    12,    14,     4,    -3,    -4,    -5,     8,     5,    -2,    -3,    -4,   -23,   -19,   -13,    -2,    -2,    -2,    -3,    -9,   -15,   -22,   -16,     2,    10,    17,    13,    11,     8,     1,     2,    -2,    -8,    -6,    -5,     0,     6,     6,    -3,    -8,   -30,   -18,   -11,    -1,     2,     0,    -1,   -13,    -8,   -11,   -12,   -12,   -13,    -1,    -1,    -2,     0,    -2,    -2,     5,     5,   -13,    -4,    12,     8,    -4,   -13,   -21,   -24,    -8,    -9,    -2,     0,     2,     1,     0,    -6,    -5,    -2,   -14,   -25,   -25,   -25,   -31,   -16,   -22,   -15,     0,    13,    16,    11,    -9,    -5,   -20,   -11,   -12,    -7,    -3,     1,     2,     2,     1,    -1,     1,    -2,    -8,   -10,   -17,   -13,    -9,   -11,     0,     8,     3,    -6,    -9,   -10,    -9,    -9,    -4,   -18,    -9,   -11,   -15,    -5,     0,     2,    -1,    -2,    -1,    -1,     0,    -4,    -6,    -1,     1,     0,     1,    -4,    -6,    -2,     2,    -4,    -5,     0,     2,    -1,     0,    -6,    -3,    -3,    -4,    -2,     0,    -2,     0,    -1,    -1,     0,     2,    -1,    -1,     1,     1,    -2,     0,    -2,     3,    -2,     0,     0,     0,    -1,     2,    -3,     0,    -2,    -3,    -1,     2,     2,    -1,    -1,     1),
		    87 => (    1,    -1,     2,     1,     1,    -1,    -2,     0,     2,    -2,     2,     1,     2,     0,     0,     0,     2,     2,    -1,     1,     1,     1,     1,     1,     2,    -2,     1,    -2,     2,     0,    -1,     2,     0,     1,    -2,    -2,     1,     0,     0,    -6,    -9,    -6,    -1,   -11,   -20,   -18,    -1,    -1,    -1,     1,    -1,    -3,     0,     2,    -2,    -1,     0,    -1,     1,     1,    -3,    -1,     1,    -2,    -2,    -3,   -12,   -22,    -3,    -3,     0,   -16,    -6,    -7,    -6,    -3,     0,    -2,    -1,    -1,    -1,     2,     2,     2,     1,     0,     2,    -4,    -3,    -5,   -11,   -19,   -14,   -12,    -7,    -9,   -14,   -12,    -9,   -11,   -12,    -9,    -6,   -14,    -5,    -5,    -7,    -1,    -1,    -3,     0,     2,     2,     2,     0,     1,   -14,    -9,    -6,   -24,   -24,   -21,   -43,   -16,    -8,    -2,    -3,    -7,   -19,   -15,   -14,   -15,   -15,    13,     1,   -13,   -16,    -8,    -3,    -1,     2,    -2,     1,   -20,    -8,    19,     2,    12,     6,     9,    -9,   -22,   -25,    -1,    -9,   -15,    -8,   -15,   -19,   -10,    -8,    -6,    -9,   -23,    -9,   -14,    -1,     0,     2,    -1,    10,    14,    11,    18,    12,    13,     7,     9,    20,    -2,     1,   -13,   -12,   -13,    -6,    -3,   -10,     1,    -1,     0,     6,   -19,    -3,   -13,    -6,    -5,     0,     4,    14,     0,    22,    20,    24,    29,     4,    26,    23,    10,     9,     6,     4,    -4,    -7,    -1,     4,     1,     3,    -1,    21,     5,    -4,   -14,    -4,    -7,    -9,    -3,     1,     2,     2,     9,     4,    19,     4,    12,    12,    10,    17,     4,     7,     6,     1,    -2,    -4,     2,    -1,    -2,    16,     0,   -11,   -20,   -12,    -9,    -2,     1,    18,     8,     7,     1,     1,     7,     6,     1,     1,     4,    19,    10,    16,     8,     2,     1,    -3,     1,     5,     0,    10,     5,   -20,     3,    15,    30,    -2,    -8,     7,    -2,    -8,    -6,    -4,    -7,     5,     1,    -4,   -10,   -10,     2,    -3,    -1,     2,     9,     7,    -4,     6,    -8,    -6,    -6,    -7,    11,    15,    28,     2,    -5,     6,    -6,    -8,   -14,    -7,    -6,    -7,    -4,   -16,    -3,   -14,   -20,    -6,    -1,    -3,    -2,    -9,    -5,     2,   -12,     1,     5,   -15,   -20,   -14,     4,     1,     6,    -9,   -11,    -9,   -15,   -15,   -17,   -20,   -26,   -31,   -12,   -16,   -12,    -9,     4,     5,     0,     3,     3,     2,    -3,    -8,   -10,   -35,    -5,   -17,     3,     0,     0,     5,   -13,   -24,    -9,    -8,   -13,   -14,   -11,   -14,   -11,    -5,   -10,    -4,    12,    -3,     5,     5,     0,   -15,     8,    -7,    -1,   -18,   -11,   -14,    -8,    -3,     2,    -2,    -5,    -7,    -5,     0,     0,    -8,    -7,     4,     2,     6,     4,     6,     5,    -8,    13,     6,    12,    -1,     8,    -2,     5,     2,   -12,   -10,    -1,     2,    -1,    -2,     0,    -2,     0,    -1,    -4,   -12,    -2,    -7,    -4,    -1,     3,     2,     3,    -9,     7,    10,     1,   -13,    16,     0,     7,    -2,   -11,    -3,    -9,     2,    -4,     0,    -8,    -3,    -3,    -5,    -3,    -6,     0,     8,    -4,     5,    10,     0,    -2,    -2,    -2,     4,     1,     5,     2,    -4,    -9,     2,   -24,   -18,    -3,     0,     2,   -14,   -14,   -15,   -10,     8,    10,     2,    10,    12,     3,     6,     0,     0,    -4,     5,    -3,   -12,    -5,     5,     1,     2,    -3,     1,   -10,     4,   -11,     3,     1,    -2,    -8,   -11,    -1,    -8,    10,     1,     2,     2,    -1,     0,    -1,    -6,    -7,    -9,    -4,   -11,    -5,    -2,   -13,    -4,    -4,    -6,   -11,     9,   -11,     0,     2,    -2,    -2,   -10,   -16,    -5,     2,     2,    -2,   -10,     2,    -2,     3,     2,    -5,   -11,    -8,   -20,   -11,   -14,   -21,    -9,    -3,    13,    -2,   -13,    -6,    -2,     9,    -3,    -8,   -26,   -22,   -11,     0,     3,    -3,    -9,     4,    -2,     1,    -3,    -8,    -5,   -22,   -26,   -16,   -15,   -17,   -22,     1,     2,   -17,   -14,    -2,    -2,    -2,    -6,   -17,   -10,   -11,   -13,   -22,   -17,   -13,    -6,    -6,     1,     2,    -6,    -7,    -8,   -16,   -20,   -14,   -18,   -12,   -17,     0,    -2,    -8,    -3,     1,    -3,    -2,    -4,   -22,     1,    -5,    -7,    -3,   -18,   -15,    -3,    -2,    -2,    -6,   -11,     1,    -3,     1,    -9,    -7,   -12,   -36,   -29,   -19,   -10,    -3,   -14,    -2,    -2,    -1,    -8,   -27,    -3,    -1,     4,     6,   -18,    -7,     0,    -2,     2,     0,    -1,     2,    -5,    -2,   -17,    -6,   -11,   -15,   -27,   -12,   -11,    -6,   -14,     1,     0,     0,     5,    -2,     7,     8,    -3,    -4,    -3,    -7,   -13,     0,    -3,     1,    -1,    -4,    -9,    10,   -11,    -5,     4,     6,   -15,   -11,   -10,    -4,    -3,     1,     1,     1,    -7,     7,    -7,    -9,    -7,    17,     8,    -5,   -11,    -7,    -5,    -3,    -2,   -10,     0,    -1,    -4,     1,    -8,    -4,    -4,    -4,   -15,    -3,    -5,     2,     2,     2,    -2,    -9,   -32,   -24,   -28,    -8,    -1,    -7,   -10,   -16,   -12,    -4,     1,    13,     0,    -7,     0,   -14,     2,    -2,    -5,    -9,    -2,     1,     0,     2,    -2,     2,     2,     0,     1,     2,     0,    -6,     4,    13,    16,    11,    -3,    -6,    -9,    10,    12,    17,    14,    -3,    -2,    -1,    -7,     1,    -1,    -2,     0,    -2),
		    88 => (   -1,    -1,     1,    -1,    -2,     0,    -2,     2,    -1,    -1,     2,     2,     2,     1,     1,     1,    -2,     1,     2,     1,    -2,     2,    -1,     0,     2,     2,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -2,     0,    -2,    -2,    -2,    -4,    -7,    -6,   -10,   -25,   -27,   -23,    -5,    -4,    -5,    -3,    -4,    -1,     1,     1,    -2,    -2,     0,     2,    -1,     0,     0,     0,    -5,    -2,   -10,   -10,   -13,   -16,   -10,    -6,    -1,   -13,   -17,     5,     7,    -1,   -11,   -15,   -17,    -2,    -3,    -4,    -1,     0,     1,     1,    -2,    -6,    -5,   -20,   -17,   -21,   -14,    -7,     5,     7,     8,     2,    -3,   -12,   -18,   -25,   -12,    -4,     4,    10,     1,     6,     6,    -6,    -3,     2,    -2,     1,     3,    -1,   -10,   -22,   -16,   -16,     8,     5,    18,    18,     3,   -17,     0,    -8,    -8,     2,    -1,   -10,    -8,     2,   -10,     3,     7,     6,     4,    -4,     0,    -2,    -8,    -7,   -20,   -17,   -19,     1,    -6,     6,    13,    11,     3,     9,     2,    10,    11,    14,     6,     0,    -1,    -5,   -15,   -13,     8,     3,    -7,    -9,     2,     2,   -16,   -15,     4,   -13,   -18,   -11,    -2,    -3,     5,     3,    -5,    -1,     7,    10,     9,     4,     6,    -9,    -4,     0,     6,     5,     2,     7,    -1,    -3,     1,   -15,    -8,     4,     8,    -7,   -10,    -1,     4,     6,     2,     0,    -4,    -2,     1,    15,    15,     5,    -2,    -6,     5,     5,    11,    14,     6,     3,     2,   -10,    -8,   -10,    -8,    20,    11,     1,     5,     6,   -11,     2,     6,     0,    -2,     2,     3,     7,     6,     4,     5,    -3,    -3,    -7,    -1,     8,    -4,     5,     8,     2,     2,    -7,   -12,    11,    22,     0,     1,    -7,    -4,     2,     2,    -8,    -4,    -5,     1,     6,    -2,    -8,    -2,     3,     1,    -1,    -6,     1,    -2,    15,    21,   -15,    -3,    -7,   -15,   -10,    11,    -1,    -3,     0,    -9,   -11,   -10,   -12,    -6,     8,     9,    -4,   -18,   -13,   -10,    -8,    -1,    -8,     4,     5,     7,     6,    15,   -13,     2,    -4,   -11,    -5,     8,    -1,     7,    -4,    -7,    -5,   -16,    -8,    -1,     7,     0,   -22,   -20,   -12,    -9,    -3,    -5,    -4,    -5,    12,     4,   -10,     8,   -12,     1,    -2,    -2,     3,   -11,    -1,   -14,   -18,   -10,   -11,    -3,     8,     8,     5,     6,     0,    -8,   -12,    -5,    -6,     3,     1,     6,     0,    -9,   -26,   -29,   -16,    -2,    -1,     0,    -6,   -13,    -7,   -12,   -10,    -6,    14,    14,    12,    17,     9,     0,     5,    -1,    -6,     2,    -5,     5,    12,     7,     2,   -17,   -23,   -22,     2,    -4,    -2,    -4,    -9,   -12,    -1,     5,    -6,     6,    17,    17,    20,    16,    10,     2,     5,    -2,    -4,     0,     9,    11,    10,    -3,   -10,    -9,     2,   -12,    -6,    -3,    -1,    -6,    -3,   -15,    -3,    12,    12,    14,    22,    25,    13,    11,    14,     5,     2,     4,     1,     7,     7,     9,     4,     5,   -12,   -10,    17,   -19,    -6,    -2,     0,    -7,    -7,   -11,    -7,    -4,    10,     5,    16,    20,    18,     6,    -2,    -1,    -1,     9,    19,    17,     4,    11,     7,     0,    -1,     0,     8,   -25,    -9,    -2,    -3,   -12,    -7,     2,   -12,   -14,     0,     2,     2,     7,     2,    -5,    -8,    -3,    11,     1,     3,     7,     6,     2,    -3,    -3,     4,     5,    -6,    -3,   -11,    -2,    -5,   -12,   -19,    -9,   -13,    -5,    -9,    -8,    -1,    -5,   -10,    -9,    -3,     8,    -2,     0,    -9,     2,    -5,   -16,   -14,    -5,     8,    -4,   -15,    -1,    -5,     1,     1,    -6,   -23,   -11,   -19,   -17,   -17,   -15,   -13,    -8,    -9,     1,     9,    11,     4,     9,    -5,    -5,   -10,    -9,    -1,     6,     2,    -8,   -19,   -11,    -7,    -2,     0,   -10,   -21,   -12,   -11,   -10,    -2,     1,   -12,    -6,    -7,     8,    10,    17,    11,     6,     3,    -8,     1,     5,     3,     1,     0,   -17,   -15,   -14,    -1,    -5,    -6,   -13,    -4,   -10,     0,     2,    -2,     0,    -1,    -7,    12,    27,    11,     8,    15,    10,     9,    -2,     1,     4,    -9,    -6,    -1,   -10,    -8,   -14,    -2,    -5,    -4,    -6,     1,    11,     5,    -2,    -6,    -7,     1,     2,    13,     7,     5,    20,    17,     6,    -2,    -2,    -9,     5,    -6,     5,     7,    -6,   -14,   -14,    -4,    -2,    -1,    -4,    -1,     5,     3,    -6,   -12,    -7,    10,    12,     1,     9,    20,    14,    11,     6,    -8,    -2,     0,     9,     2,     7,     9,   -20,   -16,    -9,     0,     0,     2,    -7,    -6,    -4,    -8,    -9,   -13,    -9,     2,    -2,     4,    17,    22,    15,     2,    -4,    -9,     3,    19,    15,     3,   -14,    -7,   -23,   -11,    -5,    -1,    -1,     0,    -7,    -1,   -25,   -17,    -1,    -7,   -16,   -16,    -2,    11,    10,    14,     5,     3,   -15,    -6,     1,     3,    -9,   -23,   -22,   -14,   -12,    -5,    -9,    -2,     2,     0,     1,   -10,    -9,   -10,   -16,   -12,    13,     8,    -9,    -5,    -3,     5,    -2,   -21,   -10,    -7,   -14,   -14,   -27,   -21,   -11,    -8,    -2,    -1,     1,    -1,     0,    -1,     1,     1,     0,    -4,    -3,     0,   -13,   -18,   -10,    -3,    -3,   -11,   -21,   -15,   -16,   -13,    -8,    -5,    -2,    -1,    -4,    -2,     2,     2,     0,    -1),
		    89 => (    0,    -2,     1,     2,    -2,     0,     2,    -1,     1,     0,     0,     0,    -2,     1,     1,    -2,     2,    -2,     0,     1,     0,     0,     0,     2,     1,     2,     1,    -1,     1,     1,     2,     2,     1,    -1,     0,    -1,     0,     2,    -1,    -6,   -12,    -8,     0,    -1,    -3,    -1,    -9,    -7,     1,    -4,    -3,     0,     2,     0,     1,     1,     2,     1,    -2,   -10,    -5,     0,    -1,    -4,    -3,     0,    -3,    -9,     0,    -3,   -14,    -6,    -4,    -3,    -5,    -5,    -7,    -4,    -4,    -1,    -3,     0,     0,    -2,     0,     2,     2,    -6,   -10,   -12,   -10,   -12,    -3,    -5,    -1,    -7,    -7,   -10,   -14,   -12,   -10,   -10,   -17,   -11,    -7,    -7,    -6,    -2,    -2,    -2,     1,     2,    -1,     2,    -1,    -2,    -6,    -3,   -13,     2,    -8,    -4,    -5,   -11,   -19,   -15,    -9,    -9,    -4,    -4,    -9,   -16,   -18,    -9,    -5,    -4,    -1,   -12,    -2,     2,    -1,     1,     1,    -5,     1,    -1,    -3,    -5,    -5,    -8,   -18,    -6,    -7,    -6,     0,    -2,     1,    -7,    -4,    -9,    -1,    -3,   -10,    -6,    -1,    -5,    -5,    -1,     1,     0,    -2,    -7,     0,    -3,   -10,   -10,   -23,   -11,    -8,    -9,    -5,     5,    17,    10,     5,     7,     0,     1,     5,     0,    -8,    -9,    -5,    -8,    -4,    -5,     1,     0,    -5,     0,    -7,   -14,   -18,   -16,   -24,    -1,    -5,     6,     7,    -1,    -5,     7,    -1,     0,    -5,    -1,    -2,    -3,    -8,    -7,   -14,    -6,    -1,    -4,    -8,    -6,    -3,    -8,    -2,   -15,   -12,   -24,    -8,   -11,     6,     0,    -6,    -1,     0,   -21,    -8,    -1,    -2,    -3,     2,    -9,    -6,   -13,   -19,    -5,    -4,     0,     1,    -1,    -4,    -6,   -15,   -18,   -11,   -18,     0,     5,    -1,     6,    -3,    -4,     3,   -10,   -10,    -4,    11,     4,     3,   -10,    -8,    -4,    -8,   -18,    -2,    -8,     2,    -5,    -8,     0,    -3,    -6,    -9,     5,     5,     2,   -12,    -8,   -18,   -14,    -8,    -9,   -17,   -11,    11,     1,    -3,   -14,    -6,     1,    -9,    -2,    -3,    -6,     0,   -17,    -2,     7,    -2,    -7,    -6,    -2,     4,    -3,    -8,   -22,   -13,    -2,    -5,    -9,   -10,     0,    -7,     0,    -1,    -5,    -3,     7,   -11,    -5,    -2,    -7,    -2,    -3,     2,     6,     3,     3,     2,    -1,     9,    -5,    -9,   -18,    -5,   -12,   -19,   -12,    -7,    -5,   -14,    -2,     0,     6,    -1,     3,   -22,    -9,    -2,    -3,    -2,   -11,    -8,    11,    10,     5,     2,     0,    -3,   -15,    -8,   -10,   -17,   -13,    -5,    -3,     4,   -13,   -13,    -2,    -2,     7,     0,    -7,   -15,    -9,    -3,    -2,    -3,    -8,   -12,    -1,     6,     4,     4,     2,    11,   -14,    -6,   -21,   -15,   -10,    -7,     4,     2,    -8,     6,     6,     0,     2,     4,   -17,   -11,    -6,     3,    -2,     0,    -2,   -11,    -3,     1,     1,     8,     5,     6,   -11,    -5,   -21,   -18,   -17,    -9,    -7,    -9,   -13,     5,     5,    11,     4,     2,   -25,   -18,    -5,     2,    -1,     2,    -1,   -12,    -9,     6,    -7,    11,    -1,     1,    -5,     6,    -5,     0,    -4,    -9,   -12,   -15,    -7,    13,     5,     7,    -6,    -4,   -20,    -8,    -9,    -1,     1,     1,    -1,    -9,    -8,     8,    -8,     0,    10,    -9,     0,    -2,    -2,    -3,   -13,    -5,    -1,     1,     0,     5,     3,     5,    -6,    -4,   -11,    -3,    -4,    -8,    -3,     0,     2,   -10,    -5,     8,     7,     6,    -2,    -6,    -2,    13,     5,     8,     2,     4,    -5,    -7,     6,     8,     3,    -5,     3,     5,    -9,   -18,     0,    -9,    -7,    -2,    -1,    -6,    -3,     4,    16,    13,    20,    -6,     2,    12,    25,     6,    -3,    -7,    -2,    -2,     1,    11,    -8,    -2,    -5,    -2,   -10,    -6,     5,   -10,    -1,     1,    -3,    -4,    -5,    -1,     7,     4,    -2,     3,     4,    -2,     0,    -1,    -7,   -17,    -8,    -6,     5,    12,    -6,    -4,     1,    -3,    -4,    13,     5,    -9,     0,     1,     2,    -9,    -6,   -14,    -4,     2,     9,     5,     1,    -1,    -3,    -7,    -7,    -6,     0,     2,    -1,     6,     2,     4,    -9,     0,     1,    16,    -4,   -19,     2,    -1,     1,    -3,    -5,    -8,    -8,   -10,   -10,    -1,    -2,    -6,   -10,    -4,   -12,     7,     3,    -3,    -3,     0,     1,     3,    -2,     6,    -3,    13,     3,   -15,     1,    -1,    -1,    -2,     3,    -9,   -10,    -9,   -12,   -12,   -21,   -23,   -20,   -17,    -4,     4,    11,    -8,    -3,    -9,     7,     2,     6,    17,    -1,    14,     5,    -9,    -1,     1,     0,    -5,     1,    -1,    -2,    -5,    -3,    -8,   -10,   -19,   -18,    -4,    14,    -3,    -1,     0,    -5,     2,     6,    10,    12,    16,    11,    12,     4,    -1,     2,    -1,    -2,     8,    -6,    -5,     2,    -2,    -7,    -6,   -10,     0,     3,     9,    13,    -1,    -8,   -10,   -13,    -4,    15,    19,    12,    20,     9,     8,    -4,    -5,     1,     0,     1,     1,     3,     6,     1,     0,     2,    -1,    -1,    -1,    -1,    -5,    -9,    -5,   -17,   -22,   -11,    -2,     2,    14,     8,     6,     7,    -1,     0,     2,     2,     0,    -1,     0,     2,    -4,    -1,    -1,     0,     0,     1,     2,     2,    -1,    -1,    -6,    -3,    -8,   -14,   -10,   -10,    -6,    -8,     1,    -3,     1,     0,     0,     1),
		    90 => (   -2,     1,    -1,     1,     1,    -1,    -2,     1,     0,    -1,     1,     1,     0,     2,     0,    -2,    -2,     2,    -2,     2,     0,    -1,     1,     0,    -2,     2,     1,    -2,    -2,     0,    -1,     2,     0,     1,    -2,    -1,    -2,     0,    -2,    -2,     2,     2,    -3,    -2,     0,     1,     0,     2,     0,     0,    -2,     0,     2,     1,     0,    -1,     1,    -2,     0,     3,     0,     1,    -5,    -3,    -4,    -6,    -5,    -3,    -5,    -6,    -5,    -2,    -1,     2,    -1,    -3,    -1,     0,    -1,    -4,    -3,     1,     0,     0,     0,    -2,     0,     2,    -3,     0,    -3,     0,     1,    -2,    -3,    -5,    -9,    -4,    -3,    -3,     2,     5,     5,     0,     0,     0,    -2,    -4,     3,     2,     0,     0,     2,    -1,     2,    -4,    -3,    -9,    -6,     4,     2,     1,    -1,    -7,    -5,    -5,    -4,    -3,     6,     9,     4,     8,     7,     0,    -1,    -3,     0,    -2,    -3,     2,     2,     1,    -2,     2,    -1,    -2,     2,    -8,    -3,    -4,    -5,    -2,     1,     1,    -4,    -3,     1,    -3,     1,    10,    10,     1,    -3,    -3,    -3,    -2,    -2,    -7,     2,    -1,    -4,    -4,    -2,    -6,     2,     4,     1,    -5,    -4,    -1,    -3,    -5,    -3,    -5,     5,     2,     1,     4,     7,     5,    -3,    -3,    -4,   -10,    -2,     0,     1,    -3,    -5,    -5,    -1,     3,     8,     2,    -4,     4,     3,     2,     4,     2,     0,     9,     2,     6,    12,     3,     0,     3,     7,     0,    -2,     0,    -6,     1,     1,    -2,     5,    -5,     4,     5,     3,     6,     3,    -6,    -4,     2,     6,    -5,    -2,    -4,     1,     4,     2,     4,     9,     8,     5,     5,    -4,    -3,    -5,    -4,    -2,     0,     3,    -1,    12,     2,    -3,    -1,     3,     4,    -3,   -12,   -13,   -10,   -10,   -10,    -5,    -2,    -1,     0,     1,    10,     6,    -2,     3,    -4,    -1,    -2,     1,     1,     1,     0,    -1,     9,     9,     8,     7,     1,   -12,   -10,   -11,    -8,    -5,     1,   -11,    -7,    -7,    -4,    -5,    -6,     7,     2,    -2,    -4,    -5,    -1,     2,     7,     1,    -2,     6,    10,     4,    -6,     1,   -10,   -12,   -17,   -13,     1,     3,     3,    -6,    -7,   -11,   -16,   -13,    -8,     1,     1,     8,     0,    -1,    -1,    -1,    -1,     2,    -2,     7,     5,     3,    -4,    -1,    -8,   -14,   -17,   -11,     1,    -2,    -4,   -15,   -18,   -11,   -11,   -12,    -5,    -1,    -3,     5,     4,    -2,     2,     2,    -2,     1,     1,    12,     2,    10,    -5,    -6,   -12,   -19,   -19,    -9,    -5,    -2,    -6,   -14,   -11,   -14,   -13,   -13,    -6,     1,     5,     6,     2,     0,    -4,     1,    -1,    -1,    -8,    13,     8,    -3,   -10,   -14,   -16,   -14,   -12,   -12,    -9,    -5,   -13,   -12,   -10,   -11,   -12,   -11,    -6,    -8,    -3,    -6,     4,    -4,    -2,    -2,     2,     0,     1,    11,     5,    -2,    -7,    -9,   -14,   -11,   -12,    -6,    -6,    -7,    -2,    -5,   -10,    -9,   -10,   -11,    -5,     1,    -1,    -4,     1,    -3,     0,     2,     1,    -4,    -1,     7,     9,     6,    -1,    -5,    -7,    -8,    -7,    -9,    -7,     6,    -5,    -5,   -15,   -15,   -14,    -6,   -10,    -3,    10,     0,     4,    -6,     3,     1,    -1,    -4,     6,    10,     8,     8,     8,    -5,    -7,     2,    -1,    -5,    -6,    -4,    -8,   -15,   -15,   -15,   -13,    -9,     0,     6,    -1,    -2,     4,   -14,     2,     1,    -1,    -2,    -1,    15,     4,     4,     8,    -2,    -2,     0,    -6,    -3,    -5,   -12,    -6,   -12,   -12,   -17,   -10,    -5,     5,     1,     3,     1,    -2,    -3,    -1,     2,     1,     2,    -1,     9,     1,     2,     4,    -2,     1,     3,    -2,     0,    -4,    -4,    -6,    -9,    -3,    -4,    -1,     6,     0,     1,    -4,     1,    -8,    -4,     1,    -2,     0,     2,     0,     7,    -4,     7,     4,     1,    -6,    -4,     2,    -4,     1,     3,    -1,     5,     6,    -7,    -2,     1,    -2,     4,    -3,    -1,    -6,    -1,     0,     1,     0,    -3,     0,     0,    -8,     1,    10,     1,     1,    -2,     4,    -4,     0,    -1,     0,    -5,     2,     1,     5,     3,     2,    -6,     0,    -5,     0,     2,     3,     2,    -1,    -1,    -4,    -5,    -3,    -7,     8,     3,    -3,     2,     4,    -4,     1,    -3,    -5,     5,     6,    -1,     2,     2,    -4,    -3,    -4,    -6,     1,     3,     3,     2,    -1,    -1,    -5,    -3,    -4,     3,     7,    -2,    -5,    -2,     0,     2,    -6,    -2,    -1,    -6,    -1,    -4,     2,     0,     0,     0,    -6,    -8,    -6,    -6,    -1,    -1,    -2,    -2,    -2,    -4,    -2,     9,     7,     5,    -5,    -1,    -2,    -5,     3,     6,     4,     1,     3,     4,    -4,    -4,     0,    -1,    -3,     0,     0,    -1,     2,    -2,     1,     1,     0,    -3,    -2,     6,    10,    10,     2,     1,     0,    -4,    -4,    -7,     1,     0,    -4,   -11,   -15,   -13,    -9,    -8,    -5,    -1,    -2,    -1,    -1,     1,     2,     2,     0,    -1,    -6,    -9,     0,    -2,     0,    -3,    -1,     1,    -6,    -5,    -4,    -7,   -19,   -11,   -10,   -11,    -7,    -3,    -8,     0,    -2,     2,    -1,     2,     0,    -2,     0,     1,    -1,     0,    -1,     0,    -2,     0,    -1,     2,    -4,    -3,    -1,    -1,     0,     0,    -2,     1,    -5,    -7,    -6,     0,    -1,     0,    -2),
		    91 => (   -1,     0,     1,    -1,     2,    -1,    -2,    -1,     2,     1,     0,     1,     2,    -1,    -1,     2,     3,     2,     2,    -1,    -2,    -1,     1,     2,     1,     2,     2,    -2,    -1,     1,     0,     1,    -1,     3,    -1,     0,     1,     0,    -1,    -1,    -1,    -5,    13,     6,     7,    -8,    -2,     0,    -1,    -1,    -2,     0,    -2,     1,     0,     2,    -1,     2,    -2,     1,     2,    -2,     1,     2,    -8,    -8,    -6,    -7,    -2,     5,     4,     9,    21,    13,    11,     4,     6,   -14,   -10,   -13,    -1,     0,    -2,     0,     0,    -2,    16,     8,    -1,    -8,   -14,     9,     2,     2,   -11,   -18,    -8,    -1,    -2,     1,     4,     1,     2,   -11,    -4,    -8,    -7,    -8,    -7,    -1,     0,    -1,     1,    -1,    15,    14,    13,     1,    -4,     5,    10,     9,     5,     1,   -12,     2,    -4,     4,    -2,    -1,    -1,   -12,   -12,    -6,    11,     9,     8,    -5,    -4,    -6,    -1,    -2,     6,     4,    17,    14,     2,     3,    10,     1,    -3,    -2,    -5,    -6,   -11,    -3,    -3,    -4,    -6,    -4,   -14,     5,    12,    15,    12,   -10,    -5,    -8,    -2,    -2,    -7,     1,    17,     7,     5,    -1,   -10,    -8,    -3,    -4,     5,    -6,    -4,    -8,   -11,    -7,    -6,   -20,    -6,     7,    13,    12,     4,    -1,    -4,    -3,     2,    -1,    -9,   -10,    -9,    -7,   -10,     6,   -19,    -4,    18,    13,    11,    -3,     3,    -7,   -16,    -8,    -4,   -13,    -4,     9,    13,    15,     3,    -7,   -10,    -3,    -2,     0,   -11,    -8,    -9,    -9,    -9,    12,   -16,    -4,    16,    -1,    11,    -1,    -4,    -6,    -7,   -13,   -11,   -11,     6,     7,     7,     2,     2,    -5,   -11,    -4,     0,    -1,   -10,     0,    -8,   -10,    -6,    14,    -5,     2,     7,    -1,    -8,   -11,    -8,    -6,   -11,   -20,   -12,   -17,     2,     1,     6,     5,     2,    -2,   -10,    -5,    -2,    -2,    -7,     0,    -7,    -5,   -10,     5,     4,    -6,    11,     2,     1,    -1,    -3,    -7,   -16,   -15,    -3,    -4,     0,     1,     6,     9,    -6,    -1,     2,     5,    -2,     1,    -1,     0,     0,    -7,   -14,     6,   -10,    -4,    -1,    -6,    -3,    -7,     7,     0,   -13,    -5,    -3,    -4,    -3,    -7,     9,     5,    -6,     1,     0,    12,    -2,     2,    -7,     0,     2,    -5,    -6,    -7,   -13,   -11,     1,     0,    -4,    -7,     3,    -4,    -4,    -3,    -2,    -4,    -5,    -7,     1,     3,    -9,     4,     7,    13,     1,    -1,    -5,    -1,    -3,    -5,    -1,    -2,     1,    -3,    -4,    -6,     2,    -6,     1,     1,    -7,    -4,   -11,    -5,    -8,   -10,    -9,   -20,   -10,     9,     3,     2,     0,     2,     3,     3,    -4,    -8,     3,    -4,    -5,    -8,   -17,   -23,    -8,     7,     5,     5,     1,    -3,    -4,   -15,   -12,   -14,   -15,    -8,    -6,   -11,    -1,     1,     2,     1,    -1,    -1,    -5,   -17,    -8,    -8,   -11,   -18,   -26,   -22,    -8,     4,     9,    -8,   -10,     4,     1,   -13,   -14,    -7,   -14,    -8,   -18,   -16,   -13,    -3,     1,    -2,     0,    -1,    -5,    -4,    -8,    -9,   -12,    -2,   -10,    -7,   -11,    -4,    12,     3,    -5,     3,     3,    -4,    -4,    -1,     0,    -6,    11,   -17,   -12,    -3,     2,    -1,    -1,    -3,    -2,    -2,    -3,    -5,     2,     1,     6,     2,    -9,    -3,     8,    -2,     6,    -5,     4,     2,     8,     7,     6,    -2,     0,   -12,    -9,    -8,     2,    -2,    -2,    -9,    -6,     1,   -10,    -1,     7,    13,     7,   -11,   -13,    -9,     4,     2,     2,     9,     2,     3,    -8,    -3,     4,     0,     3,    -1,    -8,     0,    -2,     0,     5,    -9,    -5,    -1,    15,    16,    20,    19,    15,     2,   -15,    -1,    -2,     7,    10,     1,     3,    -7,    -1,     1,     9,    22,     7,     6,    -8,    -3,     2,     1,    -1,    -5,     5,    10,    15,    17,    11,    10,     8,     0,    -6,    -2,     5,     0,     6,     1,     1,     3,    13,    12,    15,     8,     5,     0,    -6,    -1,     4,     5,    -2,    -2,    -5,   -11,    -6,     0,    -2,    -5,    -6,   -11,    -3,     2,    -8,     1,   -10,    -6,     1,     5,     5,    -2,     7,     3,    -1,     8,    -4,    -1,     7,     3,    -7,    -4,    -4,     8,    -1,    -5,   -14,   -11,   -11,   -14,     2,     2,    -1,     4,   -10,    -4,    -2,    -1,     1,     0,   -11,    -8,    -2,     0,     3,    -2,    -2,    -2,    -2,    -5,     2,    10,    13,     5,    -1,    -2,     3,     1,    11,     3,    -9,    -8,    -8,     6,    -5,    -4,     9,     1,    -5,    -7,    -7,    -9,    12,     0,     2,     1,     2,    -3,     0,     0,     0,    -4,    -4,    -4,     2,     2,    -3,     1,    -8,   -17,    -7,    -9,    -6,   -14,    -1,   -13,    -5,    -5,   -12,     8,    10,     1,    -2,     0,     0,    -5,    -4,    -6,    -2,    -5,    -7,    -4,    -8,    -3,     0,     9,     9,    -6,   -14,    -9,    -9,   -10,   -18,   -12,    -5,    -4,     2,     1,    -1,     0,    -2,    -1,     1,    -4,    -4,   -11,   -10,    -7,    -4,    -4,    -3,     0,    -3,    -7,   -10,    -7,    -6,    -9,    -2,    -2,    -4,    -4,    -2,    -2,     2,     2,     1,     1,     1,    -2,     0,     2,    -2,     1,    -2,     0,    -1,     2,    -4,    -8,     2,    -2,    -2,     1,    -1,     2,    -1,    -2,     0,     0,     0,    -1,     0,     1,     1,    -1),
		    92 => (    2,     2,     2,     2,     1,     0,    -1,    -2,    -1,    -2,     2,    -2,    -2,    -3,     5,     4,     2,    -2,    -2,    -1,     0,     0,    -2,    -1,     1,     0,    -1,     1,    -2,     2,    -1,     1,    -1,     2,    -2,     3,    -4,    -8,   -11,   -16,    -3,    -5,    -2,     7,     9,     1,    -7,   -20,   -12,   -13,    -9,    -2,     2,    -2,     0,     2,     1,    -2,    -1,    -6,    -7,     0,     2,     1,     1,    16,    16,    19,     1,     5,    14,    23,    19,     8,    -8,   -18,   -10,    -4,    -9,    -3,    -1,     0,     2,     2,    -2,     0,     1,   -13,   -16,     7,    10,    13,     0,   -11,   -17,   -22,   -28,     0,    -3,     0,     2,    -9,   -21,   -14,   -12,    -3,     1,   -14,   -15,    -1,    -2,     0,    -1,    -1,    -4,   -11,     0,     5,    23,    18,    14,    23,     6,    -5,    -8,    -8,    -6,     3,    -7,    -2,     3,    -5,    -3,   -11,     1,   -11,   -18,    -1,   -12,    -4,     1,    -1,   -10,    -6,     0,   -10,    -8,     2,    14,     4,    11,     0,     3,     3,     6,     2,    -1,     2,     6,     8,     4,    13,    -5,    -8,   -16,     5,   -21,    -6,    -1,    -1,     2,     1,     5,    -2,    -2,    -3,    10,    -2,     3,   -11,     2,    -8,     1,     0,     6,     4,     9,     4,    -1,     5,    -2,    -7,   -27,    -3,   -19,    -5,    -2,    -2,     8,     0,     9,    22,     6,     3,     6,    -2,   -15,    -7,    -1,     3,    -4,     3,     8,    -7,     2,    -3,     2,    12,    11,   -19,     4,    11,   -13,    -8,   -11,    13,     8,     3,    -2,    18,     7,    -4,     5,     4,    -4,     4,     4,     1,    -1,   -10,    -6,    -2,    -9,     2,     1,    -8,     1,    11,    -3,    -7,   -21,    -6,     1,    -9,     2,    10,   -12,     1,     1,    -6,     1,    -5,     0,     6,     7,     6,    -5,     0,    -4,    -2,     0,    -4,    -1,    -4,    10,    -2,    -9,   -27,    -4,    -5,     2,     1,    -5,     5,    -6,    13,    20,     3,     3,    -7,    12,    -4,     1,     1,    -4,     1,    -5,    13,    -7,    -8,    -2,     3,    -5,   -18,   -10,    -8,    -7,    -8,    -1,   -10,     2,     1,    -4,     6,     9,     7,     3,     6,     7,    -2,    -9,   -13,    -3,   -10,    -2,    -8,     0,     4,     4,    -2,   -13,   -10,     5,     5,    -6,   -12,    -1,    -6,   -19,     0,    -7,     2,    18,     9,     0,    12,    -3,   -13,    -7,    -6,   -13,   -10,   -11,    -6,     7,    14,    -5,    12,    10,   -11,    12,     3,     0,    -3,    -2,   -11,    -7,    -2,    -2,     8,    29,     9,    -5,     1,    -3,    -2,    -3,     3,   -11,    -8,   -10,    -3,     5,     9,    -2,     3,    11,    22,    17,    18,    19,    -3,     2,    -1,    -4,     2,     9,    10,    18,    20,   -11,     7,     2,   -16,    -8,   -11,    -8,    -5,    -4,    -1,    -1,     8,   -14,     6,    19,    33,    27,    14,    12,     6,     0,    -7,    14,    16,    -1,     4,     9,     8,    12,     2,    -5,    -3,    -4,    -9,    -3,     0,    -3,    -8,    -3,    -7,     4,    11,    10,     9,    -2,    10,    22,    18,    -1,    -1,    19,    17,   -11,    -8,     2,    18,     8,    18,     8,     2,     7,    -2,    -5,    -4,    -3,    -8,    -5,     4,    -5,    35,    28,    18,     4,    20,    24,    13,     0,    -3,    17,    12,    -4,    -6,     4,    -3,    -3,    -3,     2,     1,     1,    -1,     5,    -3,    -5,    -1,    -2,    -3,    10,    37,    20,     8,     6,     9,     9,     9,    -1,     0,     3,     6,    -4,    -3,     2,    -7,     4,    -5,    -7,     1,     3,    -1,   -11,    -6,    -9,   -12,    -1,     9,    32,    28,    22,    16,    12,    10,    -3,     5,     1,   -10,     4,    -4,    -1,    -1,    -6,     0,     5,     4,     6,     9,    -5,    -6,     2,     7,    -5,   -13,     6,    18,    20,    27,    19,     8,    -1,    -6,     4,    13,    -2,    -6,    17,    -9,    -3,    -1,    -1,     0,     0,     7,    11,    13,     0,     0,   -10,     2,   -11,    -3,     6,    21,    26,    33,    13,    10,     5,     3,     2,    -2,    -2,    -1,    16,    -6,    10,    -3,     3,     0,    12,    18,    10,     0,     5,     5,   -11,     0,    -3,   -10,    23,    37,    27,    24,    30,     4,    -5,     3,    -3,    -2,     0,     0,    -5,   -12,    -4,     4,    -8,     0,    10,     9,     4,     5,    -7,    -1,    -7,    -4,     1,     8,    31,    31,    28,    22,    21,     9,   -12,     5,    -2,    -1,    -2,     2,     0,   -15,    -1,     5,     8,     3,     4,    18,     8,     5,     3,     3,    -6,    -5,    20,    37,    30,    22,    30,    27,    20,    12,   -10,     1,     1,    -2,     1,     0,   -12,    -5,   -10,   -17,     7,    -7,     0,     9,    10,     4,   -16,   -25,    -4,     3,    23,    32,    42,    30,    17,    24,    18,    -5,     6,     2,     6,     0,     2,    -1,    -5,    -2,   -14,   -27,    10,    -8,    -8,   -10,   -15,   -14,   -19,   -19,     3,     4,     3,    16,    27,     7,     2,     4,   -11,   -10,    -6,     0,     4,    -2,     2,     2,     2,    -2,    -4,    -8,   -17,   -25,   -12,   -28,   -33,   -25,   -23,   -34,   -33,   -27,   -27,   -25,   -20,   -32,   -10,    -6,   -12,     1,     1,     0,     1,     1,     1,     2,    -2,     2,    -4,    -3,    -5,    -4,    -3,    -3,   -12,   -15,   -11,   -13,   -15,    -7,    -7,    -6,    -4,    -5,    -4,    -4,    -5,     1,    -2,     1,     2,     2),
		    93 => (   -1,     0,    -1,     1,    -1,    -2,     1,     1,     1,    -1,     1,    -1,    -1,    -3,     1,    -1,     2,    -1,    -2,     2,     2,     2,     1,    -2,     1,    -2,    -1,     2,     2,    -2,     0,     0,     2,     1,    -1,    -1,     2,    -3,    -2,    -1,    -2,    -3,    -4,    -4,    -5,    -6,    -1,    -1,    -2,     0,     1,    -2,     1,     2,    -2,     1,     0,    -2,     0,     0,    -1,    -2,    -1,     0,   -10,   -12,    15,     4,    -5,   -10,   -16,    -9,    -9,    -7,    -8,    -6,   -17,   -13,   -16,   -10,    -1,     0,     1,    -2,    -1,     0,    -1,    -1,     0,    -4,     2,     7,    -9,   -15,   -19,   -16,   -19,   -23,   -30,   -15,   -12,   -15,   -20,   -13,   -12,    -9,    -5,   -12,    -4,    -3,     1,     1,    -2,     1,     1,     0,     5,    14,    16,    -6,    -4,   -20,    -3,    -5,    -5,   -14,   -24,   -22,   -22,   -20,   -19,   -20,   -15,    -5,    -7,    -6,    -5,   -10,     0,     2,     2,    -2,     1,     3,     7,    14,     1,    -5,    -2,     6,    12,     9,     9,    -5,    -7,    -4,    -7,    -6,   -15,   -21,   -13,   -12,   -12,    -5,    -3,   -13,    -4,     2,     1,     0,     1,     9,     5,    -8,     4,    11,     0,     9,    -4,     6,     3,    -7,    -9,   -11,   -14,   -13,    -9,   -18,   -15,   -12,   -12,   -12,    -9,    -1,    -8,     1,    -1,     5,    -1,     8,     2,    -2,    11,     4,     7,    -2,    -3,   -11,    -1,     1,    -3,     6,   -10,   -15,   -21,   -24,   -15,   -14,   -10,   -12,    -8,    -2,    -6,    -3,     2,     2,    -8,     4,     0,    -1,    -3,   -10,    -3,    -2,   -12,     0,    13,    14,    16,    11,    -3,   -21,   -25,   -25,   -19,    -9,   -11,   -12,    -8,    -4,    -4,     1,    -1,    -7,    -6,     1,    -3,     5,    -8,    -6,   -10,    -3,    -5,    10,    13,    14,    17,     1,   -10,   -29,   -26,   -26,   -17,   -10,    -7,    -3,    -6,    -8,    -7,    -2,     0,   -11,    -5,    13,     2,     7,     0,    -6,   -10,     1,     1,     6,    10,     9,     2,    -9,   -14,   -29,   -32,   -25,   -20,   -19,   -10,     0,    -4,    -5,    -3,     0,    -1,   -16,    -1,    17,    10,     2,    -3,    -1,    -3,     5,     8,     4,     8,     0,    -8,   -10,   -11,   -14,   -12,   -17,   -13,   -17,   -14,    -5,    -1,   -12,    -7,     0,     1,   -12,   -15,    12,    -4,    -1,   -12,    -8,     6,     4,    13,    11,     9,     2,     2,     1,   -10,   -10,     4,     0,    -1,     7,    13,     9,   -10,    -7,    -5,    -2,     1,    -5,   -11,    13,     8,     3,    -1,    -5,     6,     9,     9,     8,     8,     7,     3,    -6,    -1,    -2,     4,    -1,    -4,     4,     8,    12,    11,   -10,    -7,     0,    -3,     5,    -1,     6,   -11,    -8,    -7,    -5,     3,     9,     4,    -2,    -2,     1,    -6,    -2,     3,    -6,    -1,    11,    -1,     2,     2,    21,     8,   -13,    -5,    -3,    -1,     6,     1,     3,   -12,   -10,    -8,    -1,     5,     1,    -5,    -9,    -8,    -8,    -2,    -9,     1,     1,     0,     8,    14,     9,     8,     8,     2,   -11,    -2,    -1,     2,     2,     0,     1,   -13,   -20,    -8,   -13,     3,    11,    -9,   -10,   -10,   -18,   -22,    -7,    -9,    -9,     0,     4,    12,    12,    12,     1,    -2,    -8,    -8,    -4,     2,     0,    -3,     9,    -4,    -9,    -7,   -15,    -7,    -7,   -19,   -10,   -10,   -11,   -20,   -20,   -10,   -10,   -16,     7,     6,    17,     9,     6,    -2,    -7,    -3,    -1,    -2,    -1,     2,     1,     1,    -6,   -12,    -8,     0,    -6,   -20,    -9,    -4,   -10,    -9,   -16,    -8,    -1,    -3,     1,     6,     9,     6,     1,     3,    -6,    -4,    -8,     2,     0,    -4,    -5,    -7,    -5,    -6,     5,    -1,    -4,    -9,    -5,     2,     5,     2,    -4,     2,     8,    -3,     0,     2,     4,     2,    -5,     4,    -2,   -11,    -6,     3,     0,    -5,   -10,    -7,    -9,   -12,     0,     4,     5,    -4,     3,     4,     6,     8,     9,    12,    -1,    -5,    -3,     7,     7,     2,    -1,     6,    -4,    -3,    -2,    -2,    -1,     0,     1,     6,    -2,   -15,   -11,    -7,    -4,    -8,    -6,   -10,    -4,     2,     1,     1,    -4,    -9,    -1,     0,   -10,    -4,     3,    -5,    -1,    -5,    -1,     1,    -1,     0,    -1,     1,    -2,   -14,   -13,   -13,   -12,    -8,   -10,     0,    -1,   -10,    -4,   -10,   -10,    -4,    -4,    -4,    -4,    -2,     4,    -7,    -5,     1,     2,     2,     1,     3,    -7,    -2,    -3,    -2,     0,    -6,    -6,    -7,     0,     5,    -3,    -7,    -3,    -8,    -6,   -13,    -5,    -7,    -6,    -5,   -11,    -3,    -4,     0,     0,     1,     1,     5,    -4,    -7,    -5,     5,     8,     4,     0,     0,    18,     3,    -7,    -2,    -3,    -9,   -13,    -8,    -3,    -8,     1,    -3,   -13,    -6,    -4,     1,     0,     2,     0,     1,   -10,    -1,    -4,     1,     5,     2,    -1,    -4,    -5,    -3,     6,     4,    -5,    -8,    -7,     1,    -3,   -18,   -11,   -11,   -16,    -1,    -1,     1,     2,     0,     2,     0,    -5,    -5,    -6,    -5,    -7,   -13,   -12,    -4,   -11,    -8,     0,   -14,    -6,     1,     0,    -7,    -6,    -6,    -2,   -12,    -2,     2,     1,     0,     2,     0,    -1,    -1,    -1,     1,    -1,    -2,    -1,    -2,    -5,    -4,    -6,    -6,    -9,    -6,   -12,    -1,     1,     0,    -9,    -5,    -6,    -3,     2,     0,     0,     2,     1),
		    94 => (   -1,    -2,     1,    -1,     1,     2,     0,    -1,     1,     2,     2,    -2,    -4,    -2,    -4,    -3,    -1,    -1,    -1,    -2,     2,     1,     0,     2,    -2,     1,     0,    -2,     2,     2,     0,     2,     1,     0,    -5,   -10,    -2,    -9,    -9,   -10,   -10,    -9,    -2,   -13,   -12,    -6,     0,     0,   -11,    -3,    -4,    -1,    -2,    -1,     0,     1,     1,    -1,     1,   -13,   -20,    -5,   -10,   -14,    -7,   -10,   -17,   -28,   -18,   -12,   -17,    -8,    -2,    -6,   -12,   -12,   -13,    -2,    -9,    -8,   -12,    -6,    -2,     0,    -1,    -2,     0,   -15,   -24,    -5,   -18,   -17,    -9,   -13,   -16,    -8,   -10,   -21,   -14,   -10,     7,    -9,   -14,     0,    -3,     2,     3,     5,   -13,    -9,     1,     2,     2,     1,    -7,   -12,     2,    -7,   -15,     1,     1,    -5,   -15,    -2,     7,    -8,    -7,   -20,    -7,   -11,   -11,    12,     8,     7,    -1,    -7,   -14,     3,    -4,     0,    -1,     0,    -7,   -13,   -14,    -7,   -10,    -1,     5,     3,    14,    -5,    -4,    -8,   -15,   -19,    -7,     3,    24,     5,     2,     4,    -8,    -9,   -14,     6,    -9,     1,     1,     0,    -2,    -3,    -8,    -7,    -2,     1,    -4,    -3,   -17,    -8,    -8,    -2,   -22,   -35,    -6,     2,    10,    14,    21,    20,   -10,    -6,   -10,    -8,    -2,    -7,     2,    -5,   -10,     0,    -8,    -1,    -3,    13,    -3,    -9,   -14,     3,     9,    -6,   -28,   -25,    -3,     5,    10,     7,     6,     6,    -7,    -7,   -15,   -12,    -4,    -7,   -10,   -11,     9,    -1,    -5,     0,     5,     7,    -8,   -13,   -10,     5,     1,   -11,   -17,   -13,   -13,    20,     2,     7,     0,   -12,   -12,   -17,   -14,    -6,   -12,    -6,    -1,   -10,     7,    -5,    -7,    -9,     1,    -2,    -6,    -4,   -15,    -1,    -5,    -4,   -10,   -18,    -1,    12,     6,    -3,     1,    10,     3,   -13,   -12,    -3,    -3,    -5,     0,    -8,     9,    12,    -1,    -8,   -12,     1,     2,    -8,     5,     0,    -4,    -2,   -12,   -25,    -6,     8,     2,    -3,    -6,     8,    -9,   -21,   -18,    -3,    -1,    -4,     1,   -16,    -5,     9,   -11,     0,    -3,    -5,     7,    -1,     5,     8,     3,    -6,   -24,   -18,     1,     9,     1,    -2,    -8,   -18,   -17,   -17,   -26,   -11,    -3,   -11,     2,    -8,     4,    -1,    -9,     0,    11,     4,     1,    -2,    12,     5,     6,   -17,   -18,   -18,     0,     2,     3,    -3,   -11,   -15,   -15,     2,     6,     3,    -7,   -11,     0,    -8,    -3,    -3,    -4,     1,    12,     3,     0,     3,     7,     7,    -4,   -17,   -19,   -15,    -6,     5,     6,    -7,   -12,     3,     9,     8,    -8,    -5,   -12,     2,     1,     1,   -14,    -4,    16,    10,     0,     6,    -4,    13,    16,    11,    -2,    -5,    -5,   -11,    -1,     2,     4,     3,     3,     9,    -1,     2,    -4,   -11,   -10,    -1,     1,    -1,    22,    -1,    13,     4,    -3,    -3,     2,     3,    11,     7,     7,     1,    -8,   -12,    -4,    -1,    -3,     7,    -2,     7,    18,    -5,   -16,   -18,    -7,     2,     0,    -2,     1,   -12,    -7,   -11,     4,     0,    -6,    -2,    -3,   -17,   -10,    -6,   -10,    -4,    -3,     2,     5,    -4,     9,     3,    -1,   -19,    -5,   -10,   -12,    -5,    -2,     2,     5,   -18,     0,    -2,     1,     6,     8,    -3,     0,    -3,   -18,    -3,     1,     7,    -2,     4,     5,    -5,     2,     7,    -9,    -6,   -13,     7,    -2,    -8,    -6,     2,     6,   -10,     4,     7,     5,    10,     0,    -3,    -6,    -7,   -18,    -3,     5,    12,    -2,     5,     3,     5,    10,     2,   -15,    -3,   -12,   -10,    -4,    -2,     1,    -2,   -11,     1,    -3,     2,    11,     0,     2,     2,    -1,   -20,   -20,    -6,    -3,    13,     2,    -8,     9,     6,     6,    10,    -9,    -7,   -12,   -16,     0,    -2,    -1,     1,    -6,    -3,     3,    -6,     1,     4,    -1,    -8,   -14,    -4,    -2,     0,     1,     2,     1,     6,     8,     8,     7,    10,   -11,    -3,    -1,    -6,    -1,     0,    -2,     1,   -13,    -2,     2,    -3,     3,     5,     4,   -12,   -11,   -12,    -2,     0,     0,     3,    -6,     7,     5,     2,     8,     9,     8,    -6,     9,    -2,    -8,    -1,     2,     2,    -1,   -13,   -19,     7,     3,    -3,   -13,   -19,   -29,   -14,    -9,     0,    -2,    -4,    -5,    -9,     3,     7,    10,    12,     3,    -4,    -2,    16,     4,    -1,     0,     0,    -1,    -8,   -13,   -10,    -2,    -5,    -3,   -19,   -25,   -13,   -11,    -8,    -2,     0,     6,   -10,     0,     7,    11,    18,   -10,    -7,     1,     5,     3,    -1,     2,     2,    -1,    -3,    -6,    -2,     0,    -2,    -7,   -12,   -15,   -13,    -7,    -2,   -12,    -7,     1,    -4,     1,    -4,     2,    -3,   -13,    -2,   -11,    -7,    -5,     1,    -1,     2,    -7,    -2,    -7,    -1,    -3,     1,    -5,   -12,   -18,    -7,     1,    -7,   -22,    -1,     3,    -3,   -12,   -23,   -11,   -16,   -19,    -9,   -13,    -9,    -6,     2,     0,    -2,     0,    -2,   -10,     1,    -1,    -3,    -4,   -12,   -21,    -2,    -7,   -14,   -22,   -14,   -23,   -17,   -17,   -16,   -24,   -18,   -20,    -3,    -2,     2,    -1,     1,     2,    -2,     2,     2,    -3,     1,    -3,    -6,    -4,    -7,   -12,   -10,   -10,    -6,    -9,     1,   -13,   -18,   -12,    -9,   -10,    -7,   -11,    -4,     2,     0,     1,    -2),
		    95 => (   -1,     1,     1,    -1,    -1,     1,     2,     0,     2,     2,    -1,    -2,     1,    -1,     0,     0,    -1,    -2,     0,     1,    -1,    -2,    -1,     1,    -2,     2,     1,    -2,     2,     0,    -1,     1,    -1,     2,     0,     2,    -1,     2,    -3,    -2,     0,     1,    -2,    -3,    -5,    -6,    -1,    -1,    -1,    -1,     2,     2,    -1,    -2,     0,     2,    -1,     0,    -1,     2,     2,    -2,    -3,    -5,    -6,   -10,    -9,    -8,   -10,    -7,    -5,     5,    -2,    -2,    -1,     5,     7,     3,     3,    10,    -3,    -2,     0,    -1,     0,     0,    -4,     3,    -1,    -3,   -10,   -14,    -4,     0,    10,     3,    10,    14,    19,     6,    -5,   -10,    14,    -4,    -3,     4,    -5,    -7,    -7,     2,     4,    -1,     1,    -2,    -6,     0,    -7,    -8,     8,    -1,   -14,    11,     0,     8,     9,    -9,   -10,    -4,     3,    -6,     3,    11,    -9,     3,    10,    12,    22,    20,     6,    -6,     1,     2,    -4,     1,     0,     2,    -6,   -11,     1,    15,    15,     1,   -12,   -13,    -8,    -4,     7,     1,     5,     1,     4,    10,    10,    10,    15,    13,    12,    -5,    -1,    -3,    -3,    -3,     6,     4,    -9,    -4,    14,     2,     5,   -13,   -11,    -2,     5,    14,     6,    12,     9,    -4,     4,     7,    14,    -3,     8,     7,    12,     0,     0,     0,     0,    -8,    -1,    -2,    -6,     7,     8,    11,     9,    -1,   -13,    -6,    13,    12,    19,    14,     5,     4,     4,     3,    -4,    -9,    -6,     9,     9,     3,     0,    -2,   -14,   -11,   -12,    -6,     0,     4,    17,    12,    11,    -8,    -5,   -12,    -2,     3,    -5,     2,     4,    -8,    -3,   -13,    -7,    -7,    -7,    -9,    15,     3,    -1,    -3,   -14,   -13,    -7,    -4,     1,     2,     9,     9,     6,     9,   -17,   -22,   -26,   -31,   -34,   -45,   -24,   -33,   -32,   -30,   -20,   -15,   -14,    -9,    15,     7,     2,    -1,    -5,   -10,    -4,    -2,    -6,     1,     7,     7,     3,    -4,   -17,   -21,   -26,   -18,   -18,   -38,   -41,   -36,   -43,   -41,   -38,   -17,   -10,    -5,     5,     9,    -1,    -1,    -1,    -2,    -1,    -5,     0,    -2,     5,     3,    -8,    -3,    -6,    -7,     0,     5,     7,     1,   -10,   -12,   -21,   -23,   -28,   -23,   -17,    -4,     1,     3,     0,    -1,     0,     7,     1,     7,     8,     3,    12,     2,     9,     1,    -5,    -6,    -6,     4,     5,     4,     5,    -5,     1,     2,   -10,    -6,   -11,    -9,    -1,     1,    -1,     2,     0,     4,     9,     4,    -7,    -6,    -3,     5,     1,     6,    -6,    -7,   -10,   -11,    -1,    -1,     3,     2,     1,     1,     2,     8,    -3,    -5,    -7,   -12,     1,    -4,    -3,     1,    13,     5,    11,     0,    -3,     8,     0,    -4,    -4,   -11,    -8,     2,    -2,    -9,    -5,   -10,    -1,    -3,     7,     3,    20,   -10,   -13,    -7,     1,     4,    -3,   -16,   -10,   -14,     6,   -12,     0,    -3,     8,     7,    -5,    -6,    -7,    -8,    -4,   -17,    -9,     1,     2,    -5,    -2,    -2,    17,     0,   -10,   -11,    -3,    -2,    -2,    -9,   -18,   -14,    -8,    -4,    -7,     2,     6,     0,    -3,    -9,    -2,    -3,    -2,    -8,   -17,    -8,    -4,     2,     4,     2,    -1,    -9,   -19,   -17,    -1,    -4,    -7,     9,     0,    -9,     4,     2,    -7,    -3,     2,     1,    -1,    -6,   -12,   -16,    -8,   -10,    -4,     6,     4,     4,     5,     1,     1,    -2,   -18,   -18,    -2,     1,     8,    13,    -6,     4,    -3,    -1,    -2,   -12,     1,    -4,    -9,   -14,   -26,   -14,   -12,   -11,    -3,     1,     0,    10,    -8,    -9,    -2,    -1,   -20,   -17,     2,     0,    14,    13,     6,     1,    -7,   -14,   -21,   -12,    -7,   -16,    -7,   -26,   -13,   -18,   -15,     3,     4,     7,    11,     5,     2,    -7,    13,     1,    -4,   -12,    -1,    -1,     7,    10,     9,    -3,    -9,    -8,    -7,    -2,    -5,    -5,    -5,     3,    -5,     7,     2,     9,     6,     5,     0,     2,     0,    -3,    -6,    -2,   -13,     2,    -2,    -1,    -4,     5,     9,    -1,     2,     1,    -9,   -16,     0,    -4,    -3,     0,    -9,    10,     4,    13,     3,    -4,     0,     6,     8,    12,     4,    13,    -2,     0,    -2,     1,    -9,     4,    -3,     4,     0,    -3,    -4,    -8,   -10,    -3,    -5,    -4,    -8,     9,     9,     2,     2,    -2,     2,     1,     3,    21,     4,    21,    19,    -1,     0,    -2,     7,     7,     0,     1,    -2,    -6,     8,     2,    -5,    -1,    -3,    -1,     3,    -6,    -5,    -5,    -6,    -8,    10,     3,    10,    10,     6,    14,    23,    -2,    -1,    -1,     1,    10,    13,     7,    10,    -6,    -3,     8,    -4,    -9,    -1,     7,     4,    12,   -10,    -2,    -1,     2,     2,     5,    -4,   -14,    -3,    -5,    -3,     1,    -2,     1,     2,    12,   -11,    -6,    15,     8,    14,    16,    11,    -2,    16,    11,    12,     9,    -8,     0,     9,    14,    12,    10,    19,    11,     8,    -2,     1,     0,    -2,    -2,    -1,    -1,    -2,    -4,    -3,    -2,     0,     1,     0,     3,     1,    13,     7,     2,   -20,    -9,    -4,     2,   -12,    -8,     3,    -6,    -4,     2,     2,    -1,     1,    -1,     1,     1,     1,    -2,     0,     1,    -2,     2,     1,    -1,    -1,     1,    -5,    -4,    -2,     0,    -1,    -4,   -10,   -12,   -10,     0,     1,     1,    -1,    -1),
		    96 => (   -1,     1,    -2,     1,    -2,    -1,    -2,    -2,     2,     1,    -2,    -2,    10,    10,    -2,     0,     2,    -2,     0,     2,     1,     0,     1,     1,     1,     2,     1,    -2,     0,     2,     0,     1,     2,     5,     5,    10,    15,     9,     7,     5,    14,    22,    -7,     4,    10,    13,    12,     4,    11,     6,     5,     4,     2,     1,     1,    -2,     0,     1,     1,    -1,    14,    16,    11,    11,     6,     7,    12,    16,    25,    18,     9,     9,    11,    12,     4,     1,     3,    -3,    -3,    -3,     4,     3,     2,     0,    -1,     1,    -2,    20,     0,     2,    17,    21,    11,     8,    12,     2,     6,    19,    13,     8,    -3,   -11,    -8,    -1,     5,    -8,    -4,    -3,    -2,    -3,     0,     2,    -1,     0,    -4,    24,     2,    18,    14,     0,    -1,     3,     3,     3,    10,     2,    -1,    -6,   -10,    -3,    -4,    -6,   -20,   -11,   -15,   -15,   -15,   -11,    -1,     3,     0,     0,    -3,    -4,     7,     5,    -1,    -6,    -8,     2,     4,     1,    12,     1,   -16,    -1,   -17,    -5,    -6,   -13,   -22,   -23,   -26,   -18,   -10,    -7,     4,     4,     2,    -2,    -2,   -12,     6,    -3,    -8,   -16,   -14,    13,     5,     9,     7,     1,    -6,   -18,   -13,   -14,   -29,   -30,   -20,   -30,   -27,   -25,   -13,    -4,     2,    -9,    -1,     0,    -2,   -15,     7,     3,   -13,   -17,    -1,    -1,     7,     6,     3,     1,   -10,   -19,   -27,   -28,   -35,   -24,   -16,    -5,   -28,   -28,   -20,    -8,     4,   -11,    -2,     1,     1,   -13,     9,     0,    -6,    -5,     8,     6,     2,    -1,    -5,     0,   -25,   -40,   -29,   -16,   -17,     0,     1,     6,    -8,   -15,   -20,   -18,     1,   -13,     0,    -3,     0,    -4,    10,    -2,   -10,    -3,     6,    -2,    -3,     4,     0,   -27,   -17,   -13,    -4,    -1,    -2,    14,    16,    13,     8,     4,    -1,   -15,   -11,    -6,    -1,    -3,    -1,    -4,     5,     4,    -7,    -1,     6,    -7,     3,    -3,    -4,   -30,   -19,     1,     4,    13,    11,     6,     7,     5,    -3,    -2,     5,    -6,   -15,   -18,     1,     2,    -3,    -8,     9,     8,   -10,     3,     2,    -5,    -6,    -7,   -12,   -26,   -13,     0,     8,     7,     7,     7,     8,    -1,     0,    -3,     2,     1,    -7,    -9,    -1,     0,    -5,   -14,     3,    -2,    -3,     0,     3,    -3,    -6,    -6,   -14,    -7,     8,    -8,     9,    -4,     7,     9,     9,     5,    10,    10,    11,     5,   -11,   -11,    -1,     0,    -5,   -13,    -4,     9,     4,    -6,     0,    -3,     3,   -13,   -18,    -5,    -1,    -1,     6,    -1,   -12,     7,     1,     7,     7,    16,    12,     4,    -9,     2,     1,    -1,    -3,   -11,    -8,     4,    12,    -4,     9,    -3,     4,     2,    -9,     0,     1,     6,     2,     1,    10,    -8,     5,     3,    11,    13,     3,    22,    -3,     0,    -2,     1,    -4,    -8,   -10,    -3,    10,    -2,     1,     2,     0,    -1,    -3,     8,     7,     3,    -3,    -4,     3,    -7,     4,     7,    -2,    -2,     5,    16,     0,   -14,     1,    -1,    -5,   -11,    -5,     2,     8,     2,    -4,     1,     6,    11,    -6,    -2,     6,     0,     3,    -1,   -13,     4,    -6,    -2,    -7,     3,    11,    16,     0,    -9,    -2,     1,     2,   -10,    -7,    -5,     0,    -2,     7,    -7,     0,    -6,    -4,     3,    10,     7,    -4,    -9,    -8,     0,   -14,    -3,    -6,     1,    17,    15,    -2,    -8,     2,     2,    -1,   -10,     6,    -6,   -13,     6,     0,    -6,   -18,   -11,    -8,     0,     5,    -3,    -3,     1,    -2,    -4,    -2,    -5,     2,     9,     9,     3,    -6,    -5,     1,    -3,    -1,    -4,    10,    -9,    -7,     3,     5,     0,     0,   -13,   -12,    -6,    11,     9,     8,    -4,   -13,    -6,     0,    -3,    -4,     0,     0,     8,    -7,     1,     1,    -2,     1,    -7,    10,     0,   -14,    -4,   -12,    -3,     2,    -9,   -13,    -6,     6,    21,    11,     4,    10,    -6,     7,    -6,   -10,   -11,    -6,     7,     2,     0,     1,    -1,    -2,    -4,     3,    -2,    -1,     5,    -9,    -4,    -6,   -10,   -12,     3,     8,     7,     3,     6,    -8,   -13,     2,    -9,    -5,   -11,   -12,    -2,     3,     1,     2,     1,    -3,    -4,    -4,    -1,     4,   -13,   -23,   -15,   -11,   -18,   -10,     2,    -2,    -8,   -11,    -5,    -9,   -13,    -7,   -19,   -21,   -22,   -22,    -6,     4,     0,     0,    -2,     0,    -3,    -6,    -2,    -2,    -7,   -10,   -19,   -26,   -19,   -15,    -3,    -3,   -17,   -32,   -33,   -28,   -17,    -4,   -15,   -17,   -11,   -19,    -1,    -1,    -2,     2,    -2,    -1,     0,    -2,     0,     0,    -4,    -4,    -1,    -1,     4,     1,    -9,   -14,   -14,   -20,   -10,   -16,   -20,    -6,    -5,    -5,     0,    -2,    -2,     0,     0,     2,     2,    -2,    -1,     1,     0,    -3,    -5,    -5,    -3,    -3,     0,    -2,     0,    -1,    -2,     0,    -1,    -2,    -6,   -14,    -6,    -9,    -8,    -2,     2,    -1,     1,     1,     2,     0,    -1,    -2,     0,     2,    -3,    -2,    -2,    -3,    -7,    -3,    -1,    -5,    -4,    -2,    -3,    -3,     1,    -4,    -1,     1,    -1,     1,     0,    -1,    -2,     1,     0,     1,    -2,    -3,     1,     2,     0,     2,    -2,    -5,    -1,     2,     1,    -1,     0,     0,     0,     1,    -2,    -1,     1,     1,     2,    -2,    -2,     0,    -3),
		    97 => (    0,     1,     2,    -2,     2,    -1,     2,     1,    -2,    -1,     0,     0,     0,     1,    -2,    -1,     2,     2,     1,     2,     1,    -1,    -2,     1,    -2,     1,     0,    -1,     1,     1,     1,     2,    -2,    -2,    -2,     2,    -2,     0,    -2,    -9,    -5,    -6,     2,    -5,   -11,   -16,    -1,    -4,     0,    -1,    -1,     0,    -2,     0,    -1,    -1,     3,    -1,    -2,    -3,    -5,    -1,    -2,    -4,    -2,    -9,   -10,   -20,    -3,    -2,    -4,    -8,    -5,     0,    -1,     0,    -5,    -4,    -6,    -7,    -1,    -1,     0,     0,     0,    -1,     2,    -4,    -1,   -12,   -11,   -25,   -22,   -19,   -22,   -27,   -24,   -27,   -14,    -6,    -6,    -5,     0,    -8,   -11,   -12,   -19,    -5,    -4,    -5,    -1,     1,     1,    -1,    -3,    -4,   -14,   -18,   -20,   -21,   -33,   -35,   -32,   -18,   -18,   -17,   -16,   -11,   -24,   -18,   -13,   -11,   -13,    -7,   -15,   -27,   -27,   -15,    -5,     2,     0,     0,     2,   -17,   -28,     5,   -13,    -4,     3,     6,    -9,    -6,     1,     8,    11,    -2,    10,     4,     0,   -13,   -22,   -14,    -9,   -30,   -21,   -26,   -13,    -1,     0,     0,    10,    10,     8,    -7,    -6,    -6,    -8,     1,    -3,     1,     5,     1,     4,     9,    -3,    -6,    -3,     3,    13,     9,     9,   -11,   -21,   -16,   -15,    -9,    -2,    12,    12,     5,    10,   -11,    -5,     2,    -3,     0,    -4,     3,     6,     3,     5,    -6,    -5,    18,     1,    -4,     1,    -1,    -3,    -4,    -1,   -17,   -22,   -11,   -12,    25,     6,    -2,     6,     0,    -7,     4,     5,    10,     9,     5,     1,    -4,    -7,     0,    -3,     7,    12,     3,     8,     0,    -6,    -7,    -9,   -25,   -29,    -9,     2,    12,    -4,     2,     8,     6,     7,     2,     8,    15,    14,     3,   -11,    -5,     5,     5,     1,     8,     9,    -1,    10,     0,     5,    -6,   -12,    -2,    -1,    26,     1,    10,     7,     0,     7,     7,    -2,     8,    14,     7,     7,    -9,   -16,    -4,     7,    17,     8,     0,     6,     4,    12,     0,    -3,   -10,    -9,     7,     1,    22,    -2,     2,    17,     4,    -5,    -1,    -2,     5,     8,     6,    -8,    -8,     6,    13,    22,    15,    10,     0,     8,    -5,     5,    -7,     0,     6,     4,   -18,   -10,    14,     0,     7,    16,     4,    -8,    -7,    -1,    -1,     6,     2,     4,    13,    10,    11,    22,    20,    13,     7,     1,   -12,    -4,     0,    16,     1,     5,    11,     9,    13,     0,     4,    15,     0,   -13,    -7,     4,    -2,     1,     4,     1,     9,    11,     8,    25,    16,    11,     4,   -10,    -9,   -17,    -6,     2,    -5,     1,    11,    -3,   -10,    -3,     6,     7,   -10,   -16,    -2,    -3,    -9,    -1,     2,    -6,     4,     2,     4,    15,     3,     4,     7,    -5,    -5,    -8,   -15,    -5,     3,    10,   -11,   -13,     0,    -1,     0,     3,   -10,   -13,    -3,     1,    -4,   -17,   -15,    -6,    -4,    -6,     1,    -4,    -7,     0,     6,    15,    -3,     2,     2,    14,     9,     9,     4,    -6,    -8,     1,    -4,    -1,    -8,    -4,    -1,     0,    -2,     0,    10,     7,    -6,   -16,    -9,    -8,    -3,    -5,    17,    27,    21,     6,    17,    11,    16,    12,   -11,   -10,    -9,     1,    -4,    -3,    -5,     0,     2,     0,    -8,    -1,     0,     0,   -11,   -19,    -7,     0,     1,    12,    18,    23,     4,    12,     8,    15,    13,     2,     8,    -3,   -14,     3,     1,     5,    -5,    -1,     9,     9,    -5,    -8,   -11,    -5,    -9,   -10,    -7,    -5,     2,     4,    26,    14,     8,     4,     2,     9,     3,     1,     3,     1,    -9,    -2,     5,     1,    -2,     4,     5,     5,     2,     6,   -10,    -5,    -6,   -10,   -13,    -6,    -7,    14,    27,     9,     9,     1,     5,     2,    -1,     8,    -2,   -10,    -3,     1,     6,    -3,    -6,   -16,     3,     1,     6,     5,     2,    -4,    -4,    -6,     0,     0,     5,     1,     6,    -2,    -1,    -1,    -1,    -7,    -6,     6,    -6,   -11,     1,     0,     1,    -2,    -5,   -11,     9,     8,     9,     6,    11,    10,     1,     3,     3,    -5,     5,     2,    -8,   -13,   -10,    -5,     4,    -5,    -4,   -11,    -9,    -3,     2,    -1,    -1,    -6,   -11,   -12,     6,    16,     7,     1,     2,     5,    -3,     5,     4,    -3,   -11,    -1,   -14,   -10,   -12,   -13,   -10,   -18,   -18,   -11,     2,   -12,    -2,    -2,     2,    -5,   -20,   -10,     8,    14,     9,     5,    -1,    11,    -1,    -4,    -1,   -19,   -16,    -7,   -15,   -18,   -15,   -10,   -10,   -21,   -19,    -7,     2,    -9,     2,     0,     1,     0,    -3,    -1,    11,     5,     9,     0,     1,     0,     3,    -2,     0,   -11,   -14,    -9,    -7,   -21,   -19,   -16,    -4,   -17,   -20,   -11,   -10,    -2,     2,    -1,    -2,    -6,    12,    -1,    -1,     1,     3,    -9,     5,     4,    -2,    -4,     3,   -18,   -16,     1,   -12,   -15,   -21,   -13,    -3,    -1,   -13,    -5,    -3,    -1,    -1,    -2,    -1,    -1,   -13,    -9,   -13,    -7,    -6,     2,    14,    -2,    -4,    -1,    -1,     1,     2,    -3,   -12,    -3,    -3,     0,     6,    -1,     0,    -2,     0,     2,     1,     0,     2,    -2,     0,     5,     7,     0,    -6,    -4,     0,     0,   -10,    -3,    -6,   -11,     3,     1,    14,     6,    -6,     0,     7,    -1,    10,    -2,     0,    -1,    -2),
		    98 => (    2,    -2,    -2,    -1,     1,    -1,     0,     2,     0,    -1,     1,    -1,     1,    -2,     0,    -2,    -2,    -1,     1,     1,     0,    -2,    -1,    -1,     0,     1,     0,     0,     0,     2,     1,     2,    -2,     0,     2,     2,     1,     1,     0,     1,    -2,    -4,    -3,    -9,    -9,    -9,    -3,     2,    -3,    -2,     0,    -2,    -1,    -2,    -1,     1,     1,     3,    -2,    -1,     0,     0,     1,    -1,    -5,   -14,   -19,   -18,    -7,    -1,    -4,   -12,   -12,    -5,    -2,     0,    -3,    -4,    -7,    -5,     0,     0,     0,     0,     2,     2,    -3,    -1,    -3,    -7,    -6,   -24,     8,    12,    15,     6,    15,    17,    11,     6,     1,     5,    -5,   -11,    -9,   -14,    -9,    -1,    -3,    -4,    -3,    -1,     1,    -3,     2,    -3,   -15,   -18,    -4,     4,     5,     7,    -5,   -11,     2,    -4,    -3,    -4,    -2,     1,    -2,     5,     1,     4,   -16,    -9,    -4,    -1,     1,    -4,    -1,    -2,     0,   -13,   -15,   -27,    -8,     5,     7,    -6,    -1,     2,   -14,    -8,     6,    -2,     3,     9,     6,     0,     7,    -1,    -6,   -10,    -8,    -3,     3,    -3,     2,    -1,   -15,    -7,    -6,    -8,     1,    21,    11,     6,     7,     3,     1,     4,     5,     9,     6,     0,    -8,     7,    -6,    -2,    -8,    -3,    -7,    -7,     1,    -1,    -2,    -9,    -5,   -12,    -4,    -1,    12,    17,   -10,    -4,     4,    -8,    -2,    -8,    -6,    -6,    -9,    -2,     0,     4,    -3,   -11,    -6,   -10,    -4,    -5,    -3,    -3,    -3,    -5,   -10,    -6,   -16,   -14,     5,    18,    -6,    -5,    10,     6,    -6,   -12,   -13,    -6,   -19,     2,     0,     3,    -4,    -5,    -2,   -13,     0,     5,     6,    -1,     2,    -1,    -4,    -3,   -19,   -14,    -2,    -5,    -6,     2,    11,    14,     6,    -7,    -9,    -5,    -2,     9,   -11,    -2,     0,     6,    -3,    -6,    -3,     3,   -16,   -15,     1,    -4,    -7,    -8,    -9,   -18,     5,    -8,   -23,    -5,     7,    25,    23,    16,     6,    -2,     1,     3,     3,   -12,    11,     6,     1,   -10,   -17,   -20,   -17,   -16,     0,    -3,    -2,   -11,    -7,    -7,     1,    -2,    -9,    -2,   -18,     1,    12,    19,    14,     0,    -4,   -10,    -4,    -4,    -3,    -3,    -8,    -8,   -19,   -14,    -4,    -6,     1,     1,    -4,    -2,    -4,    -9,    -5,   -13,   -20,   -20,   -24,   -24,     2,     1,     5,    15,     3,    -1,     5,     6,     2,     4,     4,    -2,    -3,   -11,    -7,    -5,    -2,    -1,    -5,    -2,    -6,    -4,    -2,   -11,   -20,   -28,   -21,   -16,   -12,    -1,    -1,    10,     4,    -4,    -2,    -6,   -13,     1,     4,   -14,   -13,   -10,    -9,    -3,    -1,    -2,     0,   -12,    -7,     2,    -1,    -8,   -10,   -14,    -3,     7,     3,     3,    -2,    -8,     0,     1,     0,   -11,    -6,     6,    -4,   -14,   -14,    -8,   -16,    -8,    -2,     2,    -7,    -9,   -11,    -6,    -7,     0,    -4,     3,     0,     5,    -3,   -10,    -6,    -3,     7,    -5,   -10,     1,    -1,     6,   -12,    -9,   -10,    -8,   -18,    -7,     0,    -3,    -5,    -5,    -9,    -1,     9,     7,     2,    12,     2,     1,   -10,    -3,   -16,     0,   -16,    10,    -8,     9,     9,     5,    -6,    -3,    -6,    -5,   -22,    -9,     2,    -1,    -7,   -17,     5,     2,    -5,     9,     8,     2,    -6,    -2,    -4,   -19,   -16,    -4,   -12,    -4,     4,    12,     3,    14,    11,     0,    -9,    -7,    -4,   -10,    -3,    -1,    -3,    -6,    16,     0,     5,    11,    -3,   -10,    -7,     4,    -7,   -17,    -7,    -6,   -22,    -7,     5,     8,     7,     7,     6,     4,   -15,    -8,    -1,    -7,     0,    -5,   -10,    10,    11,    15,    11,     5,   -12,    -6,     1,     4,   -16,   -10,   -11,    -3,    -7,    -1,    -6,     0,     4,     7,     1,    -9,   -13,    -5,   -19,    -6,    -2,    -1,    -8,     2,    10,     5,     8,     5,    -4,   -14,    -3,     3,   -12,    -3,    -2,     3,     7,    -7,    -7,    -5,     8,     6,     3,    -8,    -7,    -1,   -17,    -2,    -6,    -4,    -9,    -9,     2,    -1,     1,    -2,    -7,     0,    -6,    -1,     2,    -6,     7,    -4,    -5,   -10,   -15,     3,     7,     9,    -3,    -7,    -9,    -6,   -14,    -3,    -7,    -5,    -8,   -11,    -9,     1,    14,    10,    -9,    -5,     2,     4,     7,   -10,    -2,   -13,    -8,    -4,    -7,    -4,     2,    -5,   -15,    -5,     1,    -2,    -9,    -1,    -2,     2,    -2,    -4,   -14,     9,     3,    11,     3,    -9,    -5,    -9,     2,    -1,    -1,    -4,    -5,   -11,    -4,    -1,    -7,   -19,    -9,    -4,     1,     7,   -13,    -1,    -2,    -2,    -5,    -4,   -11,   -11,     5,     5,     3,     0,    -9,    -8,    -2,     0,     6,     8,    12,    -7,     1,    -1,    -1,    -7,    -7,    -2,   -11,    -2,    -3,    -1,     1,     2,    -1,    -1,    -3,    -7,     0,    -4,   -11,    -7,   -12,   -13,   -11,   -14,   -14,   -15,   -11,    -7,    -3,    -1,     0,    -6,    -2,    -3,    -3,    -1,    -3,     2,    -1,    -2,    -2,    -5,    -4,    -3,    -2,    -3,    -3,    -4,    -5,    -3,   -10,   -12,   -14,    -8,    -6,    -5,    -5,   -10,   -16,   -16,    -9,     1,     0,    -2,     2,     0,    -2,    -1,     2,     0,    -4,    -3,    -5,    -3,    -3,    -4,    -2,    -2,     0,    -9,    -3,    -2,    -4,    -4,    -4,    -3,     1,    -2,     2,    -1,    -1,    -2,    -2,     1),
		    99 => (    1,     1,    -1,     0,    -2,    -2,    -2,    -2,    -2,    -2,     0,    -1,     1,    -2,     1,     1,     0,    -2,     2,     1,     0,     2,    -1,    -3,    -2,     1,     1,    -1,    -2,     0,    -2,     1,     1,     2,     2,     1,    -1,    -1,    -4,    -5,    -7,    -7,     2,    -2,     1,    -1,    -4,     0,     0,    -1,    -4,    -2,    -1,     0,     1,    -1,     0,     2,    -1,    -2,    -2,     1,    -1,    -2,     0,    -3,     0,    -4,     0,     1,    -5,     1,     1,     1,    -2,     0,    -4,    -4,    -5,    -1,     0,     1,    -2,    -1,     1,     0,     0,    -5,    -2,    -4,    -4,    -3,    -9,    -7,    -4,    -1,     2,    -3,    -3,     1,    -1,    -3,    -4,    -4,    -9,    -2,    -7,    -4,    -8,    -6,    -1,    -2,     0,     0,    -1,    -2,    -3,    -3,   -13,    -1,     1,     1,     0,    -4,   -11,   -10,    -5,   -11,    -6,   -11,    -5,   -14,   -19,    -2,    -2,    -1,     1,   -12,    -4,    -1,     2,     2,    -2,    -5,    -2,     1,    -1,    -3,    -3,    -5,    -3,    -8,   -11,   -14,   -16,   -19,   -12,    -3,    -2,     5,    -7,    -6,    -6,    -3,    -2,    -4,    -5,     2,    -2,     2,    -1,    -6,    -1,    -6,    -8,    -7,   -12,    -4,    -7,     0,    -2,    -1,    -1,     0,    -7,   -13,    -5,    -8,   -10,    -8,    -7,    -5,    -3,     0,    -5,    -7,     1,    -2,    -3,    -5,    -5,    -8,   -15,   -18,   -19,    -9,    -7,     2,     0,     6,     1,     3,     6,    -9,    -4,   -10,    -9,   -16,    -8,     5,    -6,    -2,    -2,    -5,    -9,    -8,    -3,    -5,   -10,   -13,   -15,   -20,   -13,   -10,     0,     3,     3,    -4,     2,     0,     9,    -9,    -3,     3,    -2,     0,    -9,     0,    -1,   -11,    -3,     0,     0,    -9,    -7,    -9,   -12,    -7,   -13,    -4,     2,    -4,     1,     4,     6,     3,     4,    15,     4,    -5,     2,    10,     2,     0,     0,    -2,    -5,    -8,    -5,    -5,    -2,   -11,    -7,     0,    -6,    -9,   -12,    -6,     2,    -8,   -12,     6,     6,     3,    10,     1,     7,    -5,    10,     7,    -3,     1,    -2,    -9,    -9,    -8,    -3,    -7,     0,   -20,    13,     0,    -4,    -5,    -6,    -1,     0,    -5,   -15,     0,     3,     8,     5,    -1,    -7,   -10,    -1,     2,     2,    -3,     0,    -5,   -13,   -12,    -2,    -4,    -1,    -9,     4,    11,     9,     1,     5,     0,    -6,   -20,   -13,    -2,    -4,    -6,     1,    -1,    -3,    -1,    -2,     5,     0,     7,    -1,    -2,   -13,    -6,    -9,    -1,     2,   -10,    -4,     6,     6,     3,     6,    -2,    -7,   -24,    -6,    -3,   -16,   -15,    -9,     2,    -1,    -9,     2,     1,    -5,     9,     3,    -5,   -15,    -9,    -5,     1,    -1,    -7,    -9,     8,     7,     7,    -1,    -2,   -16,   -14,    -5,    -3,   -11,   -11,   -13,    -3,    -4,    -8,     0,     2,     5,     6,    -4,   -11,   -13,    -7,     0,    -1,    -2,     1,   -12,     8,    11,     3,     4,     0,    -9,   -17,    -4,    -8,   -10,    -2,    -1,     1,     0,   -14,     2,    -2,    -3,     4,     5,   -12,   -14,    -8,     0,    -4,     1,    -4,    -7,     8,    14,     9,    17,     6,     2,     3,     2,   -10,     2,     0,     2,     0,   -15,   -10,    -7,   -10,     0,    -2,    10,     7,   -12,    -1,    -7,    -2,     1,    -3,   -19,    -1,    -2,     0,     6,    10,    14,    11,     9,    12,     7,    -2,    -3,    -9,   -11,   -13,    -2,    -7,    -5,    -2,     9,    -3,   -12,    -4,    -8,    -8,    -2,     0,   -19,     5,    -5,    -9,    -2,     4,    -1,    -2,    12,     3,    -1,   -15,    -4,     0,    -5,    -4,    -1,   -13,    -2,    -5,     7,     7,    -6,    -2,   -10,    -5,    -2,    -3,   -11,     8,     0,   -11,   -10,    -6,   -14,   -12,    -5,    -5,     1,   -16,     5,     0,    -7,    -7,    -5,   -16,     0,   -10,    -3,     9,    11,     7,    -9,    -1,    -2,     0,    -4,     8,     6,    -2,    -7,   -10,   -14,    -8,   -11,    -6,   -18,   -13,     5,     5,    -7,   -14,    -5,    -7,     3,     0,    -3,    10,    11,    20,   -10,    -2,     0,     2,    -7,     3,     3,    -2,    -6,    -7,    -8,   -13,    -9,    -3,    -3,    -8,     8,    -6,   -25,    -7,    -3,    -5,    -4,     7,    -8,     1,     5,    12,   -13,    -1,    -1,     2,    -8,    -6,   -11,    -4,    -6,    -9,    -5,    -8,    -5,    -8,    -2,    -2,    12,   -14,   -17,    -2,     0,    -4,     0,     1,    -2,     2,    -4,   -12,    -3,    -1,     0,    -1,    -7,    -6,    -6,    -2,    -3,    -4,    -4,    -2,    -6,    -1,     0,     1,     4,    -7,     2,     5,    -1,    -5,    10,     0,    12,     5,     0,    -5,    -3,    -1,     1,    -2,    -5,    -1,    -9,    -5,     1,     4,    -9,   -10,    -6,    -3,     1,    -3,     3,     4,     8,    -5,    -1,    -1,     9,     5,     7,     5,     1,    -2,    -3,     1,     0,    -2,    13,   -10,     0,     7,     3,     0,   -12,    -5,    -4,     0,    -4,    -9,     8,     6,     4,    -2,    -4,     5,    10,     7,     8,     1,    -4,    -3,    -2,    -2,     0,     1,     2,    15,     8,     6,     7,    -1,     1,     9,    -7,    -2,    -4,   -11,     1,     4,    -1,    -2,    -1,     6,    10,    16,     8,     0,     4,     2,     2,    -1,     0,    -1,    -2,     0,    -5,    -3,     5,    10,     9,     8,     0,     2,    -3,    -8,    -1,    -3,    -3,    -2,    -7,    -4,    -3,    -2,     5,    -6,     2,    -2,     0,     0)
        );

 ---------------------------------INFO-
 -- COEF =21.569042

 -- MIN =-63.999996
 -- MAX =42.39302

 -- SUMMIN =-4547.21
 -- SUMMAX =3306.077
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
