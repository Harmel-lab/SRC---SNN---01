----------------------------------------------------------------------
---
---  producted Package by julia - Weight matrix
---
----------------------------------------------------------------------
---
----------------------------------------------------
---
-- Pascal Harmeling 2025
---
----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package WeightMatrix01 is
	-- Taille de la matrice
    constant ML01X : natural := 100;
    constant ML01Y : natural := 784;

    -- Déclaration de la matrice de poids
	type framebuffer_ML01 is array (0 to ML01X-1, 0 to ML01Y-1) of integer;

    constant ML01 : framebuffer_ML01 :=(
		     0 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,    -1,     1,     2,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     2,     0,    -1,     0,    -1,    -3,     0,    -1,     0,    -2,    -1,    -2,     0,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     1,     0,     1,     1,    -2,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -1,     2,     0,    -2,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,    -3,    -2,    -2,    -3,    -4,     0,     0,    -1,     0,    -2,    -2,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,    -4,    -2,    -3,     0,     2,     0,    -2,     0,    -2,    -3,     0,     0,     0,    -1,    -3,    -1,    -1,    -1,     1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -4,    -3,    -1,     0,    -1,     2,     1,     0,    -2,    -2,    -1,     0,    -3,    -1,    -3,    -1,     2,     0,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -3,    -4,    -4,    -1,     0,     0,     3,     1,    -3,     0,    -2,    -2,     1,    -1,    -2,    -1,    -3,     2,     2,    -3,     2,     1,     0,    -1,    -1,     0,     0,    -2,    -1,    -4,    -1,    -1,     1,    -1,     1,     3,    -1,     1,    -3,    -3,    -1,    -2,    -1,    -3,    -1,    -1,    -1,    -1,     3,     0,     0,     0,    -2,     0,    -1,    -4,    -2,     0,    -1,     1,    -1,    -1,     2,     0,     0,    -2,    -5,     0,     0,    -1,    -1,    -3,     0,     0,    -1,    -1,     1,     1,    -1,    -2,    -1,     1,     0,     0,    -1,    -1,    -1,     0,    -3,    -3,    -1,    -2,     1,    -2,    -2,    -1,    -2,    -2,    -1,    -1,    -2,     0,     0,     3,    -1,     1,    -2,     0,    -1,     0,    -1,    -1,    -2,     0,     1,    -1,    -1,     0,    -2,     1,     4,    -3,    -2,     0,    -2,    -3,    -1,    -2,    -1,     0,     0,     1,     0,     0,     0,     1,     0,     0,    -3,     0,     0,    -1,     1,    -1,    -1,    -3,     0,     2,     3,    -1,     0,     2,     0,    -3,    -2,    -2,    -2,     0,     0,     1,     1,    -1,     0,     0,     1,    -2,    -2,     0,    -1,    -2,     1,    -2,    -6,    -5,     0,     2,     3,     1,     0,     2,    -1,    -2,    -1,    -1,    -2,     0,     0,     0,     0,    -1,    -1,     1,    -1,    -2,    -2,     0,     1,     1,     3,     0,    -4,    -4,     0,     1,     1,     1,    -2,     0,     0,    -1,    -2,     0,    -2,     0,     0,    -1,    -1,    -1,     1,    -2,     0,    -3,    -2,    -3,    -1,     1,     3,     1,    -5,    -2,    -1,     1,     0,    -1,    -2,     2,    -2,    -1,     0,    -1,    -2,     0,     0,     0,    -1,    -2,     0,     0,    -4,    -1,    -2,    -3,    -2,     2,     2,    -2,    -6,     0,    -1,     4,    -1,    -1,    -2,    -2,     0,    -2,    -2,    -1,    -4,     1,     0,     0,    -2,    -1,    -3,    -1,    -2,    -2,    -2,    -5,     1,     1,     2,    -1,    -5,    -2,     0,     2,     1,     0,     1,    -1,    -1,     1,    -1,    -2,    -3,     1,     0,     0,    -1,     1,    -1,    -2,    -1,     0,    -2,    -3,     2,     2,    -2,    -3,    -5,    -1,     0,     0,    -1,     0,     0,     0,     1,    -1,     0,     0,    -2,    -1,     1,     1,     0,     1,     0,    -1,    -1,    -3,    -2,     1,     1,     2,     0,    -3,    -3,     2,     1,    -2,    -1,     0,    -2,    -1,    -1,    -1,     0,    -4,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,    -3,    -3,     1,     0,    -2,    -2,    -1,    -1,     1,     1,    -2,     0,    -3,    -2,    -2,    -1,     0,    -1,    -1,     0,     1,     0,     0,    -1,    -2,    -1,    -1,     0,    -2,    -1,    -1,     1,    -1,     0,    -1,    -1,     1,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,    -2,     0,     1,     1,     0,     0,    -1,    -4,     0,     0,     1,     0,    -1,     1,     0,     1,     0,    -3,     2,     2,     2,    -4,    -2,    -2,    -2,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,    -1,    -3,    -1,     1,    -1,     0,    -1,    -3,     2,     1,     1,     2,    -2,    -2,    -2,    -4,     0,    -3,    -2,    -1,     1,     0,    -1,    -2,    -1,     0,     1,    -1,    -1,     0,    -2,     2,     1,     0,    -3,    -3,    -2,    -2,     0,     3,     1,     1,    -3,    -1,    -1,    -2,    -2,     1,    -1,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,    -4,    -2,    -2,    -2,    -1,    -2,    -3,    -3,    -5,    -4,    -5,    -2,    -1,    -2,    -2,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,     0,     0,    -2,    -1,    -1,    -2,    -1,    -2,    -2,    -1,    -2,    -3,    -1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,     0,     0,    -1,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0),
		     1 => (    0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,     1,     1,     1,     1,    -1,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     2,     2,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,    -2,    -2,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -3,    -4,     0,     1,    -3,    -1,     0,    -1,    -1,     0,     1,     0,    -1,     4,     3,     0,     0,     1,     3,     3,     2,     2,     1,     0,    -5,    -5,    -5,    -4,    -1,    -1,     0,     1,    -2,     1,     0,    -2,     0,     0,     0,     0,     0,     3,     2,     1,    -1,    -1,     0,     0,     0,    -2,    -4,    -4,    -5,     0,     2,     0,     0,     1,     1,     1,     1,    -1,    -5,    -3,    -4,    -3,    -2,     0,    -1,     3,     4,     1,     0,    -1,    -1,    -6,    -3,    -2,    -4,    -5,    -3,     0,     4,     0,     0,     0,     1,     1,    -1,    -2,    -5,    -4,    -3,    -3,    -2,     0,     0,     0,     1,     1,    -1,     0,     1,    -5,     0,     0,    -4,    -4,    -2,    -3,    -1,     0,     1,     0,     1,    -1,    -2,    -1,    -5,    -4,    -1,     0,    -1,     0,     0,    -1,     1,     1,     0,    -1,    -2,    -5,    -1,    -3,    -4,    -3,    -1,     2,     1,     1,     0,     2,    -1,    -2,    -1,     0,    -3,    -4,    -1,    -2,    -1,     0,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -4,    -3,    -2,    -6,    -6,     0,     1,     1,     2,     1,     1,    -1,    -2,    -1,    -2,    -3,    -4,    -2,    -2,     0,     0,     0,    -1,     1,    -1,     0,    -3,    -1,    -1,    -2,    -4,    -8,    -2,     0,    -1,     0,     3,     0,    -3,    -2,    -4,    -1,    -1,    -2,    -3,    -2,     0,    -2,     0,     1,     0,    -1,     0,     0,    -2,    -3,    -2,    -3,     0,    -4,    -3,    -2,     1,     3,     3,     0,    -2,    -2,    -3,    -1,    -1,    -2,    -4,    -4,     0,     4,     0,     0,     1,     1,     1,     0,    -2,    -2,    -3,    -5,    -3,    -4,    -1,    -2,     0,     4,     0,    -3,    -2,    -1,    -1,     1,    -1,    -2,    -4,    -4,     0,     4,     0,     0,    -1,     3,     1,    -1,    -1,    -1,    -5,    -4,    -2,    -2,     0,    -1,     2,     0,     1,    -5,    -5,    -2,     2,     3,     3,     2,    -1,     0,    -1,     2,     0,    -1,     0,     1,     1,    -1,    -1,     0,    -2,    -6,    -3,    -1,    -1,     1,     3,    -1,     1,    -5,    -5,     0,     2,     0,     0,    -4,    -2,     0,     1,     0,     0,     0,     1,     1,     2,    -3,    -2,    -1,    -1,    -4,    -3,     1,     0,    -2,     3,     0,    -2,    -5,     0,     3,     3,     4,     2,    -1,    -2,     4,     4,     0,     0,     0,     1,     4,     1,     0,    -1,     0,     2,     0,    -1,     2,     0,    -1,    -1,    -3,    -2,    -4,    -1,    -3,     0,     4,     2,    -2,    -5,     1,     1,     0,     0,     1,     0,    -2,    -1,     0,     1,     0,     2,     1,     1,     3,     1,     1,    -2,    -1,    -1,    -4,    -4,    -4,     0,     3,     2,     4,     5,    -1,    -1,     0,     0,     0,     1,    -2,     1,     0,     2,     1,     1,     1,     1,     1,     0,     1,     1,    -1,    -2,    -1,     1,     2,     2,     4,     4,     5,     3,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,    -2,    -2,    -1,     1,    -2,     1,    -1,     0,     2,    -2,    -5,    -4,     1,     2,     3,     2,     0,     0,     0,     1,     3,     0,     2,     0,    -1,     2,     2,    -2,     2,     2,     1,     0,    -2,     0,     1,     1,     1,    -3,    -4,    -5,    -1,     2,     0,     0,    -1,    -3,     0,     3,     3,     1,     2,     0,     0,     2,     1,     0,     3,     1,    -2,     0,    -1,    -2,     1,     0,     1,    -2,    -4,    -4,    -1,    -1,     0,     3,    -3,    -2,     0,     1,     1,     1,     0,     3,     2,    -1,     0,     0,    -3,    -4,    -2,     0,    -1,     0,    -1,     1,    -2,     0,    -1,    -4,    -4,    -3,    -1,     2,     1,     1,     1,     2,     2,     0,     0,     2,     2,     0,     0,     0,    -2,    -5,    -1,     0,    -1,     1,    -1,     0,    -1,     2,    -2,    -1,    -3,     0,     2,     4,     1,     2,     2,     2,     3,     5,     1,    -1,    -1,    -1,     0,    -2,     0,    -2,    -2,     2,    -1,    -1,     1,     0,     0,     1,     0,     1,     1,     1,     3,     4,     0,     0,    -1,     2,     3,     5,     0,     0,     0,     0,    -1,    -2,    -3,    -1,    -2,    -1,    -2,    -4,    -1,    -2,    -5,     2,     2,    -1,     1,     1,     6,     4,     1,     0,     1,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     1,    -4,    -2,    -3,    -3,    -3,    -5,    -2,    -3,    -2,    -2,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -1,    -2,    -2,     1,     0,    -3,    -3,    -4,    -4,    -3,    -2,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0),
		     2 => (    0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -3,    -2,    -1,     0,     1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,    -2,    -2,     0,     0,    -3,    -1,    -1,    -1,    -2,    -1,    -6,    -2,     0,    -1,    -1,    -3,    -3,    -2,    -1,    -1,     0,     1,     1,     0,     0,     0,     0,    -1,    -3,    -2,     0,     3,    -1,     0,     3,     3,     0,    -3,    -3,    -2,    -3,    -3,    -1,     2,    -1,    -4,    -2,     0,    -1,    -2,     1,     0,    -1,     0,     1,     0,     1,    -1,    -2,     0,     3,     1,     0,    -3,    -2,    -2,    -4,    -4,    -3,     1,     1,     0,    -1,     1,     2,     0,    -3,     0,     0,    -2,    -1,     0,     0,    -1,     0,     3,     1,     0,     0,    -1,    -1,    -3,    -4,    -4,    -4,    -3,    -2,    -1,     0,     2,     2,     2,     3,     1,    -2,    -2,     0,    -2,     0,     1,     1,     1,     0,     1,    -1,    -1,     2,     1,    -1,    -1,    -2,    -1,    -4,    -3,    -3,    -2,     3,     1,     2,    -1,     1,     0,    -4,    -3,     3,    -2,     0,     0,     0,     3,     0,     0,    -2,     0,     2,     0,     1,     0,     1,     1,     2,    -2,    -2,    -1,    -1,    -3,    -1,     1,     1,     0,    -6,    -1,     4,    -2,     0,    -3,     3,     3,    -2,    -1,     1,     0,    -1,    -2,    -3,     0,     2,     0,     1,     1,    -4,    -5,    -2,    -2,     1,     1,     0,     0,     1,     1,     2,    -3,    -1,     0,    -1,     3,    -2,    -3,    -1,    -1,     0,    -2,    -2,     1,    -1,    -2,     0,     1,     1,    -2,    -1,     0,     3,     1,     1,     1,    -1,    -1,    -3,     2,    -1,    -1,    -1,     3,    -3,    -2,     2,     2,     2,     0,     0,     1,     0,     1,     3,     6,     2,    -2,    -1,     0,     3,     1,     1,     0,    -3,    -1,    -2,     1,    -2,     0,    -2,    -2,    -2,     2,     0,     2,     3,     3,     2,    -2,    -1,    -3,    -1,     0,     0,     0,    -3,     0,     2,     0,     1,     1,    -3,     0,    -1,     1,    -3,     0,     0,    -5,    -1,     3,     2,     2,     2,     0,     1,     0,    -4,    -4,    -2,    -2,    -2,    -2,    -2,    -2,     1,     1,     0,     0,    -4,    -1,     1,     4,     0,     0,     0,     0,     2,    -1,    -2,    -3,    -3,    -6,    -2,    -1,     0,    -2,    -4,    -3,    -3,    -2,     0,     0,    -1,    -1,    -2,    -1,    -1,     2,     2,     6,     1,    -1,     0,    -1,     0,    -3,    -5,    -2,    -2,    -4,    -4,    -3,     1,     1,    -3,    -4,    -2,     1,     1,    -1,    -2,    -4,    -3,     1,     1,     0,     2,     4,     1,     0,    -1,     0,     1,     1,    -1,    -2,    -5,    -2,    -3,     1,     1,     2,     1,     0,     1,    -1,     1,     1,     0,    -1,     0,     0,     1,     1,     1,     2,     2,     0,     0,     0,     1,     2,     1,    -1,     0,    -1,    -1,     1,     1,     1,     0,     3,     3,     3,     4,     0,    -3,    -5,    -3,    -1,    -1,    -1,     1,     3,     2,     0,    -1,     2,     2,     0,     2,     0,    -2,     0,    -1,     2,    -1,     3,     0,     0,     0,     1,    -1,    -2,    -3,    -1,    -1,     0,    -1,     0,     0,     2,     4,     0,     0,    -2,     4,     2,     4,     3,     0,    -2,    -1,     0,    -2,    -1,     1,     1,     2,     1,     0,    -1,    -1,     0,    -1,     0,     0,     4,     1,     3,     6,     0,     0,     0,     4,     5,     2,     2,     1,     0,    -1,     3,     2,     1,    -1,    -1,     1,     2,     1,     0,    -3,    -1,     0,     2,     1,     4,     2,     4,     4,     0,     1,     1,     2,     2,     2,     3,     2,     1,     0,     0,     0,    -2,     0,     0,     2,     2,    -1,    -1,     0,    -1,     0,    -1,     2,     4,     1,     4,    -1,     0,     1,     0,     0,     2,     3,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -5,    -2,     1,     0,     2,     4,     3,     2,    -3,     0,     2,     3,     3,     4,     0,     0,    -1,     2,     1,     3,     0,    -2,    -3,    -2,    -2,    -2,    -3,    -4,    -5,    -2,     0,    -1,     2,     2,     1,    -2,    -1,    -1,     1,     2,    -2,    -2,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,    -2,    -3,    -3,    -4,    -3,    -3,     1,    -4,    -7,    -2,     0,     0,     0,    -2,    -2,    -1,     1,    -1,     0,     1,     1,    -2,     1,    -2,    -2,    -1,    -2,    -1,    -5,    -5,    -4,    -4,    -5,    -2,    -2,    -6,    -8,    -4,     1,     1,     1,    -2,    -1,     2,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -3,    -4,    -3,    -3,    -4,    -4,    -2,    -1,    -4,     1,    -1,    -3,    -3,    -6,    -5,    -3,     0,    -2,    -2,    -1,     0,     1,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -2,    -5,    -3,    -1,    -1,    -2,    -1,    -3,    -3,    -4,    -5,    -5,    -4,    -3,    -3,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -4,    -4,    -1,     0,     0,     0,     0,     0),
		     3 => (    0,    -1,     0,     1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     1,    -1,     1,     0,     1,    -1,    -1,    -1,    -2,    -2,    -1,    -2,    -3,    -2,    -2,    -3,    -4,    -4,    -2,    -5,    -5,    -5,    -2,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -3,    -2,     0,    -1,    -2,    -2,     0,     3,     2,    -1,    -1,    -1,    -4,    -5,    -2,     0,     0,     0,     0,     1,    -1,     1,     3,     1,     0,     2,     2,     3,     3,     0,     0,     1,     2,     0,    -2,    -1,     2,     0,    -1,    -4,    -2,    -8,    -5,     0,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -2,    -3,     1,    -2,     1,     1,     0,     0,     0,     0,     0,     1,     2,     1,     1,     2,     1,    -1,    -2,    -1,    -1,     0,     0,     1,     0,     0,    -2,    -1,     0,     0,     1,     0,     0,     0,     1,     4,     2,     0,     0,     0,     0,     2,    -2,    -1,     0,     0,     0,    -2,    -3,     0,     0,     1,     0,    -2,    -1,     3,     0,     0,     1,     0,     1,     3,     1,    -1,     1,     2,     2,     0,     0,     0,     3,    -1,    -2,    -4,    -2,    -4,    -2,    -1,     0,     0,     1,     4,     2,     1,    -2,     2,    -1,    -3,     2,     1,     3,     1,     0,    -1,    -1,     1,     0,     0,     1,     2,    -1,    -6,    -7,    -2,    -3,    -1,    -1,    -2,     5,     4,     1,    -4,    -1,     0,    -2,    -1,    -3,    -2,    -5,    -6,    -9,    -4,     1,     0,     1,     1,     2,     1,     0,    -4,    -9,    -4,    -4,     0,     0,    -1,     6,     3,    -2,    -5,    -5,    -7,    -6,    -7,    -6,   -11,    -9,    -8,    -3,    -1,     0,    -1,    -1,     0,     1,     2,     1,    -2,    -8,    -2,    -2,    -1,     0,    -1,    -1,    -2,    -3,    -5,    -7,    -5,    -7,   -10,    -7,    -6,    -3,     2,     3,     3,     0,     1,     0,     2,     4,     3,     2,    -5,    -4,    -4,    -2,     0,     0,     0,    -2,    -3,     1,    -1,    -1,    -3,    -1,    -3,    -1,     0,     3,     3,     2,    -1,     0,    -1,     2,    -3,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,    -3,     1,     4,     2,     0,    -2,     0,    -1,     1,     3,     2,     2,    -1,     0,     0,    -2,    -3,    -4,    -3,     0,    -1,     0,    -2,    -3,    -1,    -1,    -1,     1,     0,     0,     1,     3,    -1,    -2,     3,     1,     0,     1,     1,     1,     0,     0,     0,    -1,     0,    -2,    -3,    -1,    -2,    -3,    -4,    -6,    -2,    -1,    -1,     2,     2,    -1,     2,    -1,    -4,    -6,    -3,    -2,     0,     1,     0,     3,     2,    -1,    -1,     0,    -1,     0,    -1,     0,    -3,     0,    -3,    -2,     5,     0,     0,     0,     2,     3,     1,     0,    -7,    -5,    -7,    -4,    -2,     0,    -1,     2,    -1,    -2,     0,     0,     0,     1,     1,     2,    -3,    -2,    -4,    -2,     2,     0,     0,     1,     3,     0,    -3,    -1,    -5,    -2,    -5,   -10,   -12,    -5,    -5,    -5,    -3,    -2,     1,     1,     1,     0,    -1,     1,     0,    -2,    -4,    -4,    -2,    -1,    -1,     1,     4,     1,    -2,     2,     1,     3,     0,    -1,    -4,    -3,    -6,    -6,    -2,     1,    -1,     0,    -1,     1,     2,     2,     0,    -5,    -7,    -3,    -2,    -1,    -1,    -1,    -3,     5,     1,     1,     1,     1,     1,    -1,    -1,    -3,    -2,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -3,    -5,    -2,    -2,    -1,    -1,     0,    -5,     4,     3,     0,     0,     0,     2,     0,     1,     1,     1,     1,    -1,    -2,     0,     0,    -1,    -1,     0,    -2,    -4,    -5,    -4,    -1,    -1,     0,    -1,     1,    -1,     2,     4,     0,    -1,     1,     3,     0,     2,     1,     0,    -2,    -1,    -2,    -3,     1,     0,    -3,    -1,    -1,    -3,    -5,    -4,    -2,     0,     0,     0,    -1,     0,     2,     1,     2,    -1,    -2,    -1,    -2,     0,     0,    -2,    -1,    -2,    -1,    -1,     2,    -3,     0,    -3,    -3,    -5,    -5,    -4,    -2,     0,     0,    -1,     0,     3,     3,     0,     3,    -2,     1,    -2,     0,    -1,     1,    -1,     0,     1,     0,     4,     0,     0,     3,    -2,    -4,    -7,    -5,    -2,    -4,     0,     0,     0,     0,     0,     1,    -1,    -2,     0,    -1,    -1,     1,    -1,    -1,    -1,    -3,    -1,    -2,    -2,    -3,    -1,    -4,    -4,    -3,    -4,    -2,    -2,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,    -2,    -3,    -2,     0,     1,    -3,     0,    -1,    -2,    -5,    -5,    -4,    -2,    -1,     0,    -1,    -4,    -2,     0,    -1,     0,     0,     0,     0,     0,    -2,    -1,     0,    -2,    -3,    -5,    -5,    -2,    -3,     1,     3,     2,     0,    -2,    -3,    -2,    -2,    -3,    -2,    -3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,    -2,     0,    -2,    -2,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0),
		     4 => (    0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -1,    -1,    -2,    -1,    -2,    -4,    -2,    -2,    -2,    -2,    -1,     0,    -2,    -1,    -1,    -2,     0,     0,     1,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -3,    -4,    -2,    -2,    -4,    -3,    -3,    -2,    -2,    -4,    -3,    -3,    -1,    -4,    -3,    -3,    -3,    -1,    -2,     1,     0,     0,     0,     0,    -2,    -5,    -2,    -3,    -2,    -2,    -3,    -1,    -3,    -3,    -3,    -3,    -3,    -4,    -5,    -3,    -1,     0,     0,    -1,    -1,    -3,    -2,     0,     0,     0,     0,    -1,    -4,    -1,     1,     3,     1,    -1,    -4,    -3,    -1,    -1,    -4,    -6,    -5,    -3,    -4,    -2,     5,     2,     1,     3,    -2,    -2,    -1,    -2,     0,     0,     0,    -2,    -2,     0,     1,     3,    -1,    -1,    -1,    -1,    -1,    -1,    -5,    -6,     1,    -3,     1,    -2,     1,     0,     1,     1,    -4,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     3,    -2,     1,     2,     1,    -2,    -4,    -9,    -8,    -4,    -1,     1,     3,     0,     0,     1,    -3,    -4,    -4,    -1,     0,    -2,     0,    -2,    -1,     0,    -1,    -1,     1,     0,     1,     1,     1,     1,    -4,    -7,   -10,    -4,    -2,     5,     3,     3,     1,     0,    -2,    -3,    -3,     0,    -1,    -4,    -2,    -5,     0,     0,     1,     1,     2,    -1,     1,     3,     0,    -1,     0,    -7,    -7,    -3,     4,     3,     2,    -1,    -2,     1,     0,    -1,    -2,     0,    -3,    -5,     0,    -4,     1,     1,     3,     2,    -4,    -1,     2,     0,     2,     2,     3,    -4,    -5,     0,     6,     1,     1,     0,    -3,    -1,    -1,     0,    -4,     1,    -3,    -2,     1,    -2,     0,     2,     1,     0,    -7,    -2,     1,     3,    -1,     1,     3,    -4,    -4,     3,     3,     0,     2,     2,    -2,    -4,    -2,    -5,    -5,     1,     0,    -2,     0,    -3,     1,     1,     2,     0,    -3,    -1,     1,     1,     2,     2,     0,    -6,    -6,     1,     1,     0,     1,    -1,    -4,    -4,    -2,    -3,    -1,     1,    -1,    -4,     0,    -2,     1,     2,     2,     2,     0,     0,    -2,    -2,     1,     0,     1,    -2,    -4,     2,     0,     0,     0,     1,    -2,     0,     2,     5,     5,     4,    -4,    -3,     0,    -1,    -2,     0,     3,     1,    -1,     0,    -1,     1,     3,     0,     0,     0,    -1,    -2,     1,     0,     2,     0,     1,     3,     5,     2,     1,     0,    -4,     0,     0,     0,    -2,     0,     1,     4,     1,     3,     1,     0,     0,    -1,    -1,    -1,    -3,     0,    -1,     1,     1,     2,     0,     4,     3,    -1,     2,    -1,    -2,     0,     0,     1,     1,    -1,     3,     0,     0,     3,     0,     0,     0,     1,     0,     2,     2,     2,     2,     1,     1,     2,     0,    -1,     1,    -2,    -3,    -3,     1,    -1,    -1,     0,    -4,     2,     3,    -2,    -2,     3,     0,    -1,     0,     0,     0,     1,     2,     2,     0,    -1,     2,     0,     0,     1,    -2,    -3,     0,    -1,    -1,     0,     0,     0,     3,     2,     5,     0,    -3,     1,    -2,     0,    -3,    -2,    -1,    -1,     1,    -2,    -3,    -3,     0,    -5,    -2,     1,    -1,    -2,     0,    -1,     0,     0,    -2,     0,     2,     3,     4,    -2,    -3,    -3,    -2,    -1,    -2,    -3,    -2,    -1,    -1,    -5,    -3,    -2,    -3,    -3,    -1,     0,     1,    -1,    -1,    -2,     1,     0,     0,     0,    -1,     1,     0,    -4,    -1,    -4,    -2,    -1,    -1,     0,    -2,     0,     1,     0,    -3,     1,    -2,    -1,    -1,     3,     1,     0,    -2,    -2,    -1,     0,     0,     0,    -1,    -3,    -6,    -4,    -3,    -1,    -3,    -3,    -2,     3,     1,     0,     1,     0,    -1,    -1,     2,     0,    -2,    -1,     0,    -1,     0,    -5,    -1,    -1,    -2,    -2,    -1,    -3,    -2,    -4,    -3,    -3,    -1,    -3,    -1,     0,     0,    -1,     1,    -3,     1,    -2,    -1,    -2,    -3,    -4,    -1,     1,     0,    -4,    -2,     0,    -1,    -2,    -1,    -2,    -1,     0,     0,    -3,     1,    -4,    -3,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,    -3,    -2,    -3,     1,     2,     0,     0,     1,     0,     0,    -1,    -1,    -2,     0,    -1,     2,     2,     0,    -5,    -1,    -2,    -2,    -2,    -1,    -2,     0,     0,     2,    -2,    -3,    -1,    -1,     1,    -2,     1,     0,     0,     0,     1,     0,     0,    -4,    -1,    -2,    -1,     0,    -1,    -2,    -1,    -2,    -2,     4,    -1,     2,     2,     3,    -3,     0,     0,     0,     0,    -4,     0,    -1,     0,     0,     0,     0,    -1,     0,    -3,    -7,    -4,    -3,    -2,    -3,    -3,    -3,     0,     1,    -2,     0,     1,     0,    -2,     0,     2,    -2,     1,    -2,    -1,    -1,     1,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,     1,    -1,    -4,    -6,    -6,    -4,    -2,    -3,    -6,    -1,    -3,    -4,    -6,    -5,    -4,    -1,    -2,     0,     1,     0,     1,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -2,    -2,    -4,    -2,    -2,    -5,    -1,    -2,    -3,    -2,    -3,    -4,    -3,    -3,    -1,     0,     0,     0,     1),
		     5 => (    0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     1,     0,     1,     1,     0,     1,     0,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -2,    -4,    -4,    -6,    -2,     2,     2,     2,     3,     3,     4,     3,     3,     3,    -1,    -1,     0,    -1,     0,     0,     0,     1,     2,    -1,    -1,    -1,    -1,    -3,    -4,    -3,    -1,    -3,     2,    -1,    -4,    -3,     0,    -1,     1,     2,    -1,    -1,     2,     1,     2,     1,     0,    -1,    -1,     0,    -3,    -3,    -4,    -5,    -7,    -2,    -5,    -3,    -3,     0,     3,     0,     1,     0,     0,     0,     1,     2,     2,     3,     3,     7,     2,    -1,     0,     0,    -1,     0,    -3,    -3,    -6,    -6,    -7,    -4,    -1,     0,     1,     0,     0,    -1,     1,     3,     1,     0,     5,     4,     2,     4,     4,     6,     3,    -1,     0,     0,     1,    -1,    -3,    -5,    -5,    -3,    -2,    -3,    -1,     1,     3,     0,     0,     0,     1,     2,     5,     1,     4,     0,     0,     4,     1,     3,     2,     1,     0,     1,     0,    -2,    -3,    -3,    -2,     0,    -1,     0,     0,     3,     2,     1,    -1,    -2,     1,     2,     2,     0,     2,     0,    -2,     0,    -1,     1,     2,     1,    -1,    -1,    -2,    -2,    -2,    -1,    -3,    -1,    -2,    -3,     1,     3,     2,    -2,    -2,    -4,    -8,    -4,    -4,   -10,    -5,    -6,    -4,    -1,    -1,     0,     1,     0,     0,    -1,    -4,    -4,    -4,    -1,    -4,    -4,    -4,    -2,    -2,    -1,    -1,    -2,    -4,   -10,   -12,   -14,   -15,   -14,   -10,    -8,    -7,    -4,    -2,    -2,     0,     1,     0,    -1,     0,    -2,     0,    -1,    -2,    -1,     0,    -2,    -2,     0,    -2,     0,    -3,    -1,     0,    -3,    -9,    -9,    -9,    -7,    -7,    -5,    -3,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -3,    -3,    -2,    -2,    -2,    -1,    -1,     0,    -1,    -1,     1,     0,     1,    -1,    -4,    -7,    -5,    -2,    -3,     0,     1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -2,    -1,     1,     1,     1,     1,     0,     1,    -1,    -1,     0,    -1,    -2,    -4,    -3,    -1,    -1,     0,    -2,     0,     0,     0,    -1,     0,     1,    -2,     0,    -3,     1,     2,     4,     1,    -1,     1,     0,     0,    -1,    -2,     1,     0,     1,    -2,    -1,    -2,     0,     0,    -1,     1,    -1,     0,     0,     2,    -2,    -4,    -3,    -1,    -1,     2,     0,     0,    -1,     1,    -2,     2,     0,     0,    -2,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -2,    -1,    -1,     2,    -2,    -4,    -3,    -3,    -2,    -2,    -1,     1,    -2,    -3,    -1,    -2,     1,    -1,    -1,    -2,     1,     0,     1,     1,    -1,    -1,     0,     0,     0,    -2,     1,     0,    -3,    -3,    -5,    -5,    -8,    -6,    -4,     1,     1,    -2,     1,     1,     4,    -1,     1,     1,     1,     1,    -2,    -3,    -2,    -2,    -2,     0,    -1,    -3,     1,    -2,    -2,    -2,    -5,    -2,    -6,    -9,    -3,    -4,    -5,    -4,     1,    -1,    -2,     4,     2,     2,     1,    -1,    -1,    -4,    -2,    -1,    -1,     0,    -1,     0,     2,     0,    -2,    -3,    -1,     2,    -1,     0,    -2,    -6,    -3,     0,    -2,     1,     0,     2,    -1,     0,     1,     0,    -1,    -4,     0,    -3,    -2,     0,     0,     3,     0,     0,    -2,     0,    -1,     1,     2,     1,     2,     1,     1,     1,    -1,     1,     0,     1,     1,     1,    -1,     0,    -2,    -3,     0,    -1,    -1,     0,     0,     2,     1,     6,     0,     1,     0,     3,     2,     0,     1,    -2,     3,     2,     1,     0,     0,    -1,     2,     1,    -2,     2,    -4,    -2,    -2,    -1,     0,     0,    -1,    -2,    -1,     4,     3,     0,    -1,     1,     0,     1,     2,     1,     1,    -1,     1,     1,    -1,    -2,     1,     2,     3,     2,     0,    -1,    -2,     0,     0,     0,     0,    -2,     1,    -2,    -1,    -2,    -1,    -1,    -1,     3,     1,     2,    -1,     0,    -1,     0,    -1,     1,     0,     3,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,     1,     2,    -2,    -2,     1,     0,     3,     2,     1,    -3,    -1,    -1,     0,     3,    -1,    -4,    -3,    -2,    -3,    -2,     0,     1,    -5,    -5,     1,     0,    -1,     0,    -2,     0,     3,     2,     7,     3,    -1,     2,     4,     0,     1,     1,     2,    -2,    -3,    -2,    -3,    -3,    -1,     2,     2,     0,     0,    -1,    -2,     0,     0,     0,     0,     3,    -1,     0,     2,     3,     1,     3,     2,     2,     1,     0,    -2,    -1,    -1,    -3,     1,     2,     0,     1,     2,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,     0,    -1,     1,     1,     1,    -1,    -1,    -1,     0,    -1,    -1,     0,     1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     1,     0,     0,     1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     0),
		     6 => (    0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     1,     1,     2,     3,     3,     1,     3,     2,    -1,     0,     1,     3,     0,     2,     2,     2,     2,     2,     1,     0,     0,     0,     0,     0,     1,     2,     3,     2,     2,     2,     0,     0,    -2,     2,     4,     2,     2,     4,     2,     1,     2,    -1,    -1,     0,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     5,     3,    -1,     3,     4,    -1,     1,    -2,     1,     1,     2,     1,    -1,    -1,     0,    -2,     0,     2,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -2,     3,     0,     1,     2,    -1,     0,     0,     1,     2,    -2,     0,     0,    -3,    -2,    -2,    -2,     3,     3,     1,    -2,    -3,    -2,    -2,     0,     1,     0,     0,     0,    -1,     0,    -4,    -3,    -1,    -2,     2,     0,    -2,     1,     2,    -1,    -1,    -3,     1,     1,     2,     1,     0,    -2,    -3,    -2,    -1,     1,     1,     0,    -1,     1,    -3,    -3,    -5,    -4,    -1,    -2,     0,    -3,     2,     3,     0,     0,    -1,    -1,    -2,     1,     0,    -3,     0,    -3,    -4,    -1,    -1,     2,    -1,     0,    -1,     0,    -3,    -2,    -6,    -4,    -2,    -1,    -1,     1,     4,     3,     0,     2,    -2,    -2,    -2,    -6,    -5,    -5,    -3,    -4,    -5,    -3,    -2,     1,    -3,     0,     0,     1,    -3,    -2,    -7,    -1,    -1,    -3,     2,     1,    -1,     3,     0,    -2,    -4,    -4,    -7,    -6,    -6,    -4,    -5,    -8,    -6,    -5,    -4,    -1,    -3,     0,     0,    -1,    -2,    -1,    -7,     0,     0,    -1,    -2,    -2,     0,    -1,    -3,    -3,    -5,    -5,    -7,    -7,    -6,    -4,    -7,    -6,    -5,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -2,    -3,    -6,    -4,     0,     2,     0,    -2,     0,     1,    -2,    -6,    -6,    -1,     2,     0,    -3,    -2,    -2,    -3,    -1,    -1,     2,    -2,    -3,     0,     0,     0,    -4,    -3,    -1,    -3,     0,     2,    -1,     0,     1,     1,    -5,    -5,    -1,     1,     2,     2,    -2,     0,    -4,    -2,    -3,    -3,     0,    -4,    -2,     0,    -1,     1,    -2,    -3,    -3,    -1,     2,     2,     0,    -2,     0,    -2,    -7,    -2,     0,     3,     1,     0,     2,     2,     0,    -1,    -2,     3,    -1,    -2,    -2,     0,     0,    -2,    -1,    -4,    -4,     0,     3,     2,    -4,    -3,     0,    -1,    -3,    -2,     0,    -1,    -1,     0,     3,     4,     2,    -1,     1,     1,    -1,    -2,     2,     0,     0,     0,    -3,    -5,    -2,     3,     2,     1,    -1,     1,     3,    -1,    -1,     1,    -1,     1,    -2,     2,     2,     1,     2,     3,     1,    -1,     0,    -1,     0,     0,     0,    -1,    -3,    -4,     0,     4,     2,    -1,     0,    -1,     4,     0,    -2,     3,    -1,     0,    -1,     1,     0,     0,     2,     3,     1,     0,     1,    -3,    -4,    -1,    -1,    -1,    -2,    -1,     2,     4,    -1,    -1,    -3,     2,     3,    -1,    -2,     3,    -1,    -1,     0,    -1,    -1,     1,     3,     2,     0,     1,     0,    -4,    -3,     1,     0,     0,    -1,     0,    -1,     2,     1,    -2,    -2,     0,     1,     1,    -1,     0,     0,    -1,    -2,     1,    -1,    -2,     2,     3,     0,     3,     3,    -2,    -3,     0,     0,     1,    -2,     0,    -1,     1,     2,     0,    -3,     0,     0,     2,     1,     2,    -3,    -1,    -2,    -1,     1,    -1,     3,     1,     2,     2,     4,    -2,    -3,     0,     0,     0,    -2,     2,    -3,    -3,     1,     0,    -2,    -2,     0,     2,     2,     3,     2,     0,     0,    -2,     1,    -2,    -1,    -3,     2,     1,     3,    -1,     0,     0,    -1,     0,    -2,     1,    -2,    -3,     0,    -4,    -1,    -1,     0,    -1,     0,     3,     4,     1,     0,     3,    -1,    -1,    -1,     1,     2,     3,     3,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -3,    -4,    -1,    -3,    -4,    -3,     2,     2,    -1,     1,     0,     1,     2,    -2,     2,     3,     1,     1,     1,     0,     1,     0,     0,    -1,    -1,    -1,     2,    -4,    -7,    -7,    -1,    -2,    -2,    -2,    -3,    -1,    -4,    -3,     1,    -3,    -3,    -3,     1,    -1,    -6,    -4,     1,     0,     0,     0,    -1,     0,    -2,     0,    -2,    -2,    -3,    -1,     4,     1,    -6,    -4,    -5,    -5,    -5,    -7,    -6,    -1,    -2,    -4,    -3,    -5,    -5,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -2,     0,    -1,    -3,    -5,    -4,    -2,    -3,    -4,    -6,    -3,    -3,    -1,    -2,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     1,     2,     0,     0,     0,     0,    -1,     0,    -2,    -3,    -2,    -2,    -3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0),
		     7 => (    0,     0,     0,     0,     1,    -1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -3,    -3,    -2,    -1,     0,     1,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -3,    -5,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -2,    -3,    -2,    -3,     0,    -1,    -2,    -4,    -4,    -2,    -2,    -2,    -1,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -4,    -5,    -2,    -5,    -1,     1,     0,    -3,    -4,    -5,    -5,    -4,    -3,    -2,    -2,    -3,    -5,    -3,    -3,    -2,     0,     0,     0,     0,    -4,    -1,     3,     4,     2,     4,     1,    -2,     1,     1,     1,     2,     1,     1,    -1,    -3,    -4,    -6,    -4,    -4,    -6,    -8,    -6,    -2,     1,    -1,     0,    -1,    -3,     0,     2,     2,     2,     1,     0,     2,     0,     3,     1,     1,    -2,    -2,    -2,    -3,     0,     0,    -1,    -3,    -3,    -6,    -3,    -4,    -1,     0,     2,     0,     1,     1,     2,     1,     0,     0,    -2,     0,    -2,     1,    -1,    -2,    -4,    -2,    -2,    -3,    -3,    -1,    -3,     1,     1,    -1,    -4,    -4,    -1,    -2,     4,     2,     0,     3,     4,     0,     2,     1,     1,     1,    -2,    -1,    -1,    -1,     1,     1,     1,     0,     0,     0,     0,     0,    -2,     0,    -5,    -5,    -2,     0,     3,     1,     2,     3,     4,     1,     1,     4,     1,    -2,    -3,    -2,     0,     0,     1,    -1,     0,     1,    -1,     1,     1,     2,    -1,    -2,     0,     4,     5,     0,     0,     0,    -1,     1,    -1,     2,     3,     2,     0,     0,     1,    -2,     0,    -1,    -1,    -1,     2,     2,     1,     2,     1,     1,    -1,     0,     2,     2,     4,     0,    -2,     1,     3,     0,    -1,     3,     5,     3,     2,     0,     0,     0,     1,     1,     0,    -2,     3,    -2,     3,     1,    -1,    -2,    -2,    -1,    -4,    -1,     3,     0,     1,     1,    -2,    -3,    -5,     0,     0,     1,     0,    -2,    -2,    -2,    -4,    -2,    -1,    -1,    -3,     0,     0,     0,    -1,    -2,    -1,    -1,     1,     3,     4,    -1,     1,     3,    -3,    -3,    -4,    -1,    -1,    -3,    -4,    -4,    -4,    -6,    -6,    -1,    -1,     0,    -1,     2,     1,     2,    -1,     1,     4,     2,     2,    -3,    -3,    -1,    -1,    -1,    -3,    -2,    -4,    -3,    -4,    -7,    -5,    -5,    -5,    -6,    -3,     1,     0,     1,     0,     1,     2,     3,    -2,     1,    -1,    -2,    -5,    -3,    -1,     0,     0,    -1,     0,    -5,    -2,    -2,    -6,    -3,    -2,     0,    -1,     1,     0,     2,     2,    -1,     1,     1,    -1,     3,     0,     2,    -1,    -1,    -6,    -2,    -1,     0,    -1,    -1,    -1,    -3,    -3,    -3,    -4,     0,     2,     2,     2,     2,     1,     2,    -2,    -2,     0,    -1,     1,     0,     1,     2,    -2,    -6,    -6,    -3,    -2,     0,    -1,     0,    -2,    -2,    -2,    -4,    -4,     0,     1,    -3,     0,     0,     1,     1,    -2,    -1,    -3,     1,     1,     1,    -1,     1,    -2,    -3,     0,    -1,    -1,     1,    -1,     3,    -2,    -3,    -5,    -5,    -3,    -2,    -6,    -4,    -1,     3,     3,    -3,    -3,    -2,    -1,    -1,    -3,    -2,    -3,    -1,    -3,    -2,    -1,     2,    -1,     0,     1,     0,    -1,    -2,    -6,    -3,    -4,    -3,     1,    -2,    -2,     0,    -1,    -2,    -2,    -1,    -3,    -2,    -1,    -2,    -3,    -2,    -3,    -5,    -1,    -3,     0,     0,    -1,     0,    -1,    -3,    -1,     0,     2,    -1,    -1,    -1,     0,     1,     1,    -3,    -3,    -3,    -4,    -4,    -3,    -1,     0,     1,     0,    -2,    -1,    -4,     0,    -1,    -1,     0,    -3,    -2,     3,     3,    -2,     1,     0,    -1,    -2,    -1,     1,    -6,    -4,    -5,    -6,    -3,    -4,    -3,     0,    -1,    -3,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -5,     2,     3,     3,     3,     4,     1,     1,     0,    -1,    -2,    -4,    -4,    -4,    -3,    -4,    -3,    -3,     0,     1,    -6,    -3,     0,    -1,     0,     0,     0,    -2,    -6,     2,     0,     2,     5,     0,     0,    -1,     1,    -2,    -1,    -4,    -2,    -4,    -7,    -6,    -5,    -5,     0,     0,    -3,    -2,     0,    -3,     0,    -1,     0,     1,     0,     3,     4,     3,     1,     3,     1,    -1,     1,    -1,     1,    -2,    -2,    -6,    -6,    -5,    -3,    -4,     0,    -1,    -5,    -1,    -2,     0,     1,    -1,     0,    -1,     2,    -3,     0,     0,     1,    -1,    -3,     0,     2,    -1,    -3,    -4,    -3,    -4,    -2,    -1,    -2,    -6,     0,    -1,    -4,     1,     0,    -1,    -1,     1,     0,     0,    -3,    -3,    -4,    -1,     2,     3,     1,    -2,     0,     1,     2,    -2,    -1,     0,    -1,     1,     0,    -2,     2,     2,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,     3,     2,    -1,     0,    -1,     0,     2,     1,    -1,     4,     2,     0,     1,     0,     1,    -1,     1,     3,     2,     3,     0,     0,     0,     0),
		     8 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,    -1,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,    -2,    -5,    -4,    -1,    -1,    -1,    -2,    -3,     2,     3,     1,    -2,    -2,    -2,    -2,    -1,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -4,     2,     2,    -1,    -3,    -3,    -2,    -2,     1,     1,     0,     4,     2,     0,    -1,     3,     4,     0,    -1,    -1,     1,     0,     0,    -1,    -2,    -3,    -5,     0,     2,     0,    -3,    -2,     1,    -1,     0,     1,     1,     1,     0,    -1,     0,    -1,     0,     1,    -2,    -3,     2,     2,     0,     0,     0,    -1,    -2,    -2,    -3,     0,     0,    -3,    -2,    -1,     0,     0,     1,     0,     1,    -1,    -3,    -4,     2,     0,     2,     0,    -1,    -1,     0,    -1,    -1,     0,     0,    -2,    -4,    -3,     0,    -1,    -2,    -3,    -1,     1,    -1,    -1,    -1,    -3,     0,    -2,    -2,    -2,     1,     0,    -1,    -1,    -3,    -2,    -2,     0,     0,     0,    -3,    -1,    -1,     0,     0,    -1,    -1,     0,     0,    -2,    -1,    -2,    -3,    -2,     1,    -1,    -2,    -2,     0,     0,    -1,    -2,    -2,    -2,     0,     1,     2,    -1,    -2,    -1,     0,    -1,     0,    -2,    -1,     0,     1,    -3,    -2,    -2,     0,    -1,    -1,    -2,    -3,    -2,     0,     1,     1,    -3,    -4,    -1,     0,     4,     2,     0,    -1,    -2,     0,    -1,    -1,    -2,     1,     0,    -1,    -3,     0,    -1,    -2,    -3,    -3,    -1,    -1,    -3,     1,     1,    -3,    -4,    -3,    -3,     0,     1,    -2,     1,    -1,    -2,     0,    -1,     1,    -2,    -2,     0,     0,     1,     4,    -1,    -2,     1,     0,     0,     0,     1,     2,     0,    -1,    -3,    -4,    -2,    -2,     1,     1,     0,    -1,    -1,    -2,    -1,     2,     1,     0,     1,     2,     1,     0,    -2,    -3,    -1,    -1,     1,    -1,     0,    -2,    -3,     3,    -2,    -2,    -1,    -5,     0,    -2,     0,     0,    -2,     0,     2,     2,     2,     0,     1,     2,     2,    -2,    -1,    -3,    -2,    -3,    -2,    -1,     0,    -3,     0,     1,     1,     2,     1,    -4,    -4,    -3,     1,     0,    -2,    -4,     0,     1,    -1,    -3,     2,     5,     2,     1,    -1,    -2,    -2,     0,     0,    -4,    -1,     0,     1,     3,     2,     2,     0,    -4,    -6,     1,     0,     0,     0,    -4,    -2,    -1,    -1,    -4,     1,     1,     0,     0,     1,     0,    -2,    -1,    -5,    -2,     2,     3,     3,     2,    -1,    -3,    -5,    -4,    -6,     0,    -1,     0,    -1,     1,     1,    -2,    -2,    -2,     0,     0,     1,     2,     0,     0,    -2,    -4,    -2,    -1,    -2,     1,    -1,    -3,    -4,    -2,    -1,     0,    -3,    -2,     0,     0,    -1,     2,     0,    -2,    -2,    -2,    -5,    -3,    -1,     1,     2,    -2,    -1,    -1,     0,    -1,     0,    -2,     0,     1,    -2,    -1,     0,    -1,    -3,    -2,     0,     0,    -1,     2,    -2,    -2,    -3,    -2,    -4,    -8,    -3,     1,     2,     0,     0,     0,     0,    -1,    -3,    -3,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -2,    -2,    -1,    -3,     0,     0,     1,     1,    -1,     2,     1,    -1,    -1,    -1,     0,    -2,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -3,    -4,     1,     1,     0,    -1,     2,     1,    -1,     2,    -2,     0,     0,     0,    -2,    -2,    -2,    -1,     0,     0,    -2,    -2,     1,     0,    -1,     0,    -1,    -1,    -4,    -4,    -1,     1,    -1,    -1,    -1,     1,    -2,     0,    -3,    -3,    -1,     0,    -4,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -2,    -2,    -3,    -1,    -2,    -2,    -1,     1,     3,     1,     1,     1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -4,    -4,    -2,    -2,    -2,    -4,    -2,     2,     1,     1,    -2,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,    -2,     0,     0,    -2,    -4,    -5,    -2,     0,    -2,     0,    -2,    -1,    -3,    -1,     0,    -2,    -1,     0,     1,     1,     0,    -1,     0,     0,    -2,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -4,    -1,    -2,    -2,    -1,     2,     1,    -1,     2,     1,     0,     0,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,    -2,    -2,    -2,    -3,    -1,     1,    -1,     1,     0,     0,     1,     1,     0,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,    -2,    -4,    -5,    -4,    -4,    -6,     0,     0,    -1,    -5,    -4,    -2,    -2,     1,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0),
		     9 => (    0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     1,     0,     1,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -2,     0,    -1,     0,    -1,     0,    -2,     1,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -2,    -1,    -1,    -3,    -2,    -1,    -1,    -2,    -2,    -1,     2,    -1,    -2,    -2,    -2,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -3,    -1,    -1,     0,    -1,    -1,    -4,    -5,    -6,    -5,    -3,     0,     2,    -3,    -4,    -3,    -2,    -2,    -2,    -4,    -3,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -4,    -2,    -3,    -1,    -1,     1,    -1,    -2,    -4,    -5,    -4,    -4,     1,    -2,    -3,    -3,    -2,    -2,    -4,     0,    -1,    -1,     0,    -1,     1,    -2,    -1,    -4,    -3,    -3,    -4,    -1,    -2,    -3,    -1,    -1,    -1,    -3,     0,    -2,     1,     2,     0,    -1,    -2,    -2,    -3,    -2,     0,    -1,    -1,    -1,    -2,    -3,    -4,    -4,    -5,    -7,    -6,    -4,    -2,    -2,    -2,    -4,     1,     1,     0,    -1,     5,     2,     2,     1,    -1,    -3,    -1,    -2,    -2,    -1,     1,     0,    -2,    -2,    -2,    -3,    -4,    -5,    -2,    -4,    -2,    -1,    -3,    -1,     0,     2,     2,     0,     0,     0,     0,     2,     1,    -2,    -2,    -1,     0,    -1,     3,     0,    -1,    -2,    -1,    -1,    -4,    -1,    -1,    -1,    -2,    -3,     1,     3,     0,     0,    -1,     2,    -2,     0,     1,     0,     2,     2,    -5,    -2,     0,    -1,    -2,    -2,     0,    -1,    -3,    -4,    -1,     0,    -1,     1,    -2,     1,    -1,    -2,    -2,    -2,    -5,    -4,    -2,    -1,    -2,     0,     3,     6,    -2,    -4,     1,    -5,    -1,    -1,    -1,    -2,    -2,    -1,     3,     2,     2,    -1,     1,    -1,    -3,    -4,    -5,    -6,    -3,    -1,     2,    -1,     1,     1,     4,     6,     0,    -3,     0,    -1,     0,    -3,     1,    -1,    -3,     0,     1,     1,     2,    -1,    -3,    -2,    -4,    -3,    -1,    -4,     0,     0,     3,    -1,     2,     2,    -1,    -4,    -4,    -4,     0,    -1,    -1,    -2,     1,    -2,     0,     1,     0,     1,     3,     0,     0,     1,    -2,     2,     3,     0,     0,     3,     1,     4,     1,    -1,    -3,    -2,    -2,     0,     0,    -1,     0,    -2,     2,    -2,     0,    -1,     3,     3,     3,     0,     1,     2,     1,     2,     0,     0,     0,     2,    -1,    -4,    -1,    -4,    -4,    -1,     1,     0,     0,     0,    -4,    -2,     2,    -2,    -3,    -2,     1,    -2,     0,     2,     2,     3,     0,     1,     0,     0,     2,     1,    -3,    -4,    -5,    -4,    -3,    -1,     3,    -1,    -1,    -1,    -2,    -2,     1,    -1,     0,     0,    -2,    -1,     1,     1,    -1,     1,    -2,    -3,     0,     1,     1,     0,    -4,    -1,    -1,    -4,    -2,     0,    -1,     0,     0,    -1,    -2,    -1,    -2,    -2,    -1,     2,    -2,    -3,    -2,    -2,    -1,    -1,    -2,    -1,     0,     2,     2,    -2,    -2,    -1,    -2,    -4,    -2,     2,     0,    -1,     0,     0,    -2,    -1,    -4,    -3,     0,     2,    -2,    -3,    -1,     1,    -1,    -1,     1,    -2,     0,    -1,     1,     0,    -2,    -2,     0,    -2,    -1,     3,    -2,    -2,     0,    -1,    -2,    -2,    -4,    -4,    -2,    -1,    -3,    -4,    -3,    -3,     0,    -2,     0,    -2,    -2,    -2,    -1,     0,    -4,    -2,     0,    -1,     1,     3,    -2,    -2,     0,     0,     2,    -1,    -3,    -2,    -6,    -4,     1,    -2,    -4,    -1,     2,     2,    -1,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,     0,     1,     3,    -1,     0,     0,     0,    -1,    -2,    -3,    -2,    -4,    -3,     1,     1,     0,    -1,    -1,    -2,    -2,    -5,     0,    -1,    -1,     1,    -2,    -2,    -2,    -1,     1,     2,    -2,     0,     0,     0,    -2,    -3,    -4,    -3,    -5,    -2,     1,     2,     2,     1,    -1,    -2,    -3,    -2,    -1,    -1,    -4,     0,     1,    -2,    -1,     0,     1,     0,    -1,    -1,     0,     0,    -2,    -2,    -5,    -2,    -3,     1,     3,     2,     1,    -2,    -1,    -3,    -3,    -1,     0,     0,    -1,    -1,     1,     0,     0,    -2,    -1,     1,    -1,     0,     0,     0,    -1,    -2,    -2,     0,     0,     2,     1,     2,     1,    -1,     0,    -3,     1,    -2,    -2,     0,    -2,     1,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,     1,     2,    -1,     1,     0,    -1,     0,     1,     1,     2,     0,     2,     0,    -2,    -2,     1,     3,     2,     0,    -1,    -1,    -2,     1,     0,     0,     0,     0,     0,     1,     0,     3,     2,    -1,     2,     2,    -1,     0,     1,     3,     1,     2,     2,     1,     3,     4,     2,     2,     3,     1,    -1,     1,    -1,     0,     0,    -1,     0,     0,     1,     0,    -1,    -1,     1,     3,     3,     2,     2,     4,     2,     2,     2,     2,     1,     2,     2,     3,    -1,    -1,    -1,    -1,     1,     0,    -1,     0),
		    10 => (    0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,     1,    -1,    -1,     1,     1,     0,    -1,     2,     3,     3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,    -1,     2,     2,    -1,    -1,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,    -3,     0,    -3,    -3,    -3,    -3,    -1,    -3,    -2,    -1,     0,    -1,     1,     1,     0,     0,     0,    -1,     0,    -1,     0,     1,    -2,    -5,    -3,     0,     1,     0,    -2,    -2,    -4,     0,     0,     0,    -2,    -2,    -1,     0,     0,    -4,     0,     0,     0,    -1,    -1,     1,    -3,    -2,    -3,    -2,    -3,    -3,    -3,    -5,    -5,    -1,     1,    -2,     1,    -1,     0,     0,     0,     1,     1,    -2,    -3,    -4,     0,     0,    -1,    -1,    -1,     1,    -4,    -2,    -4,    -1,     0,    -4,    -2,    -3,    -2,     0,    -1,    -2,     0,    -2,     0,    -4,    -2,     2,     0,    -4,    -2,    -3,    -2,     0,     0,    -3,     0,    -1,     0,    -2,    -2,     1,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     1,     0,    -2,     2,     3,    -2,    -4,    -4,     0,     0,     0,    -3,    -2,    -1,    -1,     0,     0,    -3,     0,    -1,     0,     0,     0,    -1,    -1,     1,    -2,     0,     2,     1,    -3,     0,    -1,    -2,    -5,    -4,    -3,     1,     5,    -4,     2,     1,    -1,    -1,    -1,    -3,    -2,    -1,     0,     0,     1,    -5,     1,     2,     0,     3,     2,    -2,    -4,    -1,    -2,    -2,    -5,    -2,    -4,    -1,     0,    -1,     3,     0,    -1,     1,    -2,     1,     1,    -1,     1,     0,     0,     0,    -1,    -2,     2,     1,     2,    -1,     2,    -1,    -2,    -2,    -2,    -5,    -4,     0,     0,     0,     2,     1,     0,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -1,     0,    -4,    -1,     1,     0,     0,    -1,    -2,     0,    -1,    -3,    -3,    -3,     0,     0,     6,    -2,    -2,    -2,     1,     1,    -2,    -4,    -3,     0,     0,    -1,     1,    -3,    -5,    -4,    -1,     1,     2,     0,    -4,    -4,    -3,    -4,    -4,    -2,     0,     0,     1,    -1,    -3,     2,     3,     1,    -2,    -6,    -1,     1,     0,     2,     0,    -4,    -5,    -2,     0,     2,     3,     1,    -3,    -4,    -1,    -3,    -4,    -1,    -1,     0,     1,     2,    -2,     5,     2,     1,     0,    -2,     2,     1,    -1,     0,    -2,    -6,    -8,    -3,     0,     1,     3,     4,    -3,    -1,     2,     0,     0,    -2,    -1,     0,     0,    -1,    -3,     0,     3,    -2,     1,     1,     2,     1,     3,     3,    -1,    -4,    -3,    -3,    -2,     2,     4,     4,    -3,     0,     2,     0,    -1,    -1,    -1,     0,     0,    -2,    -4,    -2,    -1,    -1,    -1,     1,     0,     2,     3,     6,    -2,    -6,    -3,    -1,     0,     3,    -1,     1,    -3,     0,     1,    -1,    -1,    -5,    -1,     1,     0,    -2,    -2,    -2,    -1,    -3,    -3,     2,    -1,    -1,     1,     2,    -4,    -6,    -1,     1,     1,     1,     1,    -3,    -4,    -3,    -1,    -2,    -3,    -4,     4,     0,    -1,    -2,    -3,    -1,    -2,    -3,    -1,     1,    -1,     0,     0,     1,    -4,    -3,     0,     1,     1,    -1,     1,     0,    -4,    -2,    -2,    -2,    -2,    -2,     6,     0,    -1,    -2,    -2,    -2,    -4,    -3,    -1,     0,    -1,     1,     0,    -3,    -3,    -2,     0,     3,     1,     1,    -1,    -2,    -3,     0,    -2,    -1,    -2,    -3,    -1,     0,     2,     0,    -2,    -2,    -3,    -4,    -1,     2,     0,     0,     1,    -1,     1,    -1,    -1,    -3,    -2,     2,    -1,    -1,     0,    -2,    -2,     0,    -3,    -2,    -1,    -1,     2,    -1,    -2,    -1,    -2,    -4,    -2,     1,     0,     2,     2,     2,     1,     0,    -4,    -3,    -1,    -2,     0,    -1,     1,    -2,    -1,    -3,     0,     2,     0,     0,     0,    -1,    -3,    -3,    -2,    -3,    -2,     0,     1,     3,     0,     3,     1,    -2,    -2,    -2,    -2,     0,     2,     0,    -1,    -2,     0,     0,     1,     8,     2,     0,    -1,    -2,    -4,    -3,    -2,    -3,    -2,    -1,     2,     0,     0,     0,    -3,     1,     1,     2,    -2,    -4,    -1,    -3,    -3,    -2,    -1,     0,     1,     4,     2,    -1,     0,     0,    -3,    -3,    -5,    -2,    -2,    -2,     2,     4,     1,     1,    -1,     0,    -2,     0,    -1,     0,    -1,    -3,    -3,    -1,    -1,     0,     0,    -4,     0,     0,     0,    -1,     0,     2,     1,    -3,    -4,    -5,    -4,    -3,    -2,     0,    -2,    -3,    -2,    -2,    -1,     2,    -4,    -2,    -2,    -1,     0,     1,     1,     0,     0,     1,     0,    -1,     0,    -2,    -2,    -2,    -4,    -1,    -2,    -5,    -5,    -9,    -8,    -9,    -7,    -4,    -3,    -3,    -3,    -4,    -3,    -2,    -1,     0,     0,     0,     0,     1,    -1,     0,     0,    -2,    -2,    -6,    -2,    -2,    -4,    -3,    -3,    -2,    -2,    -1,    -3,    -3,    -3,    -4,    -4,    -3,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,     0),
		    11 => (    0,     0,     0,    -1,     1,    -1,     1,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     1,     1,     0,     0,    -1,    -2,    -5,    -6,    -4,     1,     1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     2,     0,     0,    -1,    -1,     2,     2,     3,     2,     1,     0,     0,     1,    -3,    -5,    -4,     0,    -2,    -1,    -3,     1,     2,    -2,     0,     0,     1,     0,     0,     1,     1,     1,     1,     2,     2,    -1,     0,    -2,    -1,    -1,    -2,    -2,    -4,    -3,    -1,     0,     1,     2,     0,     0,    -1,    -3,    -2,    -3,    -3,     0,     0,     0,     3,     2,     2,     0,     0,    -3,    -2,    -3,    -3,    -1,    -1,    -6,    -6,    -4,     0,     1,     1,     0,     2,     2,     1,     1,    -2,    -2,     0,     0,     0,     0,     2,     4,    -1,    -2,     0,    -4,     2,     2,     0,    -6,    -6,    -8,    -7,    -3,    -2,     0,    -1,    -1,     0,     0,     0,    -2,    -3,    -2,    -1,     0,    -1,    -1,     0,    -2,    -2,    -2,    -2,    -4,     0,     3,     0,    -3,    -5,    -6,    -4,    -1,    -1,     2,     0,     0,     0,     0,     1,    -4,    -5,    -3,    -1,     0,    -2,    -2,     0,    -1,    -1,    -1,    -3,    -3,    -1,     0,    -3,    -3,    -3,    -5,    -3,     0,     1,     1,     0,     1,    -1,     0,     0,    -3,    -4,    -3,    -1,     0,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -5,    -5,    -5,    -9,    -8,     0,     2,     0,     1,     0,    -1,    -1,     0,     0,    -1,    -3,    -1,    -2,     0,     0,    -1,     0,     0,     0,    -3,    -3,    -4,    -3,    -5,    -4,    -6,    -7,    -4,     0,     3,     1,    -1,     0,     0,     1,     1,     0,     1,    -1,    -2,    -1,    -1,     0,     1,     0,    -1,     1,    -1,    -3,    -4,    -3,    -4,    -2,    -4,    -3,    -2,     4,     2,     1,     4,    -1,     0,     0,    -2,    -3,    -2,     0,    -2,     0,     0,     0,    -2,     1,     0,     1,     0,    -3,     0,    -4,    -3,    -3,    -1,    -2,     1,     3,     0,     2,     1,     1,    -3,     0,    -2,    -1,    -2,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -3,    -1,    -1,    -2,     0,     3,     2,     1,     2,     1,    -1,    -7,    -3,    -3,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,     2,     2,    -1,     0,     2,     1,     1,     2,    -3,    -4,    -8,    -9,    -1,     1,     0,    -1,    -1,    -1,     0,     0,    -1,     2,     3,     0,    -3,     0,     0,     4,     2,     1,     0,    -1,     1,     1,     1,     0,    -2,    -7,    -9,    -5,    -1,     1,     0,    -6,    -4,    -3,     0,     0,     0,     1,    -1,     1,    -1,    -2,     0,     2,     2,    -3,     0,    -1,     0,    -2,     1,     1,    -1,    -5,    -5,    -1,     1,     2,     3,     5,    -2,    -3,    -1,     0,     0,     0,    -2,     0,    -4,    -2,     1,     0,     0,    -1,     2,     2,     0,     0,    -2,     1,     0,     1,     2,     2,     4,     5,     5,     4,     0,    -5,    -2,     0,     0,     0,     0,    -2,    -6,    -4,     0,     0,     0,    -1,     2,    -1,     0,     0,    -1,    -2,     0,     1,     1,     1,     0,     3,     2,     0,     1,     0,     2,     0,     0,     0,    -2,    -4,    -1,     0,     1,     1,     0,    -1,     0,     0,    -2,    -5,    -4,    -2,    -3,    -3,    -2,    -1,    -1,     2,     2,     2,     3,     0,     1,     0,     0,     0,    -2,     1,     2,     2,     0,     1,     0,    -1,     2,    -2,    -3,    -4,    -2,     1,    -2,    -4,    -2,    -2,    -1,     2,     2,     3,     0,     1,     1,     1,     2,     0,     0,    -1,     0,     0,     1,     0,    -1,    -1,     0,    -1,    -1,    -1,     1,     2,     1,    -2,    -2,    -2,    -1,     1,     4,     3,     1,     0,     0,     2,     1,     0,     0,     1,     3,     1,     0,     1,     2,    -1,    -2,    -3,     0,    -2,     2,     3,     0,    -2,    -3,    -2,    -2,     0,     0,     1,     0,     1,     0,     0,     0,    -1,     2,     0,     0,     0,     0,     3,     2,    -1,    -2,     1,     1,     1,     2,     1,    -1,    -2,    -2,    -1,     0,     0,    -1,     2,     3,     4,     0,     0,     0,     0,     1,    -3,    -2,    -3,    -4,    -1,     2,    -1,    -2,     2,     3,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,    -2,     0,     0,     0,     0,     0,     1,    -1,    -2,    -2,    -1,    -5,    -1,     1,    -1,     1,     3,     1,    -4,    -2,    -2,    -3,    -2,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -2,    -3,    -4,    -3,    -2,    -1,    -2,    -2,    -2,    -2,    -2,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     1),
		    12 => (    1,    -1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     1,     0,    -1,    -2,    -1,    -1,     0,     1,     0,     0,    -1,     0,     1,     0,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     1,     2,     1,    -1,    -1,    -2,    -2,    -1,     1,     1,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     1,    -1,    -4,     0,    -2,    -1,    -2,     0,     2,     4,     3,     2,     0,     0,     0,     0,     0,    -1,     0,     0,     1,    -2,    -3,    -2,    -1,     0,     0,     0,     0,     0,    -1,     0,     1,     2,     3,     0,     0,     1,     3,     3,     3,     0,     0,     0,    -1,     0,    -2,    -1,    -2,    -2,    -2,    -3,    -3,    -3,    -1,     1,     0,    -2,     0,     0,     1,     2,     4,     2,     1,     1,     0,     1,     1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     1,    -1,    -2,    -3,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     3,     2,     2,     2,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,    -2,     0,     1,     0,    -2,     0,     3,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,     1,     0,    -2,    -1,     0,    -1,    -1,    -1,     1,     1,    -2,    -2,    -2,     0,     1,    -1,    -2,     1,     3,    -4,    -2,    -2,     1,    -1,     0,    -1,     0,    -1,     0,    -2,    -3,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     1,     0,     0,    -4,    -2,     0,    -2,     2,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -2,     0,    -1,     2,     0,    -2,    -1,    -1,    -1,     0,     1,     1,     0,    -1,    -2,     0,    -1,     0,     0,     1,    -1,    -2,    -1,    -1,    -3,    -4,    -3,    -4,    -1,     0,    -1,    -1,     0,    -2,    -1,    -2,    -1,    -2,     1,     1,    -1,    -2,    -1,     1,    -2,     0,    -1,    -1,    -2,    -2,    -1,     0,    -3,    -4,    -4,    -3,    -1,     0,     0,     1,    -1,    -3,    -2,     1,     0,    -1,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,    -1,    -2,    -2,    -1,     0,    -2,    -2,    -1,    -1,    -1,     1,     2,     0,     0,    -1,    -1,    -1,    -1,     0,    -2,    -2,    -1,    -2,    -3,     0,     1,     1,     0,    -1,    -1,    -2,    -2,    -3,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,     1,     0,    -1,    -1,    -2,    -2,    -1,     1,     2,     0,     0,    -1,    -1,    -1,    -2,    -3,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -2,    -2,    -2,     0,    -1,    -1,    -3,    -2,    -2,    -1,     2,     3,     2,     0,    -2,    -1,     0,    -2,     0,    -1,    -1,     0,    -2,    -1,    -1,    -2,     0,    -1,    -2,    -4,    -3,     0,     0,     0,    -1,    -2,    -2,     1,     2,     3,     2,     0,    -1,     0,     2,     2,     0,    -1,    -1,    -1,    -1,     1,     0,     1,     1,     0,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -2,     0,     2,     4,     3,    -1,    -1,     1,     2,     2,    -1,     0,    -2,    -1,    -1,    -1,    -1,     2,     0,    -1,    -1,    -2,    -2,    -1,    -2,    -3,    -2,    -2,    -3,     0,     3,     3,     3,     1,     0,    -1,     1,     2,     0,    -2,    -1,     0,     0,     0,    -2,     0,     0,     0,     0,    -3,    -1,    -2,    -2,    -1,    -1,     0,     0,     2,     2,     2,     2,     0,     0,     0,     1,     0,    -1,     0,    -1,     0,    -1,     0,     1,     0,     0,    -1,    -1,     0,    -1,     1,    -3,    -1,     1,     2,     2,     2,     2,     4,     5,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -1,     0,     0,     2,     0,    -1,    -1,    -2,    -1,    -1,     1,    -2,     0,     1,     2,     3,     3,     2,     1,    -1,     0,     0,     1,     1,    -1,     0,     0,    -1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,    -1,     1,     1,     3,     3,     1,     0,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,    -1,     0,    -1,    -2,    -1,    -1,    -1,     1,    -1,     1,    -1,    -2,     0,     0,     1,     3,     2,     1,     2,    -2,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     1,    -1,    -1,     1,     0,     0,     1,     1,     0,    -2,    -2,    -2,     0,     1,     3,     3,     0,     1,    -1,     0,     0,     1,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,    -2,     0,     1,     0,     2,     0,    -2,    -1,    -1,     0,    -2,    -1,    -2,     1,     1,     0,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,     0,    -2,    -2,    -2,    -1,    -2,    -3,    -1,    -2,    -2,     0,    -2,     0,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,    -2,    -1,    -2,    -2,    -3,    -2,    -1,    -1,    -2,    -3,    -2,    -5,    -5,    -5,    -4,    -2,    -1,    -2,    -2,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -3,    -2,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     1),
		    13 => (    0,    -1,     1,     0,     0,     0,    -1,    -1,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -3,     2,     1,     2,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     1,    -1,    -2,    -2,    -3,    -2,    -2,    -6,    -9,    -7,    -6,    -1,     1,     0,    -2,    -2,    -2,    -3,     0,     0,     0,    -1,     1,     2,     0,     1,    -2,    -3,    -2,    -1,     3,    -2,     2,     3,    -2,    -1,     0,    -1,    -2,     2,     1,    -2,    -1,     2,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     2,     0,     3,     4,     2,     2,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,    -3,    -3,    -2,    -3,    -1,    -3,    -1,    -1,     0,     0,     1,     1,     3,     3,     1,     0,    -1,     0,     0,     2,     0,     2,     1,     1,     0,     1,     0,    -6,     0,    -2,    -4,    -2,    -1,    -1,     0,    -1,     0,     1,     1,    -2,     4,    -1,     3,     1,     0,     2,     0,     1,     0,     1,     1,    -3,    -2,     0,     0,    -1,    -1,     0,    -4,    -3,    -2,    -1,    -2,    -1,     0,     0,     1,    -2,     3,     1,     0,     1,     0,     4,     2,     1,    -1,     0,    -1,     0,     0,     1,     2,    -1,    -3,     0,    -2,    -6,    -4,    -1,    -3,     1,     0,    -2,     2,     1,     3,     0,     4,     4,     2,     2,     0,    -4,    -3,     0,     0,     1,     0,     0,     0,     1,     1,    -1,    -4,    -4,    -5,    -2,    -1,     0,     0,    -2,     2,     4,     3,     2,     2,     1,    -4,    -6,    -8,    -4,    -3,     1,     1,     2,    -1,     4,     0,     0,     1,    -1,    -3,     0,    -3,    -2,    -2,     0,     0,    -1,     0,     4,     1,    -2,    -4,    -6,   -10,    -5,    -1,    -1,     2,     3,     0,     0,    -2,    -2,     1,     0,     1,     0,    -4,    -3,    -2,    -2,     0,     0,     0,     0,     3,     3,    -2,    -5,    -8,    -5,    -5,     0,     3,     2,     3,     2,     0,    -2,    -3,    -2,    -2,    -5,    -3,    -6,    -3,    -5,    -2,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -3,    -5,    -4,    -2,     0,     2,     1,     1,     1,     1,    -2,    -1,    -2,    -3,    -3,    -4,    -4,    -2,    -1,    -1,    -2,    -2,    -1,    -1,     1,     0,     2,     0,    -2,    -3,    -2,     3,     0,     1,     0,     0,     0,     2,    -1,    -1,    -1,    -3,     1,    -2,    -2,    -2,     1,     0,    -5,    -2,    -1,    -1,     1,     1,     3,    -1,    -2,    -1,    -1,     0,     1,     2,     5,     0,     1,     1,     1,     0,    -3,    -3,     0,     0,     2,    -3,     3,     0,    -2,    -1,    -2,     1,     0,     1,     2,    -3,    -4,    -2,    -2,     1,     3,     0,     0,     2,     2,     2,    -1,     0,     0,     0,    -2,     1,     4,     1,     2,    -1,    -3,    -4,    -2,     0,     1,     1,     3,    -3,    -5,    -5,    -5,    -2,    -1,    -3,    -1,     1,     2,     0,     0,     2,     0,     0,     1,    -1,     3,     3,     0,    -2,    -5,    -2,    -1,    -1,     0,     2,     4,    -1,    -3,    -4,    -6,    -9,   -12,   -10,   -10,   -10,    -8,    -5,    -7,    -2,     4,     0,     1,     1,     1,     5,     2,    -2,    -4,    -2,    -2,     0,    -1,    -4,     2,     2,     2,    -2,    -2,    -4,    -5,    -8,    -9,    -8,    -7,    -5,    -6,    -3,    -1,     1,     3,     3,     2,     3,     3,    -1,    -3,    -4,    -2,     0,     1,    -3,    -1,    -1,     2,     1,    -1,     0,    -3,    -3,    -2,    -2,    -1,    -1,    -3,    -4,    -1,     0,     2,     2,    -1,     0,     6,     0,    -3,     0,     0,     0,     0,     2,     2,     1,     0,     2,     1,     0,    -1,     0,     0,     1,     2,    -1,    -1,    -2,     0,     1,     1,     3,    -2,    -2,    -1,    -2,    -3,    -1,     0,     0,     0,     3,     2,     3,     2,     1,     2,     3,     1,     0,    -1,     0,     2,    -2,     0,     0,    -2,     1,     0,     1,     1,     0,     1,    -4,    -3,     0,     0,     0,     0,     3,     4,     3,     0,     0,     1,     1,     1,    -1,     1,    -1,     1,    -1,    -1,    -1,    -1,    -3,     0,    -2,    -1,    -3,     0,    -3,     0,     1,     1,     1,     1,     1,     0,     4,     2,     1,     4,     2,     0,     3,     2,     1,     0,     1,    -1,    -2,     0,    -1,    -2,    -4,     0,     2,     0,    -3,     0,     0,     0,     1,     0,    -1,    -2,     1,     3,     1,     1,     2,     1,    -1,    -1,    -2,    -3,    -3,    -2,    -1,    -4,    -4,    -4,    -3,    -2,    -1,    -7,    -3,    -1,     0,     0,     0,     0,     1,    -2,     0,     0,    -2,    -1,    -3,    -3,    -4,    -4,    -3,     1,    -1,    -2,     3,     0,     1,    -1,     0,     0,    -2,     0,     0,     0,     0,     0,     1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -3,    -2,    -2,     0,    -2,    -1,    -2,    -1,     0,    -1,    -2,    -3,     0,    -1,     0,     0,     0,    -1,     0),
		    14 => (    0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -5,    -4,    -3,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -5,     0,     0,    -2,    -3,    -2,    -4,    -4,    -4,     0,     1,     1,    -4,    -3,    -1,    -1,    -4,    -2,     0,     0,     0,    -3,     0,     0,     0,     0,     0,    -2,    -5,    -4,    -2,    -1,    -1,    -2,    -4,    -4,    -3,     0,     2,     0,    -3,    -4,     0,     2,     3,     2,    -1,    -3,    -4,    -2,     0,     0,     0,     0,    -1,    -4,    -2,    -2,    -1,     1,     2,     2,     0,    -4,    -4,     0,     0,    -1,    -1,    -1,     2,     0,     2,     1,     0,    -2,    -4,    -2,    -3,     0,     0,     0,    -1,    -1,    -1,     0,     2,     1,     3,     1,     0,    -3,    -3,    -2,     0,    -2,    -3,     1,     1,     2,     0,     0,     0,     0,    -1,     1,    -3,    -1,     0,     0,    -3,    -1,     2,     2,     0,     1,     0,    -1,     0,    -1,     2,     1,     3,     6,     6,     5,     3,     3,     1,     3,    -1,     0,    -1,    -2,     0,    -1,     0,    -4,    -1,     1,     1,     1,     3,     3,     0,     1,     1,     0,     2,     2,     2,     4,     4,     4,     0,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -5,    -2,    -5,     0,     0,     0,     0,     3,     2,     3,    -1,    -2,     0,    -1,     0,    -1,     1,     0,    -1,     0,     0,    -1,     0,    -1,     0,     1,     2,     0,    -4,     0,    -2,    -3,     0,     0,     1,     0,     0,     0,    -4,    -4,    -1,    -2,    -3,    -4,    -2,    -2,    -2,     0,    -2,     0,     2,     0,     1,    -1,    -1,    -1,    -3,     0,    -2,     0,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -1,    -2,    -5,    -6,    -4,    -3,    -2,     0,    -1,    -2,     2,    -1,    -4,    -5,    -3,    -2,    -1,     0,    -2,    -1,     0,    -2,     0,    -2,    -1,    -2,    -2,    -2,    -2,     0,    -2,    -5,     0,    -2,     1,     1,     1,    -1,     1,    -2,    -6,    -6,    -4,    -2,    -4,     0,     0,     0,     1,    -1,     1,     2,     0,     1,     1,     1,     0,     2,     2,    -3,     1,     1,     0,     0,     1,     1,     5,     1,    -1,    -3,    -2,    -4,    -5,     0,    -1,    -2,     0,     2,    -1,     0,     0,     2,     1,     0,     2,     1,    -1,     1,     4,     2,     2,     2,     3,     2,     1,    -1,    -1,    -4,    -2,    -3,     0,     0,    -1,    -5,    -1,     2,    -1,    -1,     0,    -1,     0,    -2,    -1,    -2,    -1,     1,     3,     1,     2,     3,     2,     3,     1,     0,    -1,     0,    -2,     3,     0,     0,     0,     3,     1,     2,    -3,    -1,     0,    -1,    -2,    -5,    -3,    -2,     2,     3,     5,     4,     4,     4,     0,     0,     1,     1,    -1,    -3,    -3,     3,    -3,     0,     0,     0,     2,     2,    -2,    -2,    -1,    -2,    -3,    -4,     0,     1,     4,     5,     4,     5,     1,     3,    -1,     0,     0,    -1,    -1,    -1,     0,     0,    -1,     1,     0,     1,    -1,     4,    -3,    -1,    -1,     0,    -3,    -1,     1,     4,     4,     3,     4,     5,     2,     2,    -2,    -1,     0,     0,     0,    -2,     0,     2,    -3,    -3,    -1,     0,    -1,     3,    -2,    -1,    -2,    -5,    -1,     1,     1,     3,     1,     3,     3,     4,     1,     0,    -2,     1,     0,    -1,     4,    -3,    -4,    -1,     0,     0,    -1,    -2,     2,     0,    -1,     0,     0,     0,     1,     2,     4,     0,    -2,     2,     2,     0,    -2,     2,     1,    -1,     1,     0,     0,    -2,    -2,    -1,     0,     0,     0,    -1,    -2,    -3,    -3,    -2,     0,     3,     2,     3,     2,     2,     2,    -1,     1,     4,     0,     3,     1,     2,     1,     0,     0,    -3,    -4,    -3,     0,    -1,    -1,    -3,    -2,    -4,     0,    -5,     0,     1,     1,     0,    -1,    -3,    -3,     3,     2,     1,     1,    -1,     1,     1,    -1,     1,     1,    -1,    -7,    -4,     0,    -1,    -1,    -1,    -3,    -8,    -4,    -1,    -1,     0,    -4,     0,    -1,    -2,    -1,    -1,     2,     0,    -3,    -1,     1,    -1,     1,     0,     1,    -2,    -3,    -1,    -1,     0,     0,     0,    -5,    -7,    -6,     2,     0,    -3,    -3,    -1,    -2,    -2,    -1,     1,    -1,    -1,    -1,     1,     2,     0,    -1,    -2,     0,    -2,     0,    -1,     0,     0,     0,    -1,    -1,    -5,     1,     0,    -2,    -3,    -3,    -3,    -2,    -1,     0,     0,    -2,     0,    -2,     0,     3,    -2,    -3,    -1,     1,    -3,     2,    -2,     0,     0,     1,     0,     0,     3,     2,    -3,    -3,    -3,     0,    -3,     1,     0,     2,     1,     1,     0,    -2,    -1,    -1,    -3,    -4,    -1,     1,    -1,    -2,    -2,     0,    -1,     0,     1,    -2,     3,     0,    -2,    -5,    -3,    -3,    -3,    -2,    -6,    -4,    -5,    -5,    -3,    -5,    -4,    -2,    -5,    -8,    -8,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -4,    -3,    -3,    -3,    -5,    -1,    -3,    -4,    -2,    -3,    -3,    -3,    -3,     0,     0,     0,     0,     0),
		    15 => (    0,    -1,     0,     1,     0,     0,     0,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     0,    -1,    -2,    -2,    -3,    -2,    -1,    -1,    -3,    -3,    -4,    -2,    -1,     0,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     1,    -1,     0,    -3,    -3,    -3,    -3,    -1,    -1,    -3,    -3,    -4,    -5,    -3,    -1,    -1,    -1,     1,     1,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     1,    -1,    -1,     0,     1,    -1,     1,    -3,    -2,    -4,    -4,    -1,     1,    -3,    -1,    -1,    -1,    -2,    -1,    -2,     1,     1,    -2,    -3,    -3,     0,    -1,    -1,     0,     0,     1,     2,     1,    -2,    -2,     1,    -1,    -2,    -3,     0,     1,    -1,    -2,    -2,    -2,     1,    -1,    -3,    -4,    -3,    -1,    -1,    -2,     0,    -1,     0,    -2,    -1,     2,     1,     0,    -2,    -2,    -1,     1,    -1,     0,     2,    -2,    -3,    -3,    -3,     0,     0,    -1,     0,    -1,    -2,     0,     0,     2,     0,    -1,    -1,    -2,     0,     1,     1,    -2,    -2,    -3,     1,     0,    -1,    -2,     1,    -2,    -3,    -3,    -6,    -6,    -5,    -2,     0,    -1,     1,     1,     1,     2,     0,    -3,    -3,    -3,    -2,     2,     0,    -1,    -4,    -1,     2,    -2,    -1,     0,    -3,    -5,    -3,    -2,    -5,    -5,    -2,    -2,    -2,    -1,     0,    -2,    -5,     0,     0,    -1,    -1,    -2,    -1,     2,    -2,    -4,    -1,     0,     1,     0,     0,    -4,    -1,    -4,     1,     1,     1,    -1,    -2,     0,    -1,     1,     3,     1,    -1,    -1,     0,    -1,     0,     0,    -2,    -1,     0,    -3,    -1,     0,     1,     0,    -1,     2,    -1,     1,     3,     3,     3,     3,     3,     1,     2,     6,     4,     5,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,     2,    -1,     0,     0,     1,     3,     0,    -1,    -1,    -1,     3,     0,     2,     2,     4,     5,     5,     5,     1,     2,     0,     0,     0,     0,     0,    -2,    -3,    -1,     0,    -1,     0,     3,     3,     0,     1,     0,     2,     0,    -1,    -1,     0,     1,     4,     2,     4,     3,     1,     2,     5,    -1,     0,     0,     0,    -1,    -4,    -1,    -2,    -2,     1,     1,     2,     1,     0,    -1,    -1,    -4,    -1,    -1,    -6,    -4,    -2,    -3,    -1,    -1,    -1,     0,     5,    -1,     0,     0,    -1,    -3,     2,     2,    -1,     0,     3,     1,     1,     3,     1,     2,    -4,    -4,    -4,    -3,    -2,    -4,    -1,    -2,    -1,    -2,    -3,    -3,    -2,     0,     1,     0,    -1,    -2,     4,     0,     1,    -1,    -1,     2,     0,     1,     3,     0,    -3,    -2,    -4,    -4,    -1,    -3,    -2,    -1,    -2,    -3,     0,    -4,    -1,    -1,    -1,    -1,    -1,     0,    -4,    -2,    -4,    -1,    -3,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -2,    -3,    -1,    -3,    -1,    -2,    -4,    -2,    -1,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -5,    -4,    -1,    -4,     0,    -1,    -3,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -4,     2,    -3,    -5,    -2,    -4,     0,     0,    -1,     1,     0,     0,     0,    -1,    -3,    -2,    -2,     1,     1,    -2,    -3,    -3,     2,     1,     0,    -2,     0,    -2,    -2,     1,    -2,    -1,    -3,    -2,     0,    -1,     1,    -3,    -1,    -3,     2,     2,    -2,    -1,     0,     0,    -1,     0,     1,     0,     2,     0,     1,     0,    -1,    -3,     1,     2,    -1,    -3,    -3,    -2,     0,    -2,     1,    -3,    -2,    -1,     1,     2,     0,     1,     2,    -1,     0,     1,    -2,     0,     2,     2,    -1,    -1,    -2,     1,     2,     0,    -1,     0,    -4,     1,     0,    -1,     0,     0,    -2,     1,     3,     3,     0,     0,     1,    -2,    -3,     1,    -2,     1,     1,     0,     2,     0,     2,     1,     0,     0,    -3,    -1,    -3,     0,     0,     0,    -1,     2,     0,    -1,     1,    -1,     1,     0,     1,     1,     3,     1,     1,     1,     0,     1,     0,     1,     2,     0,    -1,     0,    -3,     0,    -1,     0,     0,     0,     1,    -1,    -2,    -3,    -1,    -1,     2,     1,     1,     1,     2,     3,     2,    -1,     0,     0,    -2,     1,     1,    -1,    -2,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,    -3,    -3,    -3,     2,     2,     2,     1,     0,    -1,     2,     1,     1,     2,    -1,     1,     0,    -3,    -1,     1,     0,    -3,    -1,     1,     0,    -1,    -1,     0,    -2,    -4,    -2,    -4,    -3,    -4,    -3,    -2,    -3,    -4,    -2,    -2,    -3,    -4,    -3,    -2,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -3,     0,    -1,     1,    -1,    -2,    -5,    -4,    -4,    -4,    -2,    -3,    -1,    -1,     0,     0,    -2,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -4,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0),
		    16 => (    0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     2,     1,     0,     1,     1,     2,     1,    -2,     0,     1,     1,     0,     0,     3,     1,     1,     1,     0,     0,     0,     1,     0,     0,     1,     0,     1,     1,     1,     1,     1,    -1,    -1,     0,    -2,    -2,     1,     1,     4,     4,     0,    -2,    -3,     1,     3,     2,     1,    -1,     0,     0,    -1,     0,    -1,     0,     1,     2,     0,     0,     0,    -1,    -1,     0,    -3,    -1,     2,     2,     4,     2,    -1,     1,     3,     2,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,     3,     3,    -1,    -1,    -2,    -1,    -1,    -2,    -3,    -1,    -2,     0,    -1,     0,    -2,    -1,     0,    -2,     0,    -2,    -2,    -1,     2,     1,     0,     0,    -1,     0,     3,     3,     0,     0,    -1,     0,    -3,    -5,    -2,    -3,    -1,    -1,     1,     1,    -1,    -1,    -4,    -3,     0,    -2,     0,     0,     1,     1,     0,     0,     0,    -2,     2,     2,     0,     0,    -1,    -2,    -4,    -5,    -3,    -1,     1,     3,     0,    -3,     2,     1,    -1,    -4,    -1,    -1,     0,     0,    -1,     1,     0,     0,     0,    -3,     2,     2,     0,    -2,    -1,    -2,    -4,    -5,    -3,     0,     0,    -4,    -2,    -4,    -2,     0,     0,     1,     2,     0,    -1,     1,     0,    -1,     0,     0,     0,    -3,     2,     2,     0,     0,    -2,    -2,    -3,    -5,    -1,     1,     1,    -3,    -1,    -2,    -4,    -2,    -1,     3,     1,    -1,    -1,     0,    -2,    -3,     0,     0,     0,    -1,     3,     2,     0,     1,    -1,    -2,    -3,    -1,     1,     1,    -1,     1,    -3,    -2,    -3,    -3,    -2,    -2,    -2,     0,    -1,     0,     0,    -1,     1,    -1,    -1,    -2,     3,     3,    -1,    -1,    -2,    -1,     0,    -2,     1,     0,     0,    -4,    -2,    -3,    -5,    -4,    -3,    -3,    -2,     0,     1,     0,    -1,     0,     0,     0,     0,    -2,     4,     3,    -1,    -1,    -2,    -3,    -2,     1,     0,    -1,    -2,    -3,    -2,    -3,    -5,    -4,    -3,    -4,    -3,     1,     1,     0,    -1,    -1,     0,     0,    -1,    -2,     2,     3,    -1,    -2,    -2,    -1,     0,     3,     1,    -1,    -1,     0,    -3,    -4,    -3,    -2,    -1,    -3,    -3,     2,     2,     0,    -2,    -1,     0,     0,     1,    -1,     2,     2,     0,    -1,    -1,    -1,     0,     1,     0,     0,     1,     1,     3,     1,    -2,    -1,    -1,    -3,    -2,     1,    -2,    -2,    -2,     0,     0,     0,    -1,     0,     0,     2,     1,     0,     0,    -3,     0,     0,     0,    -1,    -2,     0,     2,    -2,    -3,     0,     2,    -2,    -2,     0,    -1,    -1,    -1,    -1,     1,     0,    -1,    -2,    -1,     0,     1,     0,    -1,    -2,     0,     0,     0,    -4,    -1,    -1,     1,     3,     0,     3,     2,    -2,    -1,    -1,    -2,    -2,    -1,    -2,     0,     1,     0,    -2,    -1,     1,     0,     1,     1,    -3,     0,     3,     3,    -2,    -1,    -3,     0,     1,    -2,     2,     0,    -3,    -1,    -2,    -1,    -1,    -1,    -1,     0,     1,     0,    -2,    -1,    -1,     0,     1,     1,    -3,     2,     4,     1,    -4,    -4,    -2,     0,    -2,     0,     1,     0,    -2,    -2,    -1,    -2,    -3,    -1,    -2,     1,     0,     0,     1,    -2,     0,     0,     0,    -3,    -2,     0,     0,     2,     0,    -3,    -2,     0,     1,     1,     1,    -3,    -2,    -3,    -2,    -3,    -3,     0,    -2,     0,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -3,     0,     3,     2,     2,     0,    -1,    -2,     2,     1,     1,    -2,    -1,    -3,    -2,    -2,    -2,    -2,    -1,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -3,    -4,    -3,     0,     1,     2,     0,     0,    -1,     2,     0,     1,     1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -4,    -3,    -3,     0,     2,     0,    -1,    -1,    -1,     0,     0,    -3,    -2,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,    -1,     0,    -1,     1,     0,    -2,    -4,     0,    -1,     0,     0,     2,     2,    -1,    -3,    -3,     1,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -3,    -3,    -2,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -2,     0,     1,     1,     0,     3,     5,     2,    -3,    -5,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     0,    -1,    -1,     0,     1,     1,    -1,     0,    -1,     0,    -1,    -1,    -2,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
		    17 => (    0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,     0,     1,     1,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,     0,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -2,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,    -2,     0,    -1,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -2,    -1,    -2,     0,     0,    -1,    -1,    -1,    -1,    -3,    -1,     0,    -1,     1,     0,     0,     0,    -1,     0,    -3,    -1,     0,    -4,    -4,    -2,    -4,    -6,    -5,    -5,    -4,    -2,    -1,     0,     0,     0,    -2,    -3,    -2,    -3,    -1,    -1,    -1,     0,     0,     1,     0,    -1,    -3,    -1,    -1,     1,     1,     0,    -3,    -2,     0,     0,    -3,    -4,    -5,    -9,   -10,    -9,    -9,    -5,    -1,    -3,    -2,    -1,    -1,     0,     0,     0,     3,     3,     0,     0,     0,    -2,    -2,    -3,    -4,     1,     2,     1,    -1,    -5,    -4,     0,    -1,     0,    -1,     3,     2,     1,    -2,    -3,    -4,    -1,     0,     6,     5,     4,     0,    -1,     0,     3,    -1,     0,     0,    -2,     1,     0,    -2,    -3,    -3,    -1,     0,    -1,    -2,     0,    -1,     1,     1,     0,    -3,    -1,    -4,     6,     2,     1,    -1,    -2,    -2,    -1,    -3,     0,     3,     0,     1,    -2,    -2,    -1,    -2,     1,     1,     0,    -1,    -2,    -1,     2,     4,     1,    -2,    -2,     0,     4,    -3,     0,     1,     0,     2,    -1,    -1,     0,     1,     1,     1,     0,     3,     0,    -2,     1,     2,     2,     0,     1,     1,     1,     4,    -1,    -4,     0,     1,     3,     2,     0,     1,     1,     2,     1,     1,     0,     0,     2,     2,     3,     0,    -3,    -2,     1,     0,     2,     3,     2,    -2,    -1,    -2,    -1,    -3,     1,     0,     1,     2,     3,     1,     3,     1,    -1,    -3,     3,     1,     4,     5,     0,    -4,    -3,    -1,    -1,     3,     2,     2,    -1,    -2,     0,    -1,    -3,    -1,     0,     1,     1,     1,     2,     0,     2,     1,     3,     2,     1,     3,     1,     3,    -8,    -8,    -1,     1,     1,     2,     0,     1,    -1,    -3,    -3,    -2,    -2,     0,     2,     0,     1,     3,    -1,    -1,     3,     2,     3,     2,     0,     0,     0,    -2,   -10,    -7,    -4,     2,     0,     2,    -2,     0,     1,    -2,    -4,     0,    -3,    -1,    -1,    -1,     2,     5,     2,    -1,     3,     1,    -1,     0,     2,     3,     1,    -5,   -14,    -6,    -2,     1,     0,     3,     1,     0,    -1,    -1,     0,     0,    -2,    -2,     0,    -1,     0,     1,     2,    -5,     1,     2,     2,    -2,    -1,     4,    -2,   -12,    -8,    -4,    -2,     2,     2,     1,     2,     0,    -1,     0,    -2,    -3,    -3,     0,    -1,    -1,    -1,     1,     1,    -2,    -2,     0,     3,    -1,     0,     4,    -5,   -12,    -2,     0,    -1,    -1,     0,     2,     2,    -2,     0,     2,    -1,    -1,    -2,     0,    -2,    -1,     0,     2,    -1,     0,    -2,     0,     0,    -2,    -4,    -6,    -8,    -6,    -1,     1,     0,    -1,    -1,     2,    -2,     1,     0,     2,    -6,    -8,    -1,     0,    -3,     1,    -1,     3,    -5,    -2,    -1,     1,     0,    -3,    -6,   -10,    -3,    -1,     2,     3,     0,     1,     1,     1,    -2,     2,    -1,    -2,    -7,    -7,     1,     0,    -1,     0,     2,     1,    -4,    -1,     1,     1,    -6,    -6,    -7,    -8,    -3,     0,     0,     1,     0,    -1,    -2,     1,     0,    -1,    -3,    -5,    -6,    -3,     2,     0,    -1,     0,     2,     0,    -2,    -1,    -1,    -3,    -6,    -6,    -8,    -2,     3,     2,    -2,     0,    -2,    -1,     0,    -2,    -1,    -2,    -5,    -4,    -6,    -2,     0,     0,     0,     0,     0,    -1,    -3,    -6,    -2,    -5,    -5,    -4,    -2,     4,     1,    -1,    -2,    -1,    -4,    -2,     0,     2,     0,     0,    -1,     0,    -1,     8,     0,    -1,     0,     0,     1,    -1,    -1,    -4,     0,     0,     0,     1,     1,     0,     1,    -2,     0,     0,     0,    -1,     0,     1,     2,     0,    -1,     0,    -1,     0,     0,    -2,     0,     0,     0,    -1,    -4,    -2,     2,     3,     2,     2,     0,     1,    -4,     0,     1,     0,     0,    -2,    -1,     1,    -3,    -1,    -1,    -5,    -3,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,     3,    -1,    -3,     2,     0,     0,     1,     1,     0,     2,    -1,    -2,    -1,    -4,    -2,    -1,     1,    -4,    -4,    -1,    -4,     1,     0,     0,     0,     0,     0,    -4,    -6,    -2,    -1,     0,     0,     1,     1,     1,     0,     2,     0,     1,     2,    -3,    -1,    -1,     1,     0,    -3,     1,    -1,     0,     0,     0,     0,     1,     0,    -5,    -5,    -4,    -4,    -2,    -2,    -2,    -3,     0,     2,     3,     0,     2,    -1,     0,     1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     1,     1,     1,     1,     2,     1,     1,     1,    -1,    -1,     1,    -1,    -1,     3,     3,    -2,     1,     4,     1,     2,     0,     0,     0,     0),
		    18 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -3,    -4,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,    -2,    -1,    -1,    -4,    -5,    -2,    -1,     0,    -1,    -3,    -2,    -1,     1,    -2,    -5,    -4,    -4,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -2,     0,    -2,    -2,    -5,     1,     1,    -1,    -2,    -2,    -4,    -5,     0,     1,     0,     2,     1,     5,     4,     2,     2,    -2,    -1,    -1,     0,     0,     1,     0,    -3,    -3,    -5,     0,     0,    -2,    -3,     0,    -2,    -4,    -3,     2,     0,     1,    -1,    -1,     1,     3,     4,     2,     1,     0,     4,     2,    -1,    -1,     0,    -2,    -3,    -5,    -2,     0,     0,     1,     0,     0,     0,    -2,    -2,    -1,     0,     0,    -2,    -3,    -1,     3,     2,     1,     4,     4,     2,    -2,     0,     0,     0,    -2,    -3,    -1,    -3,     1,     1,     1,     0,    -1,    -2,     1,     0,     1,     0,    -3,    -3,    -1,     2,     0,    -1,    -3,     1,     0,     5,     0,    -3,     0,    -3,    -2,    -1,     0,    -3,     1,     3,     0,    -2,    -1,    -1,     0,     0,     0,     1,    -3,    -1,     2,     1,    -2,     0,     1,     1,     1,     0,    -1,    -3,    -1,    -1,    -2,     1,     3,    -1,     2,     3,    -2,     1,    -1,     0,     1,     3,    -1,    -4,    -2,    -1,    -2,    -3,     0,     3,     2,     0,     1,     2,     2,     1,     0,     1,     0,     2,     1,    -3,    -1,    -1,    -1,    -1,     1,     2,    -1,    -1,    -3,    -4,     0,    -1,    -2,     1,     1,     1,     0,     3,     1,     1,    -3,    -7,     0,    -1,    -1,    -2,     0,    -3,    -2,    -3,     1,     2,     2,     1,    -1,    -2,    -3,    -2,     1,     3,    -1,    -1,    -1,    -1,     0,     2,     0,    -5,    -3,    -5,     0,     0,    -2,    -3,    -2,    -2,    -1,     0,    -1,     2,     0,     3,     2,     0,    -1,    -2,     0,    -1,    -1,    -4,    -2,    -5,    -2,     2,     4,     0,     4,    -3,     0,     0,    -3,     3,    -2,     3,     0,     1,    -3,    -1,     0,    -2,     1,     2,    -1,    -2,    -2,     0,     1,     2,    -3,    -1,     3,     5,     5,     2,     1,    -5,     0,     0,    -3,     3,    -1,    -2,    -5,    -2,    -2,    -3,    -1,    -1,     0,     1,     0,    -1,    -3,     1,     0,     1,     2,     4,     6,     5,     3,    -2,    -2,     1,    -1,     0,     0,    -4,     0,    -4,    -2,    -2,    -3,    -4,     0,    -2,     0,     3,     1,     0,    -3,     2,    -3,     1,     0,     3,     0,     4,     3,    -2,    -4,     0,     0,     0,    -1,     2,    -1,     1,     0,    -1,     0,    -4,    -1,     1,     2,     1,     0,    -1,     2,    -5,    -2,     1,    -2,    -4,    -1,     3,     3,     0,    -4,    -3,     0,    -1,    -1,     2,    -3,     3,    -1,     1,    -2,    -3,    -1,     0,     3,     1,     0,     1,    -3,    -1,    -1,    -3,    -4,    -3,    -2,     2,     1,     1,    -3,    -3,     0,     0,    -1,     1,    -5,    -1,     0,     2,    -1,    -2,     0,     2,     2,    -2,     3,     2,    -1,    -1,    -4,    -4,    -2,    -3,    -2,     0,     0,     0,    -1,    -2,    -1,     0,    -1,    -2,    -3,    -2,    -1,    -2,    -2,     2,     2,     3,    -2,    -5,    -1,     3,     0,    -1,    -1,     1,    -1,    -5,    -1,     0,    -3,     0,     0,    -2,     0,    -1,    -1,    -1,    -4,    -1,    -1,    -3,     3,     1,     3,     3,    -3,    -5,    -2,     1,     1,     2,    -2,    -1,    -2,    -3,     0,    -2,    -2,     0,    -2,    -1,     0,     1,    -1,    -2,    -6,    -1,    -3,     2,     1,     1,     3,     3,     1,    -1,    -1,     0,     0,    -1,     0,     0,    -2,    -2,    -2,    -2,     0,     1,    -3,     0,    -1,    -2,    -1,     0,    -5,    -6,     1,     1,     1,     1,     0,     0,     1,    -2,    -2,     1,    -3,    -1,     1,    -1,    -5,    -3,     0,    -2,    -1,     1,    -3,     0,    -1,    -1,    -1,    -2,    -3,    -7,    -3,     1,    -1,     0,     0,     1,    -1,     1,    -2,     0,    -5,     0,     0,    -5,    -7,    -3,    -2,    -2,     0,     2,    -4,     0,     0,     0,    -2,    -3,    -4,    -5,    -2,     0,     3,    -2,    -3,     0,     2,     1,     1,    -2,    -1,     3,    -3,    -7,    -7,    -3,    -3,    -1,     2,     1,    -4,     0,     0,     0,     0,     0,    -4,    -6,    -3,     0,     1,     0,     0,     1,     3,     3,     1,    -1,     1,    -2,    -3,    -4,    -2,    -2,    -2,    -1,    -2,    -3,    -3,     0,     0,     0,    -2,    -1,    -2,    -3,    -1,    -1,    -2,    -2,     3,    -3,    -4,    -2,    -1,     2,    -1,     0,     1,     2,     2,    -1,    -2,    -1,    -3,    -2,    -2,     0,     0,     0,     0,     0,    -1,    -2,    -3,     0,     0,    -2,    -5,    -3,    -3,    -4,    -5,    -5,    -2,    -1,     0,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -2,    -2,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0),
		    19 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,     0,     1,    -1,    -1,     0,    -1,    -1,    -2,    -1,    -1,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -3,     0,     0,    -2,     0,     0,     0,     0,     0,    -2,    -4,    -2,     1,     4,     1,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -2,    -2,     0,    -1,     0,     1,     0,    -2,    -3,    -4,    -6,    -6,    -6,    -4,    -5,    -6,    -3,    -3,    -4,    -2,    -3,    -2,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -3,     0,    -1,    -2,    -5,    -6,    -8,    -8,    -6,    -5,    -2,    -2,     0,    -1,    -2,    -5,    -3,    -3,    -3,     0,     0,    -1,    -2,    -2,     1,     0,    -2,    -2,    -2,    -4,    -3,    -7,    -8,    -4,     0,    -1,     0,     3,     2,    -2,    -1,    -1,    -3,    -4,    -2,    -2,    -3,    -3,     0,    -2,    -2,    -1,    -1,    -1,    -2,    -3,    -1,    -6,    -8,    -5,    -2,     1,     1,     4,     3,    -2,     2,     0,     2,    -2,    -1,     1,    -3,    -3,    -2,    -2,    -3,    -2,    -2,     0,    -1,     0,     4,    -2,     0,    -3,    -3,    -2,     1,     1,    -1,    -2,     0,     1,     1,     2,    -4,     0,     3,     2,    -4,    -4,    -2,    -1,     0,    -2,     2,     2,     2,     1,    -1,    -2,    -5,    -1,     1,     1,     2,     0,    -3,     0,    -3,    -6,    -2,     0,    -2,    -2,     5,    -2,    -2,    -4,    -1,    -2,     0,    -3,    -5,     2,     2,     1,    -2,    -4,    -2,     1,     1,     3,     1,     1,     0,     0,    -3,    -3,     0,     0,    -1,     0,     0,    -2,    -1,    -4,    -3,    -2,     0,    -1,    -2,     0,    -1,     0,    -1,     0,    -2,    -1,     0,     2,     0,     1,     0,     0,     1,    -1,     2,     0,    -1,     0,     1,    -1,    -1,    -1,    -3,    -1,     0,     0,     1,     0,     1,    -2,    -3,     0,     0,    -2,     1,     1,     1,     0,     5,     3,     2,     0,     1,    -3,    -6,    -1,    -3,    -1,    -2,    -4,    -3,    -4,     0,    -1,    -1,    -1,    -1,    -2,     0,    -2,     0,    -1,     3,     4,     2,     2,     2,     2,    -1,     0,    -1,    -8,    -7,    -3,    -4,    -1,     0,    -2,    -2,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     1,    -2,    -2,     0,     0,     0,     0,     2,     1,     0,     0,     0,    -6,    -4,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -3,    -1,    -1,    -2,     0,     0,     1,    -2,     1,     0,     1,     1,     2,     1,     3,     1,     2,    -9,    -6,    -2,    -3,     1,     1,    -1,     3,     0,     0,     0,    -2,     0,    -1,    -5,    -4,    -1,     0,     0,     5,     2,     2,    -2,    -2,     0,     0,     0,    -7,   -10,    -3,     3,     1,     0,     4,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,    -5,    -4,    -2,    -3,    -1,     2,     1,    -3,     0,     2,     0,    -2,    -2,    -5,    -5,     2,     3,    -3,    -2,     3,    -1,    -3,     0,     2,     0,    -2,    -1,    -2,    -2,    -1,    -6,    -6,    -2,     0,    -1,    -4,     1,     1,     1,    -3,    -2,    -4,    -4,     3,     3,     0,    -1,     0,     0,    -3,    -2,     0,    -2,    -2,    -1,    -3,    -4,    -3,    -5,    -8,    -6,    -5,    -5,    -1,     0,    -1,     0,    -3,    -2,    -4,    -1,     2,     4,     1,    -1,    -1,     0,    -1,    -2,     0,     0,    -1,    -2,    -3,     0,    -2,    -5,    -4,    -2,    -3,     0,     0,    -2,     0,    -4,    -3,    -3,    -3,     2,     1,    -1,    -1,    -1,     2,     1,     0,     0,    -1,     0,    -2,    -2,    -2,    -1,     1,    -1,     0,     0,     0,    -2,     0,    -1,    -1,     0,    -1,    -4,    -2,     3,     3,     0,     0,     3,    -4,     3,    -2,    -1,     0,     0,    -1,    -3,     0,     1,    -2,     0,     1,     0,    -1,     1,    -2,    -3,    -2,    -1,    -2,    -5,    -2,     2,     4,     0,    -1,     2,     4,     0,     0,     0,     0,     0,    -1,    -1,    -3,     1,    -1,     3,     0,     1,     0,    -3,    -1,    -2,    -3,    -3,    -2,    -3,    -3,     1,     5,     1,     0,    -1,     3,    -2,     0,     0,     0,     0,    -1,    -2,    -1,     1,     0,     2,     0,     0,    -1,    -2,     0,    -2,    -2,    -3,    -2,    -1,    -4,    -2,     1,     0,     0,     0,    -3,    -2,    -2,     0,    -1,     0,     2,    -1,     3,    -1,     0,     2,     0,    -3,    -2,     2,    -1,     1,    -2,    -2,     5,     2,    -2,    -1,     1,     1,    -1,     1,    -3,    -3,    -2,     0,    -1,     0,     0,     3,     4,     0,     0,     2,    -1,     2,    -1,     2,     4,     2,     3,     1,     7,     6,     0,    -4,     0,     2,    -1,    -1,     0,    -1,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     2,     4,     4,     4,     5,     3,     2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0),
		    20 => (    0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     1,     0,    -1,    -2,    -2,    -3,     1,     1,     0,     0,     2,     1,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,    -1,    -1,     0,    -1,    -2,    -2,     0,     0,    -1,    -3,    -2,     0,     0,     0,     0,     0,    -1,    -3,    -2,    -1,    -1,     0,     1,     0,     0,     0,     1,     0,    -2,    -1,     0,    -3,    -5,    -2,    -2,    -2,    -4,    -3,    -1,    -1,     0,    -1,    -1,    -3,    -3,    -2,    -4,    -2,    -2,    -3,     0,     0,     0,    -1,    -2,    -2,    -4,    -1,    -1,    -1,    -1,     0,     0,    -2,    -2,    -2,    -1,     1,     2,     1,     1,    -1,    -2,    -2,    -2,     0,    -5,    -2,     1,     0,     0,    -1,    -1,     1,    -2,    -1,    -2,    -2,     0,     1,     0,    -1,    -2,     0,     1,     3,     2,     3,     2,    -1,    -1,    -4,    -3,     0,    -4,    -2,     0,     0,     0,    -2,     0,     0,     0,     0,    -1,    -3,    -2,    -1,    -1,    -2,     0,    -1,     2,     2,     2,     2,     1,     3,     1,     0,     0,    -1,    -3,    -1,     2,    -1,    -2,    -3,    -2,    -1,    -1,     0,     0,    -3,    -1,    -1,     0,    -1,     0,     1,     0,     1,     1,     0,     1,     1,    -1,     1,     0,     0,     1,    -2,     0,     1,    -4,     1,    -2,    -2,    -1,    -2,    -1,    -3,    -2,    -2,     0,     0,     0,    -1,    -2,    -1,     0,     1,     0,     0,     1,     0,     0,     0,    -2,    -2,     0,    -1,    -1,     1,     0,    -2,    -2,    -4,    -1,    -2,    -2,    -2,     0,    -1,    -1,    -3,    -3,    -1,    -2,    -3,    -3,    -2,    -2,    -1,    -1,    -1,    -3,    -3,     0,    -1,     0,     2,     0,    -3,    -3,    -1,     0,    -2,    -2,    -3,    -4,    -4,    -4,    -2,    -3,    -2,    -1,    -3,    -3,    -5,    -5,    -1,    -1,    -2,    -1,    -3,     0,     0,     3,    -3,     0,    -2,    -1,     1,    -1,    -4,    -3,    -3,    -3,    -3,    -2,    -2,    -1,    -2,    -1,    -1,    -1,    -2,    -2,     0,    -1,    -1,    -1,    -1,    -1,     0,     1,    -4,     1,    -1,     0,     0,    -2,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     1,    -1,    -1,    -2,    -2,    -1,     0,     1,     0,     1,     0,    -1,     0,    -1,    -2,     0,    -2,    -1,    -1,     0,     0,    -2,    -1,     0,     2,     0,    -2,     0,     1,     1,     0,     0,    -3,    -2,     0,     0,    -1,    -2,     0,     0,     0,     1,     1,     0,    -3,    -2,    -2,    -1,    -4,    -3,    -2,     0,     0,    -2,    -1,    -1,     0,    -2,    -1,     2,    -3,     0,     0,     0,    -1,    -3,     1,     1,    -2,     1,     1,    -2,    -3,    -4,    -2,    -6,    -6,    -3,    -2,     0,    -1,     0,     1,     0,    -2,    -2,     0,     0,    -4,    -1,     0,     0,    -2,    -1,     3,     0,    -2,    -2,     0,    -4,    -4,    -3,    -5,    -5,    -4,     0,     0,     1,     0,     0,     2,    -1,    -2,     0,     1,     1,    -5,     1,     0,     0,    -2,    -1,     1,     0,     1,     0,     0,     0,    -3,    -3,    -1,    -2,    -1,     2,     1,     2,     0,     1,    -1,    -1,    -1,     1,     1,     0,    -4,     1,    -1,     0,    -1,     0,     1,    -1,     1,     1,     1,     1,    -1,    -2,    -3,    -2,     0,     2,     2,     1,     0,    -1,    -1,    -1,     0,     1,     0,     0,    -3,    -2,     0,     0,     0,     0,     0,     0,    -1,     2,     1,     1,    -1,    -1,     0,    -2,     0,     1,     0,    -2,    -4,    -2,     0,     2,     1,     0,     2,    -4,    -2,    -1,     0,     1,     1,     1,     0,     1,    -1,    -1,     0,    -1,     0,    -1,    -1,    -2,     0,     0,    -2,    -3,    -1,     0,     0,    -1,     0,     1,     1,    -1,    -1,    -1,     1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -3,    -2,    -4,    -2,     0,    -1,    -2,     0,     0,     0,    -2,     0,     1,     1,     0,     1,     0,     0,    -1,    -2,     0,     1,     0,     0,     0,    -1,     0,    -3,    -1,    -1,    -1,     0,    -2,     0,    -2,     0,     0,    -1,     0,     1,     1,     0,    -1,     0,     0,     0,     0,    -2,    -2,    -2,    -1,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     1,     1,    -1,     1,     1,     0,    -3,    -2,    -1,     0,     0,     0,     0,    -1,    -2,     1,    -3,    -1,    -1,    -2,    -5,    -3,    -3,    -2,    -3,    -2,    -1,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -2,    -2,    -2,    -1,    -2,    -3,    -4,    -4,    -4,    -3,    -3,    -1,    -1,    -4,    -2,    -2,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -4,    -2,    -1,    -2,    -2,    -1,    -1,    -2,    -2,    -3,    -3,    -4,    -4,    -4,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,     0,     0,     1,    -1),
		    21 => (    0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,    -2,     3,     3,     0,    -2,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -3,    -3,    -2,    -5,    -1,    -3,    -3,    -1,    -3,    -1,    -1,    -1,    -3,    -4,    -3,    -2,    -1,     0,     0,     0,    -1,     4,     3,     0,    -2,    -1,     3,     2,     3,     1,    -4,    -3,     4,    -1,    -4,    -3,    -1,    -1,    -2,    -1,    -6,    -4,    -3,    -2,    -1,     0,     0,     0,    -1,     4,     4,     0,    -1,     0,     4,     4,     3,     2,    -1,     0,     1,     0,     0,    -3,    -3,    -1,     0,    -2,    -4,    -2,    -2,    -2,    -4,    -5,    -4,     0,     0,     4,     1,     1,     2,     2,     4,     1,     3,     5,     5,     2,     3,     0,    -1,    -2,    -1,    -2,     1,    -1,    -3,    -2,     2,     0,    -7,    -3,    -3,     0,     0,    -2,     0,     2,     1,     2,     4,     1,     1,     5,     2,     1,     2,     0,     0,    -1,     0,     0,     0,     0,    -3,    -2,     2,     0,    -3,    -4,    -2,     0,    -3,    -4,    -4,    -5,     2,     3,     5,    -2,    -2,     2,     1,     2,    -1,     2,     0,     1,     1,    -2,    -2,     2,    -1,     2,     2,    -1,    -3,    -7,    -4,    -1,    -3,    -4,    -6,    -6,    -1,     3,     4,    -2,    -4,     2,    -2,     1,     3,     2,     2,     1,     2,     3,     1,    -1,     0,     1,     0,    -3,    -3,    -7,    -3,     1,    -1,    -4,    -5,    -4,    -2,     0,     3,    -1,    -1,    -3,    -3,    -1,     3,     1,     1,     0,     3,     4,    -1,     1,     1,     0,    -2,    -3,    -3,    -3,    -4,     0,    -2,    -4,    -5,    -4,    -3,    -2,     0,     2,    -2,    -3,    -3,    -1,     2,     0,     0,     3,     4,     1,    -1,     0,    -2,    -2,    -4,    -4,    -3,    -5,     0,     0,     0,    -1,    -3,     0,    -1,    -1,     3,     1,     0,    -2,    -3,    -1,     1,     0,     1,     4,     7,     2,     0,     3,    -3,    -4,    -3,    -4,    -4,    -5,     4,     0,     1,    -5,    -2,     0,     1,     3,     3,     1,    -2,    -1,     0,     1,     0,     1,     3,     3,     4,     2,    -1,     0,    -4,    -4,    -1,    -4,    -1,     0,     3,     0,    -1,    -3,     0,    -2,     2,     3,     1,    -2,    -3,    -1,    -2,    -1,    -1,     0,    -1,     0,     5,    -2,     0,     0,    -3,    -3,    -6,    -5,     1,     3,     0,     0,    -1,     0,     1,    -2,     1,    -2,    -3,     0,    -2,    -3,     1,    -1,    -1,     2,     0,    -1,     0,    -5,    -2,     1,    -1,    -1,    -2,    -4,     2,     5,     0,     0,    -1,     0,    -1,    -4,    -3,    -1,     0,    -1,     0,     1,    -2,     0,     0,     1,     0,    -1,    -3,    -5,    -4,    -1,     1,    -4,    -4,    -6,    -2,     0,    -1,     0,     0,     1,    -4,    -3,     1,     0,    -2,    -3,     2,     0,    -1,     0,     2,     2,    -3,    -5,    -5,    -1,    -2,     0,     0,    -1,     0,     2,     0,    -2,    -1,     0,     0,    -1,    -6,    -3,     1,    -1,    -2,    -2,    -3,    -2,     2,     2,     1,     2,    -5,    -4,    -5,    -4,     0,     1,     2,     3,     4,     3,     0,    -3,    -3,    -1,     0,    -1,    -5,    -4,    -4,    -6,    -4,    -3,    -2,    -1,     0,    -1,     1,     0,    -1,    -3,    -3,     3,     3,     4,     3,     1,     0,     1,     2,    -2,     1,     0,     0,     1,    -7,    -5,    -2,    -1,    -1,     0,     1,     2,     2,    -2,    -2,     1,    -1,    -1,     0,     0,     2,     6,     3,     0,     3,     4,     3,    -1,     0,     0,     0,    -3,    -5,    -1,     0,     2,    -1,     1,     3,     4,     1,     0,    -1,    -1,     0,     0,     2,     4,     4,     6,     2,     0,     0,     2,     1,     0,     0,     1,     1,    -4,     0,    -1,     1,     0,     0,    -1,     1,     3,    -1,    -3,    -2,    -1,     2,     1,    -1,     5,     4,     5,     4,    -1,    -1,     2,     1,    -2,     0,     0,     0,    -4,    -3,    -1,     1,     0,    -1,     2,     1,     1,    -1,    -2,     0,    -2,     3,    -1,     1,     8,     5,     3,     4,     1,     0,     2,     3,     0,     0,     0,     0,    -1,     0,    -3,    -1,     0,     0,    -3,    -1,    -1,     0,     3,     1,     2,     5,     2,     3,     4,     2,     3,     1,     0,    -3,    -4,    -2,     2,    -1,     0,     0,     0,    -1,    -3,    -3,    -3,     0,    -4,    -4,     1,    -2,     0,     1,     0,     2,     1,     4,     1,     1,     0,     3,     1,    -3,    -2,     1,     1,     0,     0,     0,     0,    -2,    -3,    -6,    -6,    -6,    -4,    -9,    -9,    -7,    -1,     0,    -2,     0,    -3,    -7,    -6,    -8,    -7,    -5,    -2,    -2,    -2,    -2,    -1,     1,     0,     0,     0,    -1,    -4,    -8,    -7,    -5,   -10,    -9,    -5,    -4,    -5,    -6,    -1,    -1,     1,    -4,    -3,    -1,    -2,    -3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -4,    -2,    -1,    -1,    -2,    -1,    -1,     0,     1,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1),
		    22 => (    0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -4,    -3,    -2,    -2,    -2,    -3,    -1,     0,     0,    -1,    -2,    -6,    -3,    -2,    -2,    -1,     1,     0,     0,     1,     0,     0,    -1,    -1,    -2,    -1,     0,    -2,     1,     3,     3,     3,     2,     2,    -2,    -1,    -1,    -2,    -3,    -4,    -4,    -2,    -1,    -1,     0,     3,     0,     0,     0,     0,    -1,    -3,    -3,     3,     2,    -2,     0,     5,     2,     3,     3,     1,     1,    -1,     0,     0,    -3,    -3,    -1,     2,     0,    -3,     0,     1,     0,     0,     0,     0,     0,    -1,     3,    -1,     1,     3,     1,     4,     3,     2,     2,     2,     0,     1,     1,     2,     1,    -1,     0,    -2,    -1,    -2,    -1,    -2,    -1,    -1,     0,     0,     1,     1,     2,     2,    -1,     1,     2,     1,     0,     0,     0,     1,     1,     1,     4,     1,     3,    -1,    -1,    -1,     1,    -2,    -2,    -2,    -1,    -1,     0,     0,     1,     0,     0,     1,    -1,     0,     2,     1,     1,     0,     1,     0,     3,     5,     3,     0,     1,     1,    -3,    -2,    -2,    -3,    -6,     0,    -1,    -1,     0,     0,     1,    -2,     0,    -1,     2,     2,     2,     2,     0,     1,     0,     1,     0,    -2,     0,     0,    -1,    -1,    -2,    -3,    -2,    -6,    -2,     0,    -2,     0,    -2,     2,    -2,    -3,     0,    -2,    -1,     0,    -1,     0,     3,     1,    -2,    -1,    -1,    -1,    -1,     0,     2,     1,     0,     0,    -4,    -4,    -2,    -2,    -1,    -2,     0,     0,     0,    -3,    -3,    -4,    -3,    -3,    -4,    -4,     0,     0,     0,    -2,    -3,    -3,     0,    -1,     0,    -2,     0,    -1,    -1,    -4,    -5,    -3,     1,    -1,     0,     0,     0,    -4,    -3,    -1,     1,    -2,    -4,    -5,    -3,    -4,    -3,    -6,    -4,    -4,    -1,     1,     1,     2,     1,    -2,    -6,    -2,    -1,    -1,     0,    -2,     0,    -2,    -2,    -3,    -2,    -4,    -4,    -8,    -7,    -7,    -7,    -7,    -6,    -4,    -4,    -5,    -3,     0,    -2,     2,    -1,    -2,    -1,     2,     2,     0,    -4,    -1,     0,    -3,    -3,    -3,    -5,    -5,    -5,    -8,    -6,    -4,    -3,    -5,    -1,     0,    -1,    -2,    -1,    -1,    -1,     2,    -1,    -1,    -1,    -2,    -5,     1,    -3,    -1,     0,    -3,    -1,    -2,    -4,    -4,    -2,     0,    -1,    -2,    -2,     2,     5,     3,     2,    -1,    -1,     0,     2,    -1,    -1,    -3,    -2,     0,     2,     2,     2,     1,    -1,    -3,    -3,     3,    -1,    -1,     1,     1,     2,     3,     4,     5,     5,     1,     3,     1,     1,     0,     1,    -1,     0,    -2,     0,     0,     3,     0,     3,     3,     0,    -1,     0,     2,     2,     4,     2,     0,     1,     4,     3,     3,    -1,     0,     1,     2,     0,    -1,     1,    -1,    -2,     1,    -1,    -1,    -1,     3,     3,     4,     0,     0,     2,     0,     3,     1,     2,     1,     0,     1,    -1,     2,     0,    -1,     1,     1,     1,     3,     2,     2,     3,     3,     2,     1,    -1,     5,     4,     1,     0,     0,     2,    -1,     1,     2,     3,     0,     3,     0,     2,    -1,     0,    -3,     1,     2,    -1,     2,     2,     1,     0,    -2,     1,    -1,    -5,     3,    -1,     2,     0,     0,    -1,    -4,    -2,     3,     2,     3,     4,     2,     0,    -2,    -3,     0,     1,     1,     2,    -1,    -2,     1,     2,    -2,     3,     0,     1,     0,    -1,     5,     0,    -2,     0,    -5,    -1,    -4,     1,     1,     1,     0,     0,    -4,    -3,    -3,     0,     4,     1,     1,     1,    -2,     0,    -1,     1,    -2,     0,    -1,     3,     5,     0,    -2,     2,     0,     1,     0,    -4,     0,     4,     0,    -2,    -1,    -2,    -1,    -2,    -2,    -2,    -2,     2,    -1,     0,    -2,    -1,    -2,     3,    -3,     3,     0,     1,     1,     2,     2,     2,    -1,     0,     0,     1,     0,     2,     0,    -2,    -1,    -1,    -5,    -5,    -2,    -2,     0,    -2,     2,     0,     1,    -3,    -3,    -6,     0,     0,     1,     1,     4,     2,     0,     1,    -2,    -2,     0,    -1,     0,    -4,    -2,    -5,    -8,    -2,    -3,     1,     0,    -3,    -2,     1,     1,    -1,    -4,    -7,     0,     1,     0,     1,     1,    -1,    -1,    -3,    -3,    -2,    -1,     0,    -1,    -2,    -6,    -4,    -5,    -4,    -4,    -2,    -7,    -4,    -3,     1,    -3,    -2,    -4,    -6,     0,     0,     0,    -3,    -1,    -4,    -2,    -7,    -4,    -4,    -5,    -6,    -4,    -7,    -8,    -7,    -7,    -5,    -3,    -8,    -8,    -5,    -2,    -1,    -5,     1,     1,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -5,    -6,    -4,    -2,    -4,    -4,    -4,    -4,    -6,    -6,    -4,    -6,    -4,    -2,    -2,     0,     1,     2,     3,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,    -3,    -2,    -1,    -1,     0,    -2,     0,    -1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     1,     0,     1,     0),
		    23 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,    -1,    -3,    -3,     0,     0,    -2,    -2,    -2,    -3,    -5,    -3,    -2,    -3,    -2,    -1,    -1,    -3,     0,     0,     0,     0,     0,     0,    -1,     1,    -1,     2,     3,     5,     2,     1,    -2,     0,     0,     0,    -2,     1,     2,    -1,    -6,    -4,    -1,    -4,    -2,    -4,    -1,    -1,     1,     0,     0,     1,     0,     1,     3,     3,     1,     2,     4,     3,     0,    -1,     1,     1,     1,     0,     0,     0,    -4,    -5,    -7,    -3,    -3,    -6,    -3,    -1,    -1,     0,     1,     0,     2,     0,     1,     2,     2,     0,     0,     0,     2,     2,     1,     3,     0,     1,     1,    -2,    -2,    -1,    -6,    -5,    -7,    -6,    -3,    -2,    -1,    -1,     1,     1,     1,     2,     1,     3,     3,     1,     2,     3,     3,    -1,     0,     1,     0,     1,     1,     1,     1,    -1,    -2,    -6,    -6,    -5,    -1,    -2,    -3,     0,     0,     0,     0,     2,     4,     4,     1,     1,    -1,     0,     0,    -1,    -2,     2,     1,     0,     2,     1,    -1,    -1,    -5,    -6,    -6,    -7,    -3,     0,    -3,    -1,    -1,     0,     1,     1,     0,     3,     3,     2,     0,    -5,    -2,    -8,    -5,    -1,    -1,     1,     2,     0,     0,     3,    -4,    -4,    -6,    -7,    -5,    -1,    -3,     0,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -6,    -9,    -8,    -5,    -5,    -1,    -1,     2,     2,     1,     1,     0,    -4,    -8,    -6,    -5,    -3,    -2,    -2,    -3,     0,     0,    -2,     1,     0,    -4,    -6,   -11,   -11,    -7,    -2,     2,     0,     0,     2,     3,     0,     0,     1,    -4,    -7,    -8,    -7,    -1,     0,    -2,    -1,    -2,    -1,     1,    -1,     0,    -1,    -6,    -7,    -6,    -5,     3,     2,     3,     4,     2,     3,     2,     0,    -4,    -4,    -3,    -5,    -4,    -4,    -3,     0,    -3,    -1,    -2,     0,     0,    -1,    -1,    -2,    -2,     0,    -1,     3,     3,     4,     2,     1,     0,     1,    -1,     1,    -3,    -4,    -2,    -3,    -2,    -3,    -1,    -2,    -3,     0,    -1,    -1,     0,     0,    -1,    -2,     0,     1,     3,     7,     5,     2,     0,    -2,     0,    -1,     3,     0,     0,    -3,    -1,    -1,     0,     0,    -2,    -1,    -3,    -3,    -2,    -1,     0,     0,     0,    -2,     1,    -1,    -1,     0,     1,    -1,    -1,    -2,    -2,     0,     0,    -2,    -1,    -1,    -1,     1,     0,     3,     0,     1,     0,    -6,    -1,    -2,    -1,     2,     0,    -2,     0,     0,    -1,    -5,    -2,    -3,    -2,    -3,    -2,     0,     0,    -4,     0,     2,     0,    -1,     0,     3,     1,     1,     2,    -3,    -1,    -1,     0,     0,     0,    -2,    -2,    -2,    -4,    -6,    -2,    -4,    -4,    -6,    -9,    -5,    -2,    -3,     0,     1,     0,     1,     1,     3,     3,     2,     2,    -7,    -5,    -1,     0,     1,     2,     1,    -2,    -2,    -1,     1,     3,     1,    -1,    -6,    -8,    -6,    -6,    -3,     0,     1,    -3,    -3,    -1,     1,     1,    -3,    -1,    -7,    -1,    -2,    -1,     1,    -1,     3,     2,     2,     5,    -2,     5,     1,    -1,    -1,    -1,    -3,    -2,    -1,     2,    -2,    -2,     0,     0,     0,     0,    -3,    -3,    -3,    -2,    -1,    -1,     0,    -3,     1,     1,     1,    -1,    -1,     2,    -1,    -1,     2,     3,     3,    -1,    -1,    -3,    -1,    -1,     0,    -1,    -2,     0,    -1,     1,    -2,    -3,    -2,     0,     0,    -3,     1,    -2,     1,     1,    -1,     1,     1,     0,    -2,    -2,    -2,     0,    -1,     0,     0,     1,    -2,     0,    -3,    -3,    -1,     1,    -1,    -3,    -1,    -1,     0,     1,     0,     0,     0,     1,     1,     1,     2,     0,     1,     2,     0,    -2,    -2,     0,    -2,     0,     0,    -1,    -3,    -1,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     2,     4,     1,     3,     1,     0,     1,     1,     1,     0,     0,     0,     0,    -2,    -1,    -1,     0,    -1,     0,     1,     1,     1,    -3,     0,     0,     0,     0,     1,     5,     5,     1,     1,     2,     1,     1,     1,     0,    -2,     2,    -1,     0,    -1,    -1,     1,     0,     1,     0,    -2,     0,     2,     0,    -1,     0,     0,     0,    -1,     1,    -1,     0,    -4,     2,    -1,    -2,    -1,     1,     0,     0,     0,    -1,    -2,    -1,    -1,    -2,    -2,    -3,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     1,    -1,    -1,    -1,     2,     3,     3,    -1,    -1,    -3,    -6,    -2,    -3,    -2,     1,     0,     0,     3,    -1,    -3,    -5,    -3,     0,    -1,     0,    -1,     0,     0,     1,    -1,    -1,    -2,    -1,     0,    -2,    -3,    -2,    -2,    -3,    -4,    -5,     0,     1,    -1,    -1,     0,    -2,    -2,    -3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -4,    -2,    -4,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     1,    -1,     0,     0),
		    24 => (    0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -2,    -2,    -1,    -3,    -4,    -2,    -5,    -1,     2,    -2,    -3,    -2,    -3,    -1,    -2,    -1,    -1,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -6,    -6,    -1,    -2,    -4,    -4,    -3,    -4,    -6,    -5,    -2,    -1,    -4,    -3,    -3,    -2,    -4,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     1,     0,    -1,    -5,    -5,     0,    -2,    -5,    -4,    -6,    -1,    -3,    -6,    -4,     0,     0,     2,     2,     2,     0,    -2,     0,     2,     1,     2,    -2,     0,     0,     0,     1,     0,    -1,     1,    -4,    -1,    -2,    -1,     0,    -1,     1,    -1,     1,    -2,     0,     1,     0,    -2,    -3,     2,     2,     5,     5,     3,     0,    -2,    -1,     0,     0,    -1,     1,    -2,    -1,    -2,    -3,    -2,    -2,     0,     2,     1,    -1,    -2,    -2,    -4,    -5,    -2,    -1,     1,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     1,    -2,    -3,    -1,     1,     1,    -2,    -3,    -1,    -2,    -1,    -9,   -11,    -5,     0,     3,     1,     2,     1,    -3,    -1,     0,    -2,     0,    -1,     0,    -2,    -1,    -1,    -2,    -1,     1,     0,     0,     0,     0,     1,    -1,    -6,   -11,    -9,    -3,     2,     1,     3,     5,     4,    -2,    -4,     3,    -2,    -1,    -2,     2,    -1,    -3,    -3,    -2,    -1,    -1,    -3,     0,    -2,    -1,     2,    -2,    -5,    -9,    -7,    -1,     1,     0,     1,     3,     2,    -2,    -1,     2,    -3,     0,    -1,     2,    -2,    -2,    -1,    -1,    -2,     0,     0,    -1,    -2,     1,     1,    -4,    -8,   -10,    -6,    -1,     4,     2,     0,     3,     1,     0,     0,    -2,    -1,     0,     0,     1,     2,    -1,    -2,    -2,    -1,     1,     0,    -1,     1,     1,     0,    -7,    -9,    -6,    -3,     3,     3,     1,    -1,     0,     1,     1,    -1,    -1,    -2,     0,    -1,    -1,     1,    -1,    -2,    -1,    -2,     0,    -1,     1,     1,     0,    -1,    -3,    -6,    -4,    -1,     1,     3,    -1,     0,     0,     1,    -1,    -2,    -2,    -3,     0,     0,     1,    -2,    -1,    -3,    -1,     0,     0,    -1,     0,     0,     1,    -2,    -6,    -3,    -4,    -1,     3,     2,     0,    -2,     0,     1,    -2,    -3,    -2,    -3,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     1,    -1,     0,    -2,     0,    -3,    -3,    -3,    -3,     0,    -1,    -1,    -1,     1,     1,     0,    -5,    -1,    -2,     0,     0,     0,    -3,     4,     1,     5,    -1,     1,    -3,     1,     0,     0,    -2,    -3,    -2,    -2,    -2,     0,    -3,     1,     0,    -1,     0,    -1,    -2,    -4,     0,     0,     0,     1,     6,     3,     1,     2,    -2,     0,     0,     3,     3,     0,    -2,    -1,    -3,    -3,    -3,     1,     0,     0,     0,    -3,     2,    -1,    -6,    -4,    -3,    -1,     0,     1,     2,     0,    -5,    -1,     2,     3,     5,     3,     6,     0,    -2,     0,    -2,    -1,     0,     0,     0,     0,     1,     0,     2,    -4,    -3,    -4,    -2,    -2,    -1,     0,     0,    -3,    -3,    -2,     1,     3,     4,     2,     4,     2,    -2,     0,     1,     0,    -1,     1,     4,     3,     1,     2,     2,     0,    -4,    -3,     1,    -2,    -1,     0,     0,    -6,     1,     1,     0,     1,     1,     0,     0,     0,     2,     0,     1,     2,     1,     2,     3,     2,     1,     2,     1,    -2,    -5,    -3,     0,     0,     0,     0,    -1,    -4,    -1,     2,     3,     0,     0,     0,    -1,    -1,    -2,    -1,     0,     2,     0,     0,     1,     3,     0,    -3,    -2,    -2,     0,    -5,    -1,     0,     0,     0,     0,    -5,    -4,    -1,    -2,    -2,    -3,    -4,    -5,    -4,    -1,    -2,     1,    -1,    -2,    -1,    -2,     3,     1,    -1,     1,     1,     1,    -3,    -2,     0,     0,     0,    -1,    -4,    -1,    -2,    -2,    -1,    -4,    -7,    -7,    -3,    -2,    -1,     0,    -1,     0,     0,     0,     2,     0,    -1,     2,     2,     0,    -4,    -2,     0,    -1,     0,    -1,    -3,    -4,    -2,    -3,    -4,    -5,    -5,    -5,     2,     0,    -2,    -2,    -1,     0,    -2,    -1,     0,    -2,     2,     2,     3,    -2,     0,    -1,     0,     0,    -1,     0,    -1,    -3,    -1,    -3,    -4,    -1,    -1,     0,     2,     1,    -1,     0,    -2,     1,    -1,    -1,    -1,    -4,     2,     0,     1,    -3,    -2,    -1,     0,     0,     0,     0,    -1,    -1,     1,     0,    -3,    -1,     0,     0,    -1,    -1,     0,    -2,     0,     2,     1,    -3,    -2,    -4,     0,     3,     2,    -3,    -2,    -1,     0,    -1,     0,    -1,     1,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,     0,     0,    -4,     0,    -1,    -3,     1,    -1,    -3,    -4,    -1,     1,    -2,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     1,     2,     1,     2,     1,    -7,    -4,    -2,    -2,    -3,    -1,    -4,    -5,    -4,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,     0,    -3,    -3,    -1,    -2,    -1,    -3,    -2,     0,     0,    -1,    -1,     0),
		    25 => (   -1,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -1,    -2,     0,    -2,     3,     2,    -2,     1,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     1,     1,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -4,    -1,     1,     1,     2,     2,    -2,     1,     2,     1,    -2,    -2,    -1,     2,     0,     0,     0,    -1,     1,    -1,     0,     0,     0,    -1,     0,    -2,    -6,    -4,    -4,     0,     2,    -2,     1,     2,     0,    -1,     0,    -1,     1,     1,     1,     0,    -3,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -4,    -5,    -3,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,    -2,    -1,     2,     1,     4,    -1,    -2,     0,     0,     0,    -1,    -1,    -2,     0,    -2,    -1,    -2,    -3,    -7,    -1,    -1,     3,     0,     0,    -2,     0,     2,     1,    -1,     3,     3,     3,     3,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     0,    -2,    -6,    -1,    -5,    -2,    -1,     0,     1,     1,     0,    -1,     0,    -1,     1,     3,     3,     2,     4,     1,     0,    -1,    -2,    -2,    -1,     0,    -1,     1,    -2,    -2,    -2,    -1,     0,     3,     0,    -1,     0,    -2,    -1,     1,     0,    -1,     1,     3,     4,     4,     4,     0,     2,     0,     0,    -2,    -1,     0,     1,    -2,    -2,     0,     0,     2,    -1,     1,    -2,     0,     0,    -2,     0,    -1,    -1,    -1,     0,     3,     4,     7,     4,     0,     3,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,    -4,     2,    -1,     1,     1,     3,     0,    -1,    -2,     1,     2,     2,    -2,     1,     1,     4,     3,     2,     3,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,     2,     0,     0,    -1,    -2,    -2,    -4,    -4,    -3,     1,    -4,    -2,    -1,     1,    -1,     1,     3,     1,     0,     0,     0,     0,    -1,     0,     1,     1,     2,     0,     1,    -1,     1,     2,    -1,    -4,    -8,    -9,    -8,    -9,    -8,    -8,    -5,    -2,    -3,     0,     2,    -3,     0,    -1,     0,     0,    -2,     0,     2,     1,    -1,     0,     1,    -2,     1,     0,     0,    -3,    -5,    -6,    -8,    -7,    -7,    -7,    -7,    -4,     0,     0,     3,    -2,     1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,    -1,     2,    -2,     0,     0,    -1,    -1,    -3,    -7,    -8,    -6,    -6,    -5,    -4,    -3,     1,     1,     0,    -2,     0,    -1,    -1,     0,    -1,    -3,    -3,    -3,     0,    -1,    -1,    -1,     2,    -1,     1,     1,     0,     0,    -4,    -5,    -6,    -5,    -4,    -2,    -1,     0,     0,    -1,     1,    -1,    -1,     2,    -1,    -3,    -5,    -5,    -2,    -2,    -1,    -1,     0,     0,     1,     0,     1,     0,    -3,    -5,    -6,    -4,    -3,    -3,    -1,    -1,    -2,    -1,     0,     0,    -3,     4,     1,    -3,    -5,    -5,    -2,    -3,    -4,    -1,     2,     0,     1,     0,     2,     3,    -3,    -4,    -5,    -3,    -2,    -3,    -3,    -1,    -2,    -2,     0,    -1,     0,     4,     3,     2,     0,    -1,    -3,    -4,    -3,    -3,    -2,     1,    -1,    -1,    -2,    -1,    -3,    -2,    -5,    -3,    -2,    -2,    -1,    -1,    -2,    -1,     0,     0,     1,     0,     3,     2,     3,     4,    -1,    -3,     0,    -2,    -2,     2,    -2,     0,     0,     2,    -3,    -2,    -2,    -1,    -1,    -2,    -1,    -3,    -2,    -1,    -1,     0,     0,     1,    -1,     2,     2,     4,     2,     0,     0,     0,     1,     2,     0,     1,     3,     0,    -1,    -3,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -2,     2,     2,     1,     0,     1,     1,     1,     2,     1,     1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     1,    -1,     2,     0,    -2,     0,     1,     0,     0,     0,     3,     2,     0,     0,     1,    -2,     0,     0,    -2,    -2,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     2,     1,     2,    -1,     0,     4,     3,     3,     1,     3,     2,     1,     1,     0,     0,     2,     0,     0,    -1,     0,     0,     0,     1,    -1,    -2,     0,     0,     0,    -1,    -1,     0,    -2,     1,     2,     0,     4,     3,     3,     2,     1,     0,    -1,    -2,     1,    -1,     1,     0,     0,     0,     0,     0,    -3,    -1,     1,     0,     0,     0,     0,    -3,    -3,     0,    -2,    -1,     2,     0,    -1,    -1,     0,    -3,    -3,    -2,    -1,     2,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -4,    -4,    -2,    -1,     1,     2,     3,     1,    -4,    -4,    -1,     0,    -1,     0,     0,     0,     1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     1,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,     0,    -1,    -1,     0),
		    26 => (    0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     2,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     2,     2,     3,     2,     5,     5,     1,     2,    -2,     0,    -1,     0,     2,     2,     6,     2,     1,     3,     1,     0,     0,    -1,     0,     0,     1,     2,     3,     5,     2,     3,     6,     5,     3,     3,    -5,    -3,     0,     0,     0,     3,     2,     0,     2,     2,     4,     2,     0,    -3,     0,     0,     1,     0,    -5,    -1,     0,     4,     4,     1,     1,     0,    -1,    -3,    -5,    -1,     2,     1,    -1,     2,     2,     1,     0,    -2,     0,     5,     2,    -4,    -3,     0,     0,     0,    -5,     0,     0,     4,     0,    -1,     3,     3,    -1,    -3,    -7,    -2,     0,    -2,     1,    -1,    -3,     0,    -1,     2,     2,     4,     0,    -5,     3,     4,     1,     0,    -4,    -3,     1,    -2,    -5,     2,     2,     1,    -3,    -7,    -3,    -2,     0,     0,    -4,    -1,    -4,    -2,     0,     0,     1,     3,     1,    -2,     6,     4,     0,    -1,     2,    -1,     1,    -2,    -3,     2,    -1,    -4,    -3,    -3,     0,    -3,    -3,     0,    -1,    -1,     0,     1,    -1,    -2,     2,     0,     1,    -2,     2,     2,     0,     0,     0,    -2,     1,    -1,    -2,    -1,    -2,    -3,    -3,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -3,    -1,    -1,     0,     0,     0,     1,     0,     1,     2,     0,     1,    -2,    -2,     1,    -2,    -3,    -3,    -2,    -4,     0,    -1,    -2,    -1,    -3,    -3,    -2,    -3,    -5,     0,    -5,     0,    -1,    -1,     2,    -6,    -1,    -4,     1,     0,    -3,     1,     1,    -5,    -1,    -3,    -3,     0,     0,     1,    -2,    -2,    -1,    -4,    -7,    -6,    -6,    -3,    -4,    -3,    -9,    -3,     1,     0,    -1,    -4,     0,     0,    -4,    -3,    -2,    -4,    -5,    -5,    -3,     1,    -2,    -1,     1,     0,    -2,    -3,    -5,    -4,    -2,    -2,    -2,    -2,    -3,     2,     3,     4,    -3,    -6,     0,     0,     0,    -2,    -1,    -2,    -3,     0,    -1,     1,     2,     1,     1,     3,     1,    -1,    -1,    -2,    -3,    -4,     1,    -2,    -2,     1,     1,    -1,    -3,    -1,     0,     0,    -1,    -2,    -2,    -4,     0,     2,     3,     4,     4,     1,     0,     1,     0,    -1,     1,    -1,    -3,    -6,    -5,    -1,     2,     4,     3,     0,    -5,    -1,     0,     0,    -1,    -2,    -2,     0,     4,     2,     1,     3,     4,     1,     0,    -1,    -1,     0,     0,     0,    -2,    -2,    -3,    -2,     1,     4,     3,     1,    -2,     1,     0,     1,    -1,    -4,    -3,     3,     1,     1,     3,     4,     1,     3,     0,    -2,     0,     0,     1,    -1,    -1,    -1,    -1,     2,     3,     3,     1,     1,    -4,    -3,     0,     0,    -2,    -4,    -4,     3,     3,     4,     6,     5,     3,     2,     2,     1,    -1,    -2,    -1,     0,     0,     1,     1,    -1,     3,     3,    -3,    -2,    -5,    -3,     0,     0,     0,    -4,    -1,     2,     2,     4,     7,     6,     4,     4,     4,     0,     1,     0,     1,    -1,    -1,     3,     2,     1,     2,     3,    -2,    -3,    -5,    -3,     0,    -1,     0,    -4,    -4,     1,     2,     3,     2,     2,     5,     2,     4,     5,     0,     0,    -1,    -1,    -1,     1,     1,     2,     0,    -1,    -1,    -4,    -6,    -4,     1,     0,    -1,     0,    -2,    -1,     0,     2,    -1,     1,     1,     0,     4,     5,     2,    -3,     0,     0,    -2,    -3,     0,    -1,    -1,    -2,    -6,    -4,    -3,    -3,     0,     0,    -3,     0,     0,    -4,    -3,    -1,    -3,     0,    -1,     2,     2,     1,     0,    -1,    -1,     2,    -2,    -1,    -1,     0,    -1,     0,    -3,     1,    -2,    -4,     0,    -1,     0,    -4,     1,    -3,    -3,    -2,    -2,     1,    -1,     0,    -1,    -2,     2,     0,    -3,    -2,     0,    -1,    -1,    -1,     3,     0,     2,     4,    -1,     0,     0,     0,    -1,    -2,    -2,    -2,    -3,    -1,    -1,     1,     0,    -3,     3,     3,     0,    -2,    -1,     0,     0,     2,    -1,     0,     3,     3,     3,     1,    -1,    -1,     0,     0,     0,    -1,    -2,    -6,    -6,    -3,     2,    -2,     0,    -2,     3,     3,     1,     2,     2,     0,     1,     1,    -1,     2,    -1,     0,    -2,    -5,    -1,    -1,     1,     0,     1,    -1,    -3,    -4,    -5,    -4,    -2,    -1,    -1,     0,    -2,     0,    -1,     1,    -2,     0,     2,     3,     0,    -3,    -5,    -4,    -3,    -3,    -5,     0,     1,     0,     0,     0,    -2,    -1,    -1,    -3,    -4,    -5,    -6,    -4,    -1,    -3,     0,     2,     2,     3,     1,    -6,    -3,    -6,    -4,    -3,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -2,    -2,    -3,     0,     3,     0,    -2,    -1,    -3,    -2,    -1,    -2,    -4,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -2,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     1,    -1,     0,     0,     1,    -1,    -1,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0),
		    27 => (    1,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,     0,    -3,    -2,    -2,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,    -3,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -2,    -1,     0,    -1,    -2,    -1,     0,    -2,     0,    -2,    -2,    -1,     0,     0,     1,     0,     0,     0,     0,     0,    -3,     0,    -1,    -3,    -3,    -4,    -5,    -5,    -5,    -5,    -4,    -4,    -3,    -1,    -1,    -1,     0,    -2,    -3,    -3,    -2,    -2,    -1,     0,     0,     0,     0,    -2,     1,     1,    -1,    -3,     2,     2,    -3,    -2,    -4,    -3,    -3,    -4,    -5,   -10,   -12,    -8,    -6,    -2,     0,    -5,    -4,    -4,    -2,     0,     0,     0,     1,     5,     4,     3,    -1,    -3,     3,     0,    -2,     0,     2,     2,     0,    -4,    -1,     0,     2,     0,     1,     5,     0,    -7,    -5,    -5,    -3,     0,     0,     4,     0,     4,     4,    -1,     0,     0,     0,     2,     3,     3,     2,     0,    -1,    -1,     1,     1,     0,     3,     2,     3,     4,     4,     0,    -2,    -4,    -2,    -3,     5,     1,     3,     2,    -3,    -2,     1,     2,     0,     0,     1,     1,     1,     0,     1,     1,    -1,     1,     1,     1,     2,     1,     1,     1,    -3,    -5,    -1,     0,     3,    -2,     1,     2,     1,     0,     2,     2,     3,     3,     2,     3,     0,    -1,     0,    -1,     1,     0,     2,     1,     4,     1,     0,    -1,    -1,    -5,     0,     0,     2,     0,    -2,     3,     3,     0,     1,     1,     1,     1,     3,     1,    -1,    -4,    -2,     0,     3,    -1,     2,     2,     1,     1,    -1,    -3,    -3,    -3,     1,     0,    -1,     4,    -1,     3,     1,     1,     2,     0,     0,     4,     5,    -1,    -6,    -9,    -2,     1,     2,    -1,     0,     2,    -1,    -1,    -1,     1,    -4,    -1,     0,     0,     2,     1,     0,     0,     3,    -2,     2,     0,     0,     2,    -1,    -6,   -14,    -9,    -1,     1,     0,     1,    -4,     0,     1,    -1,    -5,     0,    -2,    -1,     1,     0,     2,     0,     0,    -2,    -1,     1,     2,     2,     2,     1,     0,    -9,   -15,    -6,    -2,     1,     0,    -3,    -4,     0,     1,    -4,    -5,    -2,    -1,    -2,    -1,     0,     0,     2,     0,    -1,    -1,     3,     1,     1,     1,     3,    -5,   -13,   -13,     0,     0,     1,    -1,    -3,    -1,     0,    -2,    -2,     0,     2,    -1,    -1,     0,     0,     0,     2,    -1,    -2,     1,     0,     2,     0,    -1,     0,    -8,   -14,    -3,    -2,    -3,     0,    -1,    -1,     0,     1,    -1,     0,     1,     2,     0,     0,     0,     1,     0,     2,    -2,    -2,     0,    -1,     0,    -1,    -3,    -4,    -8,    -5,    -2,    -2,    -2,    -2,    -1,    -2,    -1,     0,     0,    -1,    -4,    -4,    -2,     0,    -1,     0,     0,     0,    -2,    -2,    -1,    -6,    -3,    -2,    -2,    -2,    -1,    -4,    -4,    -2,    -1,     0,     0,     2,     1,     0,     1,     0,    -4,    -5,    -2,     0,    -3,     1,     0,     3,    -4,    -4,    -1,    -2,    -3,    -3,     0,    -1,    -3,    -4,    -2,    -1,    -3,     0,     1,     1,     1,     0,    -3,    -2,    -3,    -6,    -5,     0,    -2,     1,     2,     0,    -4,     1,     2,    -1,    -5,     2,     2,    -1,     0,    -2,    -1,     1,    -1,    -1,    -2,    -2,    -1,     0,    -3,     1,    -3,    -3,    -2,     0,    -1,     0,     3,    -1,    -1,    -2,    -4,    -4,    -1,     0,     1,     0,    -1,     3,    -1,     0,    -1,    -3,    -2,    -3,     0,    -3,    -6,    -5,    -5,    -4,     0,    -1,     1,     0,     1,     0,    -2,    -4,    -4,    -3,    -5,    -1,    -2,     1,     3,     1,     0,     0,    -1,    -1,    -3,    -1,     0,    -1,     1,     1,    -2,     0,     0,    -2,     0,     0,     0,    -1,    -2,    -3,     1,    -3,    -2,    -1,     0,     0,    -1,    -1,     1,    -1,     1,    -2,    -1,     1,     1,    -2,    -1,    -2,    -2,    -1,     0,    -5,     0,     0,     0,    -1,    -2,     1,     3,     1,     0,    -2,     1,     2,    -2,    -3,     0,    -2,     0,     0,     0,    -2,     0,    -3,     0,    -3,    -2,    -1,     0,    -3,     0,     0,     0,     2,     3,     7,     4,     0,    -1,     0,    -2,     3,    -1,    -1,    -4,    -5,     1,    -1,    -1,    -2,     0,    -2,     1,    -2,    -1,     0,    -1,     0,     0,     0,     1,    -3,     2,     1,    -4,    -3,     0,     1,     0,    -3,    -1,     3,     0,     2,     1,     0,     1,     0,    -1,     1,     4,     2,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -4,    -2,     3,     3,    -1,    -3,    -3,    -2,     1,     0,     2,     1,    -1,     0,     3,     2,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     3,     3,     1,     0,     2,     2,     1,     0,     0,     3,     3,    -1,     0,     3,     1,     2,     2,     1,     1,     4,    -1,     0,     0,     0),
		    28 => (    0,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -5,    -4,    -5,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,     0,    -1,     0,    -2,    -4,    -7,    -6,    -3,    -2,    -1,    -6,    -6,    -5,    -2,    -4,    -2,    -3,    -3,    -3,    -1,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,    -4,    -7,    -9,   -10,   -11,    -7,    -6,    -2,     3,    -2,     0,    -2,    -3,    -7,    -7,    -2,     1,     2,     3,     2,     0,    -1,     0,     0,    -2,    -1,    -4,    -5,    -8,    -4,    -4,    -1,    -2,     0,    -3,    -3,     1,     1,     0,    -1,    -2,    -3,     1,     2,    -3,    -2,    -2,     2,    -3,     3,     0,     0,     0,    -4,    -3,    -3,    -7,     0,     0,     1,     0,    -2,     0,    -1,     0,     2,    -2,    -1,     0,    -4,    -1,    -1,     3,     2,    -1,     5,     4,    -3,     1,     0,     0,    -1,    -6,    -2,    -3,     2,     0,     0,     0,    -1,     1,     1,    -2,    -2,    -1,     1,     0,     2,    -2,     1,     2,     2,     3,     1,    -3,    -3,     0,    -1,    -2,    -1,    -5,     0,     1,     0,     2,     0,    -1,     2,     0,    -1,    -2,    -3,     0,     0,     0,     1,     0,    -3,     2,     4,     1,    -1,    -2,    -4,     1,    -2,    -3,    -4,     0,    -1,    -1,     1,     1,     0,     2,    -1,    -2,    -1,     1,    -2,    -4,    -3,     1,     2,     0,     0,     0,     3,     2,     3,    -2,     2,     2,     0,    -2,    -5,     0,    -4,    -1,    -1,    -1,     2,    -1,    -1,    -1,    -2,    -1,    -3,    -4,    -1,     1,    -3,     2,    -1,    -1,    -1,     3,     3,     0,     2,    -2,    -1,    -1,    -6,    -6,     1,    -1,    -1,     2,     0,     2,    -1,     0,    -1,    -2,     4,     1,    -1,    -2,    -1,     1,     1,     0,     1,     5,     3,    -3,     1,    -1,     0,    -1,    -4,     4,     1,     1,    -1,     0,     1,     0,     0,     0,     1,     2,     4,     4,     0,     0,    -1,    -1,     1,     1,     0,     2,     6,     6,     3,    -3,     0,     0,    -3,     5,     3,     2,    -1,     0,     0,    -3,    -3,     3,     4,     4,     2,     3,     1,     4,    -1,     4,     1,     0,    -4,    -1,     2,     4,     2,    -3,     0,     0,    -2,     6,     0,     1,    -1,     1,    -2,     0,     1,     4,     3,     4,     4,     3,     2,     2,     2,     3,    -1,    -4,     1,    -2,    -4,     0,    -1,     0,     0,     0,    -1,     4,     1,     1,     1,    -2,    -3,    -1,     5,     3,     2,     4,     2,     0,     2,     2,     2,     1,    -4,    -5,    -3,    -2,    -3,     4,    -4,     0,     0,     0,    -1,     0,    -5,    -4,    -1,     1,     1,     3,     4,     3,     2,     4,     3,     1,     2,     2,     0,    -2,    -3,    -4,     1,     1,    -4,     4,    -9,    -3,    -1,    -1,    -1,    -1,    -1,    -1,     1,     1,     1,     2,     5,     1,     4,     0,     1,     1,     4,    -3,    -2,     0,    -3,    -2,    -1,     4,    -5,     2,    -7,    -3,     0,     0,    -1,    -3,     3,     1,     5,    -1,    -2,     2,     4,     5,     4,     5,     3,     0,     4,     0,    -3,    -1,    -2,    -1,     1,     6,     2,    -4,    -2,    -5,    -1,    -1,    -1,    -4,     4,     0,    -1,     1,    -1,     1,     2,     3,     6,     7,     3,     3,    -1,    -2,    -2,    -4,    -1,    -2,    -1,     1,    -1,    -4,    -2,    -2,    -1,     0,    -5,    -2,    -2,     0,     2,    -1,     2,     1,     1,    -2,     1,     4,     1,    -2,    -5,    -3,     0,    -1,     1,    -1,     2,    -2,    -1,    -5,    -7,    -2,     0,     0,    -2,     0,    -1,     0,     2,     1,    -4,    -1,    -2,    -3,    -2,    -2,    -1,    -2,    -1,    -3,     0,    -1,     2,    -2,     2,    -3,    -2,    -4,    -4,     0,    -2,     0,    -3,     1,    -1,     1,     0,    -2,    -3,     0,    -4,    -5,    -4,    -3,    -2,    -3,    -3,     3,     3,    -1,     0,    -1,    -1,    -3,    -6,    -4,    -7,    -1,    -1,    -1,    -2,     0,     1,    -3,    -1,     0,     1,    -1,    -1,    -3,    -2,    -4,    -3,    -1,    -2,    -3,    -1,    -1,    -1,     3,    -2,    -4,    -5,     1,    -3,     0,     0,     0,    -2,     1,     0,     0,    -4,     0,     1,     2,    -2,    -2,    -2,     0,    -3,     0,     0,     0,     0,     2,     4,    -2,     1,     2,    -2,     1,    -4,     0,     1,     1,    -2,    -1,    -7,    -5,    -5,    -6,    -4,     0,     0,    -1,     0,    -1,    -3,    -2,    -3,    -4,    -2,     3,    -1,    -4,    -1,     1,    -2,    -2,    -1,    -1,     0,     0,    -2,    -2,    -1,     0,     3,     2,    -1,     0,     4,     1,    -4,    -2,     0,     2,     2,     0,     1,    -3,    -2,    -3,    -4,    -3,    -4,    -3,    -2,     0,     0,     0,     0,    -2,    -2,    -4,    -5,    -5,    -6,    -9,    -7,    -3,    -3,    -3,    -3,    -9,    -5,    -3,    -4,    -7,    -5,    -3,    -2,    -2,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,    -2,    -4,    -4,    -3,    -1,    -1,    -3,    -4,    -5,    -3,    -3,    -2,    -2,     0,    -1,     0,     0,     0,     0,     0,     0),
		    29 => (    1,     0,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,     0,    -1,    -2,    -3,    -2,    -1,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,     0,     0,    -4,    -3,    -2,    -1,    -1,     0,    -5,    -2,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -4,    -4,    -3,    -4,    -4,    -7,    -8,    -5,    -6,   -11,    -4,    -5,    -8,    -6,    -4,    -6,    -7,    -5,    -3,    -2,    -1,     0,     0,     0,     0,    -2,    -2,    -2,    -7,    -9,    -3,    -4,    -5,    -2,    -2,    -1,    -1,    -2,     1,    -1,    -4,    -1,    -9,    -8,    -2,    -3,    -2,    -1,    -4,    -3,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -3,    -2,     0,     1,     3,     1,     2,     1,    -1,     1,     2,     3,     3,     1,    -4,    -4,    -4,    -1,    -3,    -2,     0,    -1,     0,    -1,    -3,    -2,    -4,    -2,    -3,     0,     3,     1,    -1,    -3,     1,     1,     2,     1,     0,     4,     2,     3,    -1,    -1,     2,     0,    -1,    -2,    -4,     0,    -1,    -3,    -2,    -3,    -3,    -4,    -4,     0,     1,     1,    -1,     0,    -2,     0,    -1,    -1,     0,     0,     1,    -1,    -3,    -3,    -1,     1,     2,    -2,    -1,    -2,    -2,    -1,    -1,    -1,    -3,     1,    -1,     1,     3,     2,    -1,    -1,     0,    -1,    -1,     0,    -1,     0,    -2,    -4,    -3,    -4,    -2,     1,     0,    -3,    -1,     0,    -2,     1,     4,     4,     1,     2,     0,     1,     3,     0,    -1,    -1,    -2,    -2,    -2,     1,     3,     2,    -1,    -1,    -1,    -3,    -5,    -3,    -4,    -7,    -2,     0,    -3,    -3,     2,     8,     4,     4,     3,     1,     1,    -1,    -1,     1,    -1,    -1,     1,     6,     4,     1,    -2,    -2,    -1,    -2,    -2,    -2,     1,    -2,    -1,     0,    -6,     0,     0,     4,     4,     4,     1,    -2,     0,    -1,     1,    -1,     2,     3,     2,     6,     4,     0,    -3,    -2,     0,     2,     1,     0,     3,    -1,    -2,     0,    -1,     1,    -1,     3,     2,     3,    -1,     0,    -1,    -1,     0,     0,     1,     6,     4,     3,     0,     1,    -1,     1,     0,     1,     1,    -2,    -2,    -2,    -2,     0,    -2,    -1,    -2,     2,     4,    -1,     0,    -1,    -2,    -1,     1,     0,     5,     6,     6,     3,     1,     1,    -1,     0,     1,     1,     1,     0,    -1,    -2,    -1,     0,    -2,    -3,    -2,     0,     1,     2,     0,     0,     1,    -1,     1,     2,     6,     6,     4,     4,     1,     2,     2,     2,     0,    -2,    -3,    -2,    -2,     0,     0,     0,     0,    -4,    -2,    -1,    -1,     1,    -1,    -2,    -1,    -1,     0,     2,     6,     6,     3,     4,     1,     4,     2,     3,     1,    -2,    -4,    -4,    -2,     0,    -1,     0,    -1,    -4,    -3,    -1,    -2,     2,     1,     2,    -2,     2,     1,     3,     3,     5,     4,     0,     2,     4,     3,     5,     0,    -1,    -2,    -5,    -4,    -1,    -2,     0,     0,    -4,    -1,    -2,    -3,     3,     3,    -1,     1,     0,     4,     3,     2,     5,     2,     1,     2,     3,     2,     3,     0,    -1,    -2,    -5,    -2,    -3,    -1,     2,     0,    -4,    -2,    -4,    -4,     3,     4,     4,     2,     2,     1,     0,     1,     1,     1,     0,     5,     2,     3,     2,    -1,     0,    -3,    -6,    -3,    -3,    -3,     0,     0,    -5,    -1,    -5,    -4,     2,     4,     3,     3,     2,     1,    -1,     0,    -2,     0,     4,     3,     2,     0,     0,     0,     1,     0,    -2,    -1,    -1,    -1,     0,    -1,    -5,    -2,    -5,    -3,    -2,     1,     3,     1,    -1,     0,     1,    -1,    -2,    -1,     2,     1,     0,     0,    -1,    -1,    -1,     0,    -1,     2,    -2,     0,     0,     0,    -4,    -2,    -4,     0,    -2,     0,    -2,    -1,    -2,     0,     1,    -2,    -2,     2,     0,     0,    -3,    -2,    -1,    -1,    -2,    -1,     1,     0,    -4,     0,     0,     0,    -3,     2,    -2,    -4,    -1,    -2,    -2,    -1,    -1,     0,     1,    -3,    -1,     1,    -3,    -3,    -4,    -2,    -2,    -4,    -3,    -2,     1,    -3,    -1,     0,     0,     0,    -2,     1,    -2,    -2,    -1,    -3,    -3,    -3,    -3,     0,     1,     0,     0,    -2,    -4,    -3,    -3,    -2,     2,    -2,    -3,    -4,     1,    -1,    -2,     0,     0,     0,    -3,    -4,    -1,     1,    -3,    -3,    -1,    -1,    -1,    -1,     0,     0,    -2,    -4,    -3,    -2,    -3,    -3,    -2,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     2,    -1,    -1,    -1,    -3,    -5,    -3,     0,    -2,    -2,     0,    -1,    -1,    -4,     0,    -1,    -1,    -3,    -2,    -2,     0,     2,    -1,     0,    -1,     0,    -1,     0,     0,     4,    -2,    -4,    -3,    -3,    -2,    -2,    -2,     0,     0,     0,     0,    -1,     3,     2,     2,    -3,     0,     1,     0,     1,     1,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     2,     2,     1,     1,     1,     0,     0,     2,     1,    -1,    -1,    -2,     0,     0,    -1,    -2,    -1,    -2,     0,     0,     0,     0),
		    30 => (    1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -3,    -2,    -4,    -2,     2,     1,     1,    -2,     3,     3,     3,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     4,     3,     0,     0,     0,    -2,    -3,    -5,    -6,    -3,    -5,    -4,    -8,    -7,    -7,    -5,    -4,    -3,    -3,    -4,    -3,    -1,    -1,     0,     0,     0,     0,     0,     2,    -1,    -2,    -2,    -4,    -3,    -1,    -4,     1,     2,     3,    -2,    -5,    -2,    -1,    -5,    -6,    -2,    -3,    -3,    -3,    -4,     0,    -2,     0,     0,     0,    -2,    -4,    -1,    -5,     1,     0,    -1,     0,     1,     0,     1,     1,    -2,    -2,    -4,     0,     0,     2,     0,     0,    -2,    -3,    -5,    -6,    -2,     0,    -1,     0,    -1,    -3,    -1,    -1,     2,     1,     0,    -2,     1,    -1,    -3,    -3,    -1,    -2,    -3,    -1,     1,     1,    -2,    -2,     0,    -4,     0,    -8,    -5,    -1,     0,     0,    -1,     0,    -1,     0,     0,     2,     1,    -5,     0,    -2,    -4,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     0,     1,     0,     2,    -6,    -2,     0,     1,    -1,     0,    -2,    -1,    -1,     0,     0,    -3,     0,    -1,     3,    -1,     2,     0,    -2,     1,     0,     2,     3,     1,     3,     2,     4,     1,     0,    -4,     0,     5,    -4,     3,     1,    -2,    -4,    -3,    -2,    -1,     0,     3,     0,     1,     0,     0,     4,     3,     4,     1,     3,     3,     3,     3,     0,     0,    -3,    -6,    -2,     0,     0,     4,    -3,    -3,    -2,    -2,    -3,     0,     1,     1,     0,     0,     0,     2,     1,     2,     2,    -2,     1,     4,     2,    -1,     0,     1,    -5,    -3,    -1,    -1,    -1,     4,     2,    -4,    -2,     2,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,     3,     1,     3,     0,     0,     2,     2,     1,    -3,    -2,    -5,    -6,     0,     0,     4,    -3,    -1,    -7,     0,     1,     1,     1,    -2,    -1,    -3,    -3,     0,    -2,    -2,    -1,    -1,    -2,    -2,     0,     3,     1,    -4,    -5,    -5,    -4,     0,     0,     1,    -3,    -1,    -1,     1,     2,     2,     0,     1,    -1,    -4,    -1,    -1,    -4,    -2,    -1,    -1,    -2,    -1,     0,     2,     3,     0,    -3,    -1,    -2,    -2,     0,     1,     0,     2,     3,     1,     5,     3,     0,     2,     0,    -2,    -1,    -3,    -2,    -4,    -1,     2,     0,     1,    -3,     1,     0,     0,    -3,    -1,    -3,    -3,     0,     0,     0,    -1,     5,     6,     6,     3,     2,     3,     3,     1,     0,    -2,    -3,     0,    -3,     0,     0,     2,    -1,    -4,     0,    -2,     2,    -4,    -5,     0,     0,     0,    -2,    -2,     4,     7,     2,     4,     5,     7,     4,    -1,     3,    -2,    -2,    -1,    -2,     0,     0,    -1,    -1,    -3,     0,     1,     0,    -3,    -6,    -3,     0,     0,    -1,    -5,     4,     4,     3,     3,     5,     6,     2,     5,     3,    -2,     1,     1,    -2,    -1,     0,    -2,    -1,    -3,    -4,     2,    -4,    -6,    -8,     4,     0,     0,    -1,    -6,     2,     2,    -1,     2,     1,     3,     4,     4,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -4,     1,    -1,    -4,    -5,    -4,     6,     0,     0,    -1,    -7,     0,    -1,    -1,     0,     3,     1,     2,     0,     2,     0,     0,     0,    -1,    -2,    -2,    -2,    -2,    -2,     0,    -2,    -2,    -4,    -4,    -2,     0,     2,    -2,    -5,    -2,    -1,    -1,    -1,    -1,    -3,    -2,    -1,     3,     1,     0,     0,    -1,    -3,    -1,     0,    -2,     0,     0,    -2,    -2,    -7,    -4,    -2,     0,     2,    -2,    -6,    -1,     0,    -1,    -2,    -3,    -4,    -1,     1,    -1,     1,     2,     1,     0,    -2,     0,    -2,    -2,    -1,    -1,    -1,    -2,    -6,     0,    -1,     0,     0,    -5,    -3,    -3,    -1,     2,     1,    -2,    -2,    -1,    -1,     1,     4,     3,     3,     3,     1,    -1,    -4,    -3,    -1,     0,    -1,    -2,    -2,     4,     1,     0,     0,    -7,    -2,    -6,    -2,     0,     1,     4,     0,     2,     2,     5,     2,     4,     4,     0,     0,    -2,    -2,     0,     1,     2,     2,    -3,    -2,     2,     1,     0,     0,    -2,    -7,    -5,    -1,     1,    -1,     0,    -1,     1,     1,     1,     1,     2,     1,     2,    -2,    -2,    -2,    -1,     2,    -1,    -2,    -3,    -2,    -5,     0,     0,     0,    -1,    -1,    -1,     2,    -2,    -3,    -4,    -6,    -6,    -4,     1,     4,     4,     4,     3,     0,    -1,    -6,    -4,    -2,    -3,    -4,    -2,     0,     0,     1,     0,     0,     0,    -2,   -10,    -8,    -2,    -1,    -1,    -6,    -5,    -3,     0,    -1,    -2,    -3,    -1,     0,    -4,    -7,    -5,    -5,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -5,    -4,    -6,    -2,    -3,    -5,    -5,    -3,    -3,    -3,    -5,    -4,    -3,    -7,    -7,    -3,    -4,    -5,    -2,    -3,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -1,     0,     0,     0,    -2,     0,     0,    -1,    -1,    -2,    -2,    -1,    -2,    -2,    -2,     0,     0,    -1,     1),
		    31 => (    0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,    -1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,    -2,    -3,    -2,    -2,    -4,     2,    -1,     0,     1,     0,     1,     3,     3,    -6,    -5,    -3,    -1,    -1,     1,    -1,     0,     0,     3,     2,     0,    -3,    -4,     2,     3,     3,     0,    -4,    -2,    -2,     0,     3,     0,     0,     0,     3,     2,    -1,     0,    -2,    -3,    -1,    -1,     0,     0,     0,     3,     3,     2,     3,     0,     0,     2,     1,     2,     0,     0,     2,     0,     0,     0,     3,     4,     3,     0,    -1,     1,     0,    -2,    -3,    -4,    -3,     0,     1,     1,     1,     3,     4,     3,     3,    -1,    -3,    -1,    -1,     0,    -1,    -2,     0,    -1,    -1,     0,     3,     1,    -1,    -1,     2,    -1,    -4,    -3,    -3,     0,    -1,    -3,     1,     4,     3,     4,     2,    -2,    -2,     0,    -1,    -2,    -1,    -2,    -2,     1,     0,     1,     1,     1,    -2,    -2,     0,     0,    -2,    -4,     0,     0,    -2,    -4,    -2,    -6,     0,     3,     4,    -2,    -2,    -2,    -1,     0,     1,     1,     0,     0,    -3,     0,     1,     1,    -1,     0,     2,    -1,    -4,    -8,    -5,     0,    -4,    -5,    -6,    -6,    -2,     1,     0,    -3,    -2,     0,    -1,     3,     3,     3,     0,    -1,    -1,     1,     0,    -2,    -1,     2,     0,    -1,    -3,   -11,    -2,     0,    -1,    -4,    -6,    -5,    -3,    -3,    -1,    -3,    -2,    -1,     1,     4,     4,     3,    -1,     0,    -1,     0,     1,    -2,    -3,     0,    -1,    -3,    -3,    -5,    -3,     0,    -1,    -4,    -2,    -5,    -4,    -4,    -2,    -3,    -4,    -2,    -1,     4,     4,     2,     0,    -1,     1,    -1,    -2,    -2,    -3,    -3,    -4,    -3,    -2,    -2,    -1,     0,     1,     0,    -3,    -3,    -4,    -5,    -5,    -4,    -3,    -4,    -3,     0,     3,     1,     2,    -2,    -1,    -1,    -2,     0,    -2,    -1,    -4,    -4,    -2,    -3,     3,     0,    -1,    -5,    -2,    -1,    -3,    -3,    -6,    -4,    -4,    -2,    -2,     0,     4,    -1,     0,     2,     0,    -1,    -1,     1,    -3,    -3,    -2,    -3,    -1,     0,     3,     0,     0,    -5,     1,    -1,    -4,    -2,    -4,    -3,    -2,    -2,    -3,     0,    -1,     1,     1,     4,     3,     0,    -1,    -1,    -6,    -4,    -4,    -4,     0,     0,     0,    -1,     0,     1,     0,    -2,    -3,    -3,    -2,    -3,    -2,    -3,    -3,     1,    -1,     0,     1,     1,     1,    -1,    -4,    -1,    -4,    -3,    -2,    -3,    -3,    -1,     0,     0,     0,     1,    -2,    -4,    -3,    -4,    -4,    -3,    -1,    -1,     0,     0,     1,     1,     0,     2,     2,     1,    -2,    -4,    -6,    -5,    -4,   -11,    -5,    -3,    -2,     0,     0,     1,    -4,    -4,     0,    -2,    -3,    -2,     1,    -1,    -2,    -1,     1,     0,     0,     2,     0,    -1,    -1,    -3,    -5,    -3,    -2,     1,    -3,    -2,    -3,     1,     0,    -2,    -5,    -2,    -2,    -3,    -5,     1,     0,     2,     2,    -2,    -1,     3,     2,     2,     1,     0,     0,    -1,     1,     1,    -1,     1,    -2,    -3,    -3,     0,     0,     0,    -5,    -3,    -4,    -7,    -5,     0,     2,     2,    -1,    -3,    -2,     1,     4,     3,    -1,     1,    -4,    -2,    -1,    -1,     1,     1,     0,    -2,     0,    -1,     0,    -1,    -6,    -6,     0,     0,     0,     2,     3,     3,    -1,    -2,     1,     1,     1,     1,    -1,    -2,    -4,    -3,     0,     2,     2,     3,     1,    -3,    -1,     0,     0,    -2,    -6,    -1,     3,     4,     5,     1,     3,     3,     0,     2,     2,     1,     1,     1,    -2,     1,    -1,     1,     2,     3,     3,     3,     0,    -1,     0,     2,     1,    -1,     0,    -1,     2,     3,     3,     5,     5,     2,     0,     2,     4,     0,    -2,     1,    -1,     1,     0,     2,     2,     3,     1,     1,     1,    -2,     0,     1,     1,    -2,    -1,    -1,     3,     3,     3,     3,     4,     2,     2,     2,     4,    -4,    -3,    -1,    -1,     1,     2,     3,     2,    -2,    -1,     2,     0,     0,     0,     0,     0,    -1,    -1,    -2,     1,     1,     0,     1,     5,     3,     3,     3,     0,    -3,    -2,    -3,     1,    -1,    -1,     1,     0,    -1,    -3,    -3,    -2,     4,    -1,     0,     0,     1,    -1,    -3,     0,    -1,     0,    -1,     2,     1,    -3,    -1,     0,    -4,    -3,    -3,     1,    -1,    -3,    -1,     2,     0,    -4,    -4,     0,     1,     1,    -1,     0,     0,    -1,    -3,    -5,    -3,    -6,     1,    -3,    -1,    -3,     2,     0,    -3,    -4,    -5,    -6,    -7,    -6,   -10,    -4,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -3,    -7,   -10,   -10,    -7,    -7,     1,     0,    -4,    -4,    -4,    -4,    -3,    -5,    -3,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -4,    -3,     0,    -1,    -3,    -1,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,     1),
		    32 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -4,     0,     1,    -1,    -1,    -3,    -1,    -1,    -2,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,    -1,     1,     1,    -1,     1,    -1,    -1,    -1,    -2,    -2,     1,     0,    -3,    -1,    -1,     0,     0,     1,     1,     0,     0,    -1,     0,    -1,    -2,     2,     1,     1,    -2,    -2,    -3,    -2,    -4,    -5,    -3,    -1,    -5,    -6,    -4,    -1,    -4,    -4,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     2,     3,     4,     3,     3,     2,     0,     1,     1,    -2,    -2,    -1,    -1,    -3,    -1,    -1,    -3,    -3,    -4,    -2,    -1,    -1,    -2,     0,     0,    -1,     1,     1,     1,     0,     1,     1,     1,     2,     2,     1,    -1,    -2,    -3,    -4,    -1,    -1,    -2,    -2,    -2,    -1,    -3,    -2,     0,     0,    -1,    -1,     0,     0,    -2,     2,     2,     2,     4,     0,    -1,     0,     0,     0,    -2,    -1,    -2,    -2,     0,     0,     0,     0,    -2,    -1,    -1,    -3,    -1,    -2,    -1,     0,     0,     0,     0,     4,     4,     1,     4,     2,     4,     0,    -2,     0,     2,    -1,    -3,    -1,    -1,    -2,     0,    -1,    -1,    -1,    -2,    -5,    -3,    -2,    -2,    -1,    -2,     1,     0,     1,     2,     1,     3,     2,     2,     2,     1,    -1,     2,    -1,     2,    -1,    -4,    -2,    -2,    -1,    -1,    -3,     0,    -2,    -4,    -2,    -3,    -1,     0,    -1,     0,    -1,     0,     2,     1,     1,    -1,    -1,    -4,    -2,    -2,    -2,     1,     0,    -1,    -3,    -1,     0,     0,    -1,     1,    -1,    -3,    -2,     1,     0,     0,    -1,     0,    -4,    -2,     0,     2,     0,    -1,    -3,    -3,    -7,    -6,    -3,    -1,     0,    -1,    -1,    -1,    -1,     1,    -2,    -2,     0,    -1,    -1,    -2,     0,     1,    -1,    -2,    -2,    -3,    -2,    -1,    -1,    -1,    -3,    -1,    -2,    -6,    -3,    -2,    -1,     0,    -2,    -1,     0,    -1,    -2,     0,    -1,     0,     0,    -4,    -1,     0,     0,    -1,     0,    -3,    -6,    -4,    -4,    -3,    -3,    -2,    -1,    -2,    -3,    -2,    -3,    -1,    -1,    -2,     0,    -2,    -1,     2,     1,     4,     1,    -1,    -1,     0,     0,     0,    -1,    -1,    -6,    -7,    -6,    -4,    -4,    -3,     0,     0,    -1,    -1,    -4,    -2,    -3,    -2,     0,     1,    -1,     3,     4,     5,     3,     0,    -1,     1,    -1,    -1,    -1,    -3,    -5,    -7,    -5,    -4,    -2,     2,     1,    -1,    -3,     0,    -2,    -3,    -4,    -1,     3,     0,     1,     2,     2,     1,     1,     1,     2,     1,    -2,     2,     2,    -2,    -4,    -4,    -1,     0,     1,     2,     0,     1,     2,     2,     0,    -1,     1,     1,     5,     4,     2,     0,     2,     3,     3,     2,     4,     0,    -1,     2,     0,    -2,    -5,    -1,     0,     0,     0,     1,     0,     1,     0,     0,    -1,    -3,     0,     3,     4,     1,     3,     3,     3,     1,     5,     1,     2,     0,    -1,     3,    -1,    -3,    -1,     1,     2,     1,     3,     0,     0,    -2,    -2,     1,    -1,    -4,     2,     4,    -1,     0,     2,    -1,     0,    -3,     3,     0,     2,     0,     0,     1,     3,    -4,     0,     2,     1,     1,    -1,    -2,    -1,     1,    -2,     0,    -1,     1,     3,     2,    -2,    -3,    -1,    -2,    -1,     1,     4,     1,     5,     0,    -3,    -1,    -1,    -4,     0,     1,     2,     1,    -1,    -2,     0,    -1,     0,    -1,     0,     2,     3,     0,    -2,    -3,    -4,     0,    -2,    -3,     0,     3,     4,    -1,    -2,     0,     0,    -3,     0,     1,     1,     1,    -2,    -3,     0,     0,     2,    -1,     0,     1,    -1,    -1,    -2,    -3,    -3,    -2,    -3,    -4,    -1,     1,     0,     0,     1,     1,     1,    -4,    -2,    -1,    -2,     1,    -1,    -1,     1,     0,     1,     0,     2,     2,     0,     0,    -2,     0,     0,    -2,     0,    -2,    -1,     1,    -1,     0,     0,     0,     2,    -3,    -5,    -2,    -3,    -2,    -2,    -1,     2,     0,     3,     3,     0,     0,     1,     0,    -1,     1,     0,    -3,     0,     0,     0,    -2,     0,     0,     0,     0,     2,    -3,    -4,    -3,    -2,    -2,     0,     1,     1,     4,     2,     0,     0,     1,     2,    -1,    -1,    -1,    -1,     1,     1,     1,     1,    -2,     0,     0,     0,    -3,    -2,    -5,    -3,    -4,    -2,    -3,    -4,    -4,    -3,    -3,    -3,    -1,    -1,    -4,    -1,     0,     1,     1,    -1,     0,     1,     2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -2,    -4,    -6,    -5,    -4,    -8,    -1,     0,    -2,     0,    -1,     2,     2,     1,    -2,     0,     1,     1,     0,     0,     0,    -1,     0,     0,     0,    -2,    -2,    -2,    -2,    -4,    -1,    -1,    -2,    -2,    -3,    -2,    -3,    -4,    -3,    -2,    -2,    -1,    -2,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,     0,     1,     0,     0,     1),
		    33 => (    0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -2,    -2,    -4,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -2,    -2,    -1,     0,     0,     0,     0,     0,     2,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,    -2,    -1,    -1,    -1,     0,     0,    -4,    -2,    -1,     0,     0,     0,     0,     1,     2,     0,     1,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -1,     0,     2,     2,     1,     0,    -1,    -2,    -1,    -1,    -3,    -1,     0,     0,     0,     2,    -1,     2,     1,     1,     1,     0,     0,     1,     0,     1,    -1,    -1,    -1,    -2,    -3,     0,     1,    -1,    -3,    -2,    -1,     0,     0,    -2,     0,     0,     1,     3,     0,    -1,     1,     0,     2,     2,     2,     0,     1,     0,    -2,    -1,    -2,    -2,    -1,    -2,    -4,    -2,    -2,    -2,    -2,    -1,    -1,    -3,    -1,    -1,     1,     2,     2,     1,     0,     2,     2,     2,    -1,     1,    -1,    -2,     0,     1,     1,     0,     1,     0,     0,    -2,    -1,    -1,     0,    -1,    -2,    -3,     0,     0,    -3,     5,     1,     2,     0,     3,     1,     0,     2,     1,    -2,    -2,     0,     2,     0,    -4,     0,     1,     0,     0,     1,    -1,     0,    -3,    -3,    -1,     0,     1,    -2,     5,     1,    -1,    -1,     1,     0,    -2,    -3,    -2,    -2,     0,     0,     3,    -3,    -3,    -1,     1,    -1,     1,     1,     0,     0,    -3,    -1,     0,     0,     0,     0,    -2,    -2,    -1,    -2,    -3,    -3,    -3,    -4,    -1,     0,     1,    -1,    -2,    -2,    -1,     0,     1,     0,     1,     1,     1,    -1,    -1,    -3,    -1,     0,     1,     0,    -2,    -1,    -1,    -3,    -4,     0,    -1,    -1,    -1,     0,    -1,    -4,    -2,     0,     0,     1,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -2,    -1,     0,    -2,    -2,     0,     0,     1,    -1,     0,    -1,     1,    -1,    -1,    -1,     1,    -1,    -1,    -2,     0,     1,    -1,    -2,    -1,    -2,    -1,     0,     2,    -1,    -1,     0,     0,    -1,    -2,    -1,    -2,     0,    -1,    -2,     1,     2,     1,     0,    -2,    -3,    -2,    -2,    -1,    -1,     0,    -1,    -4,    -2,    -1,     0,     1,    -1,    -1,     1,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     1,     1,    -1,     0,     0,    -2,    -3,    -1,    -1,     1,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     2,     0,    -1,    -1,     0,     0,    -1,     0,    -2,     0,     0,    -1,     0,     1,     0,    -1,     0,    -2,    -2,    -1,     1,    -1,     2,     0,    -1,     0,    -1,     0,     2,     0,     1,     1,    -1,    -1,     0,    -1,    -3,    -3,    -1,    -1,     0,     1,     0,    -2,    -1,     0,    -1,    -1,     0,     0,     2,     2,     1,     0,    -2,     0,     1,     3,     0,     0,     2,     0,    -1,    -1,    -3,    -3,    -1,     0,     1,     2,     1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     2,     1,     0,    -1,    -1,     0,     1,    -1,     1,     0,    -1,    -1,    -2,    -2,    -2,    -1,     1,     1,     3,     2,    -2,    -1,    -1,    -1,     0,     0,    -1,     1,     1,     1,     1,    -1,    -2,     0,     0,    -3,     0,     2,     0,    -2,     0,    -1,    -2,     0,    -1,     1,     3,     2,    -2,    -2,     0,    -1,     0,     0,     0,     1,     1,     0,     0,    -2,    -3,    -1,    -2,    -3,    -3,    -2,    -3,    -1,     1,    -1,     0,     0,     0,     0,     0,     2,    -2,    -2,     0,     0,    -1,     0,     0,     1,     2,     1,     0,    -1,    -3,    -2,    -1,    -3,    -5,    -3,    -4,    -3,    -1,    -1,     2,     3,     1,    -1,     0,     2,    -1,    -2,     0,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -1,    -1,    -2,    -2,    -3,     0,     2,     1,     1,    -1,     0,     1,     1,     0,    -1,    -2,     1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     1,    -2,    -2,    -3,    -1,    -4,    -1,     2,     4,     2,     0,    -1,    -1,     0,    -1,    -1,     1,    -2,    -1,    -1,     0,     0,     0,     1,    -1,    -3,    -3,    -1,     0,     2,     0,    -1,    -1,     1,     4,     6,     1,     2,    -1,     0,     0,     1,     0,    -2,    -6,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -2,    -4,    -3,    -2,    -4,    -2,    -2,     2,     4,     3,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -3,     1,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,    -1,     1,     0,    -2,    -2,    -1,    -1,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0),
		    34 => (    0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -2,    -2,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,    -2,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -2,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -3,    -1,    -2,    -1,     0,    -1,    -1,    -2,    -4,    -4,    -2,     1,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -4,    -2,    -1,    -1,    -3,    -3,    -1,    -2,    -2,    -1,     1,     0,    -1,    -1,     0,     1,     0,    -1,    -1,     0,    -1,     0,    -2,    -2,    -1,    -3,    -4,    -2,     0,     2,    -1,    -5,    -5,     0,    -2,    -1,    -1,     2,     2,     0,    -2,     0,     0,     0,     0,    -2,    -1,     2,    -2,     0,    -2,    -1,    -2,    -2,    -1,     0,     4,     0,    -8,    -9,    -3,     0,     3,     0,     2,    -2,     1,    -1,     2,    -3,    -1,    -3,     0,     0,    -1,     3,    -1,     0,     0,    -1,    -4,    -2,     2,     1,     1,    -6,    -8,    -6,    -1,     2,     1,     0,     2,     1,     1,     1,     0,    -2,    -1,    -3,     1,    -1,     0,     0,     0,     2,     0,    -1,    -4,     1,     2,     2,    -3,    -3,    -7,    -2,     0,     0,     1,     0,     2,     1,     1,     0,    -1,    -3,     0,    -3,     1,    -1,     0,    -1,    -2,    -1,    -2,    -3,    -2,     3,     0,     0,    -2,    -6,    -5,    -1,     1,     2,     1,     0,     1,     0,     0,    -1,     0,    -1,    -1,     0,    -2,     0,     0,    -3,    -3,    -1,    -3,    -3,    -1,     3,     0,    -2,    -4,    -2,    -1,    -1,    -1,     0,    -1,    -3,    -4,     0,    -3,     0,    -1,    -1,     0,     0,    -2,    -1,    -2,    -2,    -1,    -3,    -1,    -1,     1,     2,     0,    -2,     0,     2,    -1,     0,     0,     2,    -1,    -1,    -2,    -3,    -2,    -1,    -2,    -3,     1,     0,    -4,    -2,    -4,    -2,    -3,    -2,    -2,     0,     1,    -1,     0,     0,     1,    -1,     0,    -1,    -1,     0,    -1,     1,    -1,    -3,    -2,    -2,    -5,    -3,    -1,     0,    -3,    -2,    -4,    -2,     0,    -1,     0,     0,     4,     1,    -1,     1,     2,     2,     2,    -1,    -2,     1,     2,     1,    -3,    -3,    -3,    -4,    -5,    -1,     0,     0,    -2,    -4,    -4,    -1,    -2,    -1,    -2,     0,     1,     0,    -1,     1,     0,     2,     2,    -2,     0,     1,     3,     1,    -2,    -1,    -2,    -2,    -2,     0,     0,     0,    -1,    -1,     1,    -2,    -2,     0,    -1,     1,    -1,    -1,    -1,     0,     0,     3,    -2,     0,    -1,     3,    -2,     0,     0,     1,    -2,    -1,    -1,     1,    -1,     0,    -1,     0,     0,     1,    -2,     0,     1,     2,    -2,    -2,    -1,     1,     0,     0,    -1,    -3,    -4,    -2,    -2,    -2,    -1,     1,     1,     0,    -1,    -1,     1,     0,    -2,     0,    -1,    -2,     0,    -1,     1,    -1,    -2,    -1,    -2,    -2,    -1,     0,     1,    -3,    -3,    -3,    -2,     0,    -1,     1,     0,     0,     0,    -1,    -1,     0,    -2,     1,     2,     0,    -1,     0,    -3,    -4,    -3,     0,    -1,    -1,     0,    -1,     0,    -3,     0,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,    -2,    -3,     1,     2,    -1,    -3,    -3,    -3,    -2,    -3,     0,     0,    -1,    -1,     0,     0,    -2,     0,     1,     0,    -1,    -2,     0,     0,     1,     0,    -1,     0,    -1,     0,    -1,     0,    -2,    -5,    -3,    -5,    -2,    -1,     1,    -2,    -2,    -2,    -4,    -1,    -3,    -1,    -1,    -2,    -2,     0,     1,     1,    -1,    -1,     0,     0,     0,    -1,    -2,     0,    -2,    -6,    -4,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -4,    -2,     0,     0,    -1,    -2,     1,     1,     1,    -3,    -1,     0,    -1,     1,     0,    -2,    -2,     0,    -2,    -3,     0,     0,     1,     2,     0,    -1,    -3,    -1,    -2,    -1,     1,    -2,    -1,     0,     1,     0,     1,     0,     0,    -1,     0,     1,    -1,    -1,    -1,    -3,    -2,    -2,     1,    -1,     1,     0,    -2,    -4,    -2,    -1,    -1,    -1,     3,     2,    -3,     0,     0,     2,     1,     1,     0,     0,     0,     0,     0,    -1,    -3,    -1,     0,    -1,     1,     1,     2,     1,    -3,     0,    -1,     1,     0,    -1,     3,     3,     2,     1,     2,     1,     0,     3,     0,     1,     0,     0,    -2,     0,    -2,    -1,    -3,    -1,    -3,    -2,     1,     0,     1,     1,     0,    -1,    -2,     0,     2,     3,     1,     0,     2,     1,     1,     0,    -1,     1,     0,     0,     0,    -1,    -2,     0,    -2,    -2,    -2,    -3,     0,    -1,     1,    -1,    -3,    -1,     0,    -1,    -3,    -1,    -2,    -5,    -4,     0,    -1,     0,     0,    -1,     0,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -4,    -4,    -3,    -2,    -3,     0,    -2,    -3,    -1,    -2,    -2,    -1,    -1,    -1,    -1,     0,     0,     0),
		    35 => (    1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,     0,    -2,    -1,    -1,    -3,    -3,    -2,    -3,    -3,    -7,    -5,    -3,    -2,    -1,     1,     0,    -3,    -1,     1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -3,    -3,    -2,    -5,    -5,    -4,    -1,    -1,     0,    -1,    -1,    -2,     1,     3,     1,    -2,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0,    -1,     1,    -2,    -1,    -3,     0,    -1,     0,     2,    -1,    -3,    -1,     2,     2,    -1,    -2,     0,    -2,    -2,    -1,    -3,    -4,    -4,    -3,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,    -2,    -4,    -3,    -2,    -2,    -1,    -3,    -3,    -1,    -3,    -3,    -5,    -6,    -1,     1,    -2,    -2,    -1,    -3,    -4,     1,     1,     0,     0,     2,    -3,    -3,     2,    -2,    -2,    -1,    -2,     1,    -1,    -3,    -1,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,     0,    -1,     0,    -4,    -1,     0,     0,    -1,     2,    -2,    -4,     1,    -3,    -2,    -1,    -1,     4,     1,    -1,     0,     0,     1,    -3,    -3,    -5,    -5,    -2,    -1,     0,     1,    -2,    -1,     0,     2,    -1,     0,    -3,     0,    -1,    -1,    -2,     0,     0,     0,     1,     1,    -1,    -1,     1,     1,     2,     1,     0,     2,     2,     2,     3,     3,     3,     2,    -2,     1,     0,     0,    -3,    -2,    -1,    -4,     1,     2,     0,     0,    -1,    -2,    -1,     0,     2,     1,     3,     5,     4,     5,     3,     4,     3,     2,     5,     4,    -3,     1,     0,     0,    -1,    -2,     0,    -1,     1,     1,    -1,     0,     0,     2,    -1,     0,     1,     1,     0,     2,     5,     4,     4,     5,     3,     2,     6,     4,     2,     3,     1,    -1,     0,    -1,     1,     0,    -1,    -3,    -1,    -2,     1,    -1,    -1,    -2,    -4,    -4,    -3,    -3,    -2,    -4,    -3,     1,     1,     2,     1,     5,     4,     0,     0,    -1,     0,     1,    -1,    -2,    -2,    -1,     0,     2,     2,     3,     2,     0,    -2,    -3,    -5,    -4,    -9,   -14,    -9,    -6,    -6,    -3,    -3,     3,     4,    -1,     0,     0,    -1,     1,    -1,    -3,    -3,     1,     0,    -1,     4,     1,     2,     0,     1,     0,    -2,     0,    -3,    -6,    -8,    -5,    -7,    -7,    -2,    -1,     3,    -1,     1,     0,    -1,    -1,     2,     0,     1,     1,     2,     2,     0,     0,     0,     0,    -1,     0,    -1,     1,     0,    -5,    -5,    -4,    -3,    -2,    -2,    -3,    -1,    -1,     1,     0,    -3,     2,     4,     2,     1,     3,     2,     2,    -1,     0,     1,     0,    -2,    -2,    -4,    -1,     1,     0,    -2,    -2,    -4,    -2,    -3,     1,    -1,    -2,     0,     0,    -2,     0,     2,     4,    -1,     2,     0,     1,     0,    -2,    -1,    -1,    -4,    -1,    -2,    -1,     1,     0,     0,    -2,    -1,    -2,    -1,     1,    -2,    -2,     0,    -1,    -4,     1,     1,     1,     1,    -2,    -1,     1,     0,    -1,    -3,    -3,    -3,     0,    -1,     0,    -2,     0,    -1,    -3,    -1,    -1,    -4,    -5,    -4,    -4,    -1,    -1,    -2,    -5,    -2,    -1,     0,    -1,    -1,    -2,    -5,     2,     2,    -1,    -2,     1,    -2,     0,    -1,     0,     1,    -3,    -1,     2,     0,    -2,    -5,    -3,     0,     0,    -1,    -4,     2,     3,    -1,    -2,    -1,    -3,    -4,    -4,     0,     2,    -3,    -2,    -1,     1,     1,     2,     0,    -3,     1,     4,     4,     4,    -4,    -3,     0,     0,    -1,    -3,     2,     0,    -2,     0,    -2,    -2,    -2,     0,     1,     2,    -5,    -2,     1,     0,     0,     2,     1,    -2,     1,     1,     5,     5,    -3,     0,     0,     0,    -1,    -2,    -1,     1,    -2,    -2,    -1,     0,     1,     1,     1,     1,    -2,     3,    -1,     0,    -1,     0,     1,    -1,    -2,     0,     3,     6,     3,    -1,     0,     0,    -2,     0,    -1,     1,     1,    -2,    -3,     0,     0,     1,     2,     1,     0,     2,     1,     2,     0,    -2,     0,     0,    -2,     4,     7,     7,     7,     1,    -1,     0,     2,     0,     0,     0,    -1,    -3,    -3,     2,     3,    -1,     0,    -2,     1,     1,    -1,     0,     0,    -2,     0,    -2,     0,     6,     7,     6,     8,     0,     1,    -1,     0,     0,    -3,    -4,    -3,    -2,    -1,    -2,     0,     1,     2,    -1,     2,    -1,    -1,    -1,    -2,    -1,     0,     2,     4,     2,     2,    -5,    -2,     0,     0,     0,     0,     0,    -4,    -5,    -3,    -4,    -3,    -2,    -2,     0,     4,     2,    -1,    -3,    -2,    -2,     1,     0,    -2,     2,     3,     3,     4,     0,    -1,     0,     0,     0,     0,     0,    -2,    -5,    -7,    -7,    -6,    -6,    -5,    -4,    -4,    -6,    -9,    -2,     0,    -1,    -1,     1,     0,     1,     0,    -3,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -5,    -3,    -1,    -2,    -3,    -2,    -1,    -2,    -5,    -3,     0,     0,     0,     0),
		    36 => (    0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     2,     2,     2,     1,     3,     0,     0,     1,    -2,     0,     0,     1,     3,     2,     5,     2,     2,     2,     1,     0,     0,     0,     0,     0,     2,     1,     3,     2,     3,     3,     2,    -1,    -2,    -2,    -3,    -3,     0,     1,     2,     5,     2,     1,     1,     5,     5,     3,     2,     3,    -1,     0,     0,     0,    -4,     1,    -1,     2,     3,     3,     0,    -1,    -2,    -5,    -6,     0,     3,     2,    -2,    -2,     1,    -2,    -1,     0,    -2,     1,    -4,    -2,    -3,     0,     0,     0,    -5,    -1,     2,     4,     3,    -1,    -3,    -3,    -4,    -6,    -8,    -3,    -4,    -2,     0,    -2,    -1,     5,     4,     1,    -4,    -5,    -8,    -6,    -2,     2,     0,     0,    -2,    -3,     1,     3,     1,    -1,    -2,    -1,    -2,    -7,    -5,     0,     1,    -2,    -1,     0,     2,     2,     3,     2,    -1,     0,    -4,    -5,     0,     0,    -1,     0,     2,     1,     1,     3,     3,     0,    -1,    -4,    -4,    -3,    -2,    -2,    -2,     3,     2,     1,     0,     0,     0,     0,     1,    -2,    -2,    -4,    -2,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -2,    -4,    -7,    -5,    -2,    -2,     1,     2,    -2,    -3,    -1,    -5,     0,    -1,     2,    -3,    -6,    -6,    -1,    -2,     0,     0,    -2,    -2,    -1,     1,     2,    -2,    -4,    -7,    -7,    -1,     0,    -1,    -1,     1,     0,    -2,    -6,     0,    -2,    -3,    -3,    -7,    -6,    -3,    -2,    -3,     0,     0,    -2,    -2,     3,    -1,    -1,     0,    -4,    -4,    -2,     0,    -1,     1,     2,     1,    -3,    -4,    -6,    -8,    -9,    -9,    -8,    -7,    -6,    -3,    -3,    -1,     1,     0,    -2,    -1,    -2,    -2,    -3,    -3,    -6,    -2,     1,     0,     1,     1,     0,    -1,    -3,    -1,    -1,    -5,    -5,    -5,    -7,    -7,    -5,    -4,    -3,    -2,     0,     0,     1,    -4,    -2,    -1,    -1,    -1,     1,     0,     1,     1,     2,     2,    -1,    -4,    -3,    -1,    -2,    -1,    -1,    -3,     0,    -6,    -7,    -6,    -4,    -3,     1,     0,    -1,    -3,    -2,    -1,     0,    -2,     0,     1,     2,     2,     1,     4,    -1,     0,    -3,     2,    -1,     0,    -1,    -2,     1,     1,    -3,    -6,    -6,    -3,     0,     0,    -1,    -3,    -3,    -1,    -2,    -3,     1,     0,     1,     4,     1,     2,     0,     0,    -1,     1,     4,     0,     1,     0,     4,     4,    -3,    -7,    -3,     0,     0,     0,     0,    -4,    -3,     1,    -3,     0,    -1,     2,     2,     1,     0,    -1,    -1,     0,     0,    -5,     1,     2,     0,     4,     3,     0,     1,    -2,    -3,     0,     0,     1,     0,    -3,     0,     1,    -2,     0,     2,     1,     1,    -3,    -1,    -1,     0,    -4,    -3,    -4,     1,     3,     1,     4,     2,     1,    -3,    -4,    -5,    -3,     0,     0,     0,    -1,    -1,     1,     0,     2,    -1,     2,     0,     2,     3,     2,     2,     0,     1,     0,     0,     0,     2,     4,     2,     0,    -4,    -5,    -5,    -4,     0,     0,     0,     0,     1,     1,     0,     1,     3,     0,     1,     2,    -2,     0,    -1,    -2,    -2,    -1,     0,     0,     1,     3,    -1,    -1,    -4,    -3,     0,    -4,     0,    -1,     0,     0,     3,    -1,    -2,    -1,    -1,     3,     2,    -2,    -1,    -1,     0,     3,    -1,     1,     2,     1,     1,    -1,    -6,    -5,    -4,    -3,    -1,    -2,     0,    -1,    -2,     1,     2,    -2,    -1,     0,    -2,     1,     1,     3,     0,    -5,    -2,     1,     0,    -1,     2,    -1,    -1,    -2,    -6,    -3,    -1,    -1,    -2,    -1,     0,    -2,    -1,    -4,     3,     1,    -1,    -1,    -1,    -2,     1,     2,     2,    -1,     0,    -1,    -4,    -2,    -3,    -1,     0,     0,    -1,    -3,    -2,    -2,    -3,     0,     0,     0,    -2,    -2,    -2,    -2,     0,    -1,     0,     0,    -1,     3,    -1,    -1,    -1,    -3,    -1,    -2,    -1,    -2,    -1,     0,    -3,    -2,    -2,    -2,    -2,    -1,     0,     0,    -1,    -1,    -3,    -3,    -4,    -2,    -2,    -1,     0,     0,     1,     2,     0,     1,    -1,    -3,    -1,    -2,    -4,    -4,    -1,    -2,    -5,    -2,     0,    -1,     0,     0,     0,    -1,    -2,    -2,    -2,    -4,    -3,    -4,     0,     2,     1,     0,     1,     2,    -2,    -5,     2,     4,     2,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     1,    -1,     0,     0,    -2,    -3,    -4,    -4,    -5,    -2,    -1,     1,     3,     4,     0,     0,    -5,    -3,    -1,    -1,     0,     0,     0,     1,     1,     0,     0,     1,     1,     1,     0,    -1,    -2,    -1,    -1,    -2,     1,     3,     1,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,     0,     0,    -1,     1,     0,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0),
		    37 => (    0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -3,    -2,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     1,     0,     0,     1,    -1,     0,    -1,     0,     0,    -2,    -2,     0,     0,    -2,    -3,    -1,     0,    -3,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,    -1,    -1,    -1,    -1,    -2,    -5,    -4,    -1,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -3,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -3,    -2,    -2,    -3,    -5,    -5,    -5,    -5,    -5,    -3,    -5,    -4,    -3,    -2,    -3,    -1,    -1,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -4,    -6,     1,    -2,     2,     5,     2,    -3,    -5,    -3,     2,    -2,    -1,    -6,    -7,    -5,    -7,    -6,    -3,    -3,    -3,    -1,    -3,     0,     0,     0,     0,     1,     1,    -1,     0,     0,    -2,     0,    -1,    -4,    -2,    -3,    -3,    -1,    -2,    -5,     0,     1,     0,     0,     3,     0,    -3,    -4,     0,    -4,    -1,     0,     1,     1,     2,     2,     1,     2,     2,     0,     0,     1,    -3,    -2,    -1,    -2,    -4,    -3,    -1,     0,    -6,    -4,    -1,    -1,    -2,    -4,    -2,    -2,    -1,    -1,     1,    -2,     0,     2,     2,     4,     1,     0,     3,     0,     1,     1,     0,    -3,    -2,    -2,    -1,     2,    -3,    -1,     0,    -1,     1,     0,    -2,    -4,    -1,     0,     1,     0,     1,     5,     0,     1,     0,    -1,     1,    -2,     1,     3,     2,     3,     2,    -2,    -2,     0,    -1,     0,     3,     2,     4,     1,    -3,    -2,     3,     0,     3,     2,     2,     6,     2,     3,    -2,     0,     2,     0,     2,     1,     0,     2,     2,    -1,     0,    -1,     0,    -1,    -1,     5,     2,    -4,     0,    -2,     3,     0,     2,     5,     4,     5,     1,    -2,     0,    -1,     0,     1,     2,     0,     1,     1,     1,    -2,    -2,    -1,     0,    -2,     2,     2,    -1,    -6,    -5,    -1,     4,     1,     1,     1,     5,     2,     1,    -1,    -1,    -1,    -1,    -1,     1,     0,    -1,     1,     1,     0,    -2,     1,     1,     0,     2,     3,    -3,    -3,     1,    -1,     3,     1,     2,     2,     5,     2,     1,    -2,    -1,    -3,    -2,     2,     1,    -1,    -3,     1,    -2,     0,    -1,    -1,    -1,     4,     3,     1,    -1,     0,     3,    -2,    -2,    -1,     1,     5,     5,     0,     2,    -2,    -3,    -2,     0,     2,     2,    -2,    -6,    -1,    -1,     0,     2,     0,     3,     2,     2,     1,     4,     4,    -2,    -2,    -1,     0,     1,     3,     3,    -2,     0,     1,     0,    -1,     0,     2,     0,    -3,    -4,     0,    -2,    -2,     1,     1,     4,     2,     1,     3,     2,     2,    -3,    -1,    -1,     0,     0,     1,     1,     4,     1,    -1,     1,     1,     4,     0,    -1,    -6,    -3,    -2,     0,    -1,     0,     0,     2,     0,     4,     5,     5,     2,    -7,    -3,     0,    -1,     0,    -1,     0,     2,     1,    -2,     0,     2,     1,    -2,    -3,    -5,    -4,     1,     1,     1,    -1,     0,    -1,     1,     2,     5,     3,     0,    -7,    -2,    -5,     2,     0,     2,    -5,     0,     0,    -2,     1,     2,     1,    -2,    -4,   -10,    -4,     3,     2,     1,     0,     0,    -2,     1,     1,     3,    -1,    -4,    -2,     0,    -2,     0,     2,    -1,    -5,    -1,     1,     2,     1,     0,    -1,    -6,   -11,    -9,    -3,     3,     0,    -2,     1,    -2,    -1,    -2,    -5,    -7,    -4,    -3,    -3,     0,     0,     0,     1,     0,    -1,     1,     3,     2,     2,     0,    -6,    -8,   -11,    -3,    -1,     0,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -5,    -5,    -1,    -2,     0,     0,     0,     0,    -1,    -1,    -3,     2,     1,     1,    -3,    -6,    -7,    -6,     0,    -3,     1,     2,     2,    -2,    -2,    -2,    -3,    -2,    -3,    -4,    -4,    -2,     0,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,    -4,    -4,    -6,    -3,    -1,    -1,     1,     0,     0,     0,     1,     1,     1,    -1,    -2,    -3,    -2,    -2,    -3,     0,    -1,     0,    -1,    -1,     1,     1,    -1,    -2,    -4,    -4,    -5,    -3,     1,    -1,     3,     1,     0,     0,     3,     0,     0,    -2,    -3,    -4,     0,    -1,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,    -2,    -3,    -3,    -4,    -2,     1,    -1,     0,    -1,    -1,     1,     1,     2,     0,     0,    -1,    -4,     0,     0,    -1,     1,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -2,    -3,    -5,    -3,    -3,    -2,     2,    -1,     2,     2,     2,     2,     1,     0,     1,    -5,     0,    -2,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     1,     1,     1,    -1,    -5,    -3,    -2,    -5,    -2,     2,     1,     2,     3,     1,     1,     1,    -1,    -1,     1,     0,     0,     0,    -1,    -1,     0,     0,     2,    -2,    -2,     0,     3,     2,     0,    -1,    -3,    -4,    -2,     2,     3,     1,    -3,     0,     3,     2,     3,     0,     0,     0,     0),
		    38 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,    -1,     0,     0,     0,     1,    -1,    -1,    -2,    -3,    -1,    -1,     0,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,     0,    -1,     0,    -1,    -1,    -2,    -1,     0,    -2,    -2,    -3,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -3,    -3,     0,     0,    -2,    -2,    -2,     0,     2,     2,     2,     1,    -1,    -1,    -1,     0,     0,     0,     0,    -2,     0,     0,    -1,     1,    -1,    -4,    -2,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,     1,     1,     0,     1,     1,     2,     2,    -2,    -1,    -4,    -2,    -1,    -1,    -1,     0,    -1,    -3,    -3,    -1,     0,    -1,    -2,    -2,    -2,    -2,    -3,    -3,    -2,     1,    -1,    -1,     1,     2,     2,     0,     0,    -2,    -1,     0,     0,    -2,     0,     0,    -1,    -2,     0,     1,    -1,    -1,    -1,    -3,    -4,    -4,    -3,    -2,     0,     1,     0,     0,    -1,     2,    -1,     2,     0,     0,    -2,    -1,     0,     0,     0,    -2,    -2,    -1,     1,     0,     0,     0,     1,     0,     1,    -1,    -1,     2,     1,     1,     0,    -2,    -1,     0,     0,    -2,     0,    -1,    -2,     1,     2,     1,    -1,    -1,    -1,     0,     0,     0,     0,     1,    -1,     1,     1,     0,     0,     0,     3,     3,     1,     0,    -2,     0,    -2,    -1,    -2,    -1,     2,     5,     3,     1,     1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -3,    -2,     0,    -2,    -1,     0,     1,     2,     0,    -2,    -3,     0,    -1,     0,     1,     3,     3,     3,     1,    -4,     0,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,     1,    -2,    -3,    -3,    -2,     0,    -1,    -1,    -1,    -3,    -2,     0,     3,     3,     1,     0,    -4,    -2,    -4,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -3,    -1,    -2,     1,    -1,     1,    -2,    -1,     1,    -2,     0,     3,     0,    -1,    -2,     1,    -2,     0,     0,     0,    -2,    -1,    -2,    -1,    -3,    -4,     0,     1,     0,     1,     0,    -1,     1,    -1,     1,     1,     0,     2,     1,     0,     0,     0,    -4,    -2,    -4,     0,     0,    -2,    -3,    -1,    -1,    -4,    -3,    -2,    -1,    -2,    -1,    -1,     1,     0,     0,     1,     2,    -1,    -1,    -2,    -2,     0,     0,     0,    -2,    -1,     1,     0,     0,    -1,    -4,    -2,    -2,     2,     1,    -2,    -5,    -4,     1,     0,     2,     1,     1,     2,    -2,    -2,    -4,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     4,     1,    -2,    -2,    -1,     1,     2,     1,     0,    -1,     0,    -3,    -5,    -2,    -2,    -1,     0,    -2,    -3,     0,    -2,    -1,     0,     0,    -1,    -1,    -1,     1,     2,     0,     1,     3,     2,     2,     1,    -2,    -3,    -3,     0,    -4,    -6,    -3,    -2,    -1,    -2,    -3,    -2,     0,    -4,    -2,     0,    -1,     0,    -1,     0,     1,     3,     5,     4,     3,     2,     0,    -3,    -2,    -3,    -2,    -3,     0,    -3,    -2,    -2,    -4,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     2,     3,     3,     3,     2,    -2,    -3,    -4,     0,     2,    -2,    -3,     0,     0,    -1,    -2,    -3,    -3,    -1,    -1,    -1,     0,    -2,     0,     0,     0,    -2,     1,     4,     2,    -1,     0,    -2,    -4,    -3,    -1,     1,     0,    -1,    -2,     0,     1,    -3,    -2,    -3,    -3,    -2,     0,     0,    -2,    -1,     0,    -1,     0,    -3,    -1,     3,    -1,     1,     1,    -3,    -3,    -2,    -3,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -4,    -3,    -3,    -1,    -1,     0,    -2,     0,    -2,    -1,    -1,    -2,     0,     3,     0,     0,     2,    -2,    -1,     0,    -2,    -2,    -2,    -3,    -2,    -2,    -3,    -4,    -4,    -3,    -1,    -1,     0,     0,    -2,     0,    -2,    -1,     0,    -1,     1,     0,     0,     1,     2,    -1,     0,     0,    -3,    -2,    -1,    -3,    -1,    -2,    -3,    -2,    -4,    -3,    -1,    -1,    -1,     0,    -2,     0,     0,     0,     0,    -2,    -1,    -2,    -2,     1,     0,     1,     0,     0,    -1,     0,    -2,     0,     1,    -2,    -4,    -3,    -3,    -2,     0,    -1,    -1,    -1,    -3,     0,     0,     0,    -1,    -1,    -2,    -1,     2,     3,     3,     4,     1,     1,     1,    -1,    -2,     0,    -2,    -2,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -1,    -3,     0,     2,     1,     0,    -1,     0,     1,    -1,     2,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,    -2,    -1,    -2,    -3,    -2,     1,     0,     1,     0,     1,    -1,    -2,    -2,     0,    -1,     0,     0,    -2,    -1,    -2,     0,     0,     1,     1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0),
		    39 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,    -2,    -2,     0,    -1,    -1,    -1,    -2,    -1,     0,    -1,     0,     0,     0,     0,     1,     0,     1,     0,     1,    -1,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,     0,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -3,    -4,    -2,    -4,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -3,    -2,    -1,     0,    -1,    -1,     0,     0,     1,     0,     0,    -1,    -2,    -3,    -5,    -1,    -2,    -2,     0,    -1,    -2,    -3,    -4,    -5,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,    -1,    -4,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -3,     1,     2,     0,     0,     1,    -2,    -4,    -2,    -3,    -6,    -3,    -2,    -3,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -2,    -3,    -5,     1,    -2,     2,     2,     3,     1,     0,     4,     0,    -3,    -4,    -3,    -5,    -2,    -5,    -2,     1,     1,    -3,    -1,     0,    -1,     1,    -1,    -3,    -2,    -4,    -4,    -3,    -2,     0,     3,     1,     0,     0,     1,    -1,    -4,    -1,    -4,    -2,    -3,    -6,    -2,     1,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -3,    -2,    -3,    -2,    -3,    -2,     0,    -1,    -1,    -2,     0,     1,     2,    -1,    -3,    -2,    -3,    -2,    -3,    -3,     0,     0,    -1,    -2,    -1,     0,     0,    -1,    -3,    -1,     0,    -1,     1,     3,     1,    -2,    -3,     1,     0,     2,     1,    -1,    -2,    -1,    -2,    -4,    -2,    -4,    -2,    -2,    -3,    -3,    -1,    -1,     0,    -2,    -3,     0,     3,    -1,     2,     0,     1,    -2,     0,    -1,    -1,    -1,    -2,     1,     0,    -1,    -1,    -3,    -2,    -1,    -6,    -6,    -3,    -2,     0,    -2,     0,    -4,    -1,     2,    -1,     0,     4,     3,    -2,    -3,    -2,    -3,    -1,     1,     1,     2,     1,     2,    -2,     0,    -1,    -2,    -5,    -4,    -3,    -5,     0,    -2,     0,    -3,    -2,     1,    -1,     2,     3,    -1,    -2,    -1,    -2,    -4,    -1,    -1,     2,     1,    -1,     2,     0,    -1,     0,     1,    -2,    -2,     0,    -4,    -3,    -1,     0,    -3,    -1,     0,    -2,     3,     0,     0,     0,    -1,     1,    -3,    -2,    -1,     0,    -2,    -1,     0,     1,     0,     2,     1,     0,    -3,     0,    -3,    -2,    -1,    -1,    -1,    -1,     3,     0,     1,     0,     0,    -1,     2,     3,     3,     0,     1,    -1,    -4,    -2,     1,     2,     0,    -1,     1,     1,     0,     1,    -4,    -2,     0,     0,     0,    -1,     3,     1,     2,     2,    -2,     1,     1,     0,     1,     3,    -3,    -1,    -3,    -5,    -1,     1,     1,     1,    -1,    -1,     0,     1,    -4,    -2,    -2,     0,    -1,    -2,     1,     4,    -2,     2,    -1,     0,    -1,    -1,    -1,     0,    -1,    -4,    -4,    -3,     0,     3,     3,    -1,    -1,    -3,     0,     2,     0,    -2,    -3,     1,     0,    -2,     0,     1,    -1,     0,    -2,     0,    -1,     0,     0,     1,     1,    -1,    -2,    -1,     1,     0,     3,    -1,    -1,    -4,    -1,    -1,    -3,    -3,    -3,     0,     0,    -2,     1,    -2,     2,     1,     1,    -1,     0,     1,     2,     0,     0,     2,     2,     2,    -2,     0,     1,     1,    -4,    -3,    -2,    -1,    -3,    -3,    -2,     0,     0,    -2,     0,    -2,    -1,     1,     2,     0,     2,     1,     1,     4,     2,     0,     0,     0,    -4,    -3,     1,     1,    -1,    -1,     1,     0,    -4,    -2,    -1,    -1,    -1,    -1,     0,     1,     0,    -3,    -3,     1,    -2,     0,    -2,    -3,    -2,    -2,    -4,    -3,    -4,    -1,     3,     1,    -1,    -1,     1,     5,     0,    -4,     0,     0,     0,    -2,    -1,     0,     0,    -1,    -3,    -6,    -6,    -2,    -2,    -3,    -3,    -4,    -4,    -6,    -3,    -2,     2,     0,     0,    -1,     0,     3,    -2,    -5,     0,    -1,     0,    -2,     1,    -1,    -1,    -1,    -2,    -4,    -5,    -1,     2,    -1,     2,    -1,    -3,    -1,    -3,     0,     1,     1,     0,     1,     0,     2,    -4,    -2,    -1,     0,    -1,     0,     2,     1,     0,    -1,    -2,    -2,    -2,    -2,    -2,     0,     1,     0,    -1,    -2,    -2,    -1,    -1,     1,     0,    -1,     3,     4,    -3,    -2,     0,     0,     0,    -2,     0,    -1,     0,    -1,    -1,    -2,    -3,    -2,    -3,     0,     0,     0,    -2,    -1,     0,     1,     3,     5,     1,     4,     6,     1,     1,     0,    -1,     0,     0,     2,    -1,    -1,     1,    -1,    -2,    -2,    -2,    -1,     1,     0,     1,    -3,    -4,    -4,    -3,    -1,     3,     2,     1,     0,    -2,    -2,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     1,     1,     1,     0,     0,    -1,    -1,     1,     1,    -1,    -3,    -3,    -3,    -3,     0,     0,     1,     3,     2,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     0,     0,     0,     1,     1,     1,     0,    -2,    -2,     1,     1,    -2,    -3,     0,    -2,     0,     0,     0,     0),
		    40 => (   -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     1,     0,     0,     1,     2,     2,     0,     0,     1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     1,     2,     1,     0,     0,     0,    -2,    -4,    -3,    -2,    -3,    -5,    -4,    -5,    -1,    -2,    -2,    -3,    -3,    -1,    -3,    -2,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,    -2,    -1,    -1,     0,     0,    -2,    -1,     0,     0,    -1,    -1,    -2,    -4,    -5,    -1,    -1,    -3,    -2,    -2,    -1,    -2,     0,     1,     0,     0,    -1,     0,    -4,    -3,    -2,    -1,     2,     0,    -1,    -3,     0,     0,    -1,     1,    -2,    -3,    -2,    -2,    -1,     1,    -3,    -2,    -2,    -3,     0,     0,     0,    -1,     1,     0,    -2,     0,     0,     2,    -1,     0,    -2,    -2,     1,     0,    -2,    -1,     1,     0,    -2,    -3,    -2,    -1,    -2,    -1,    -2,    -2,    -2,     0,     0,    -1,    -1,     2,     2,     1,     0,    -4,    -3,     0,    -1,    -2,     1,    -1,    -2,     1,     1,    -2,     2,     0,     2,     1,    -4,    -2,    -4,    -2,    -1,     0,     0,    -1,    -1,     2,     2,     0,    -1,    -4,     1,    -1,    -2,     0,    -1,     0,     0,     1,     2,     4,     3,     1,     1,     1,     1,    -3,    -2,    -5,     2,     4,    -2,     2,     0,     2,     1,    -1,     0,     0,     0,    -1,    -1,     3,     0,     2,     1,     2,     2,     3,    -2,     0,     1,     1,     2,    -4,    -5,    -4,    -1,     0,    -1,     3,     0,    -4,     0,    -1,    -1,     1,     0,    -2,    -2,     0,    -1,     1,     0,    -2,     1,     2,    -1,     4,    -1,     0,    -1,     0,    -5,    -5,     0,     0,     0,     3,     0,    -2,    -3,     0,    -1,     0,    -1,    -2,    -3,     0,     0,     2,     0,    -1,     1,     0,    -1,     3,     2,     3,    -1,     0,    -4,    -4,     0,    -1,     6,    -2,    -1,    -3,    -3,     2,     3,     1,     1,    -1,    -1,     1,    -1,     1,    -2,    -2,     1,    -2,    -1,     2,     3,     2,    -2,    -2,    -4,    -4,     0,     0,     1,    -1,    -1,    -3,    -2,     4,     2,     1,     1,     0,     1,     0,    -2,    -3,    -2,    -4,    -3,    -1,    -1,     1,     3,     1,     0,     0,    -1,    -4,     0,     0,     1,     1,     2,    -1,     1,     2,     3,     4,     2,    -1,     1,    -3,    -3,    -1,    -5,    -4,    -4,     1,     0,     1,     2,     3,     2,     1,     2,    -2,    -1,     0,     1,     0,     1,     1,     4,     3,     5,     3,     1,     0,     1,    -1,     0,    -3,    -3,    -5,    -2,    -1,     2,     1,     0,     0,     3,    -1,     0,    -3,     0,     0,     0,    -1,    -1,     0,     2,     0,     2,     5,     2,     0,     0,    -1,    -2,    -3,    -3,    -2,    -4,    -1,     0,     2,     3,     2,     4,     3,     1,    -5,    -1,     0,     0,    -1,    -2,     2,     0,     3,     4,     1,     1,     1,    -2,    -3,    -3,    -4,    -3,     0,    -1,     1,    -2,    -1,     3,     2,     0,     2,    -2,    -5,     3,     0,     0,    -2,    -4,     1,    -2,     0,     0,     2,     3,     0,    -3,    -5,    -3,    -1,     2,     0,    -1,    -2,    -2,     1,    -2,     3,    -1,     1,    -3,    -4,     4,     1,     0,    -1,    -4,    -1,    -3,    -1,     2,     5,     3,     1,    -2,    -5,    -2,     2,     1,     0,    -1,     0,     0,     1,     0,     2,    -2,     0,     0,    -2,    -2,     0,     2,    -2,    -2,    -1,    -2,    -2,    -1,     4,     2,     1,    -4,    -2,    -2,    -2,    -1,     0,    -2,    -1,    -2,     3,    -1,     1,     0,     0,    -5,     0,     0,     0,     1,    -3,     0,    -1,     1,    -1,    -1,     2,     3,     5,    -2,     0,    -1,    -1,    -2,    -2,    -1,    -2,    -1,    -3,    -2,    -1,    -4,    -3,    -2,     1,     0,     0,    -1,    -4,    -2,    -1,     0,    -2,    -2,     1,    -1,     0,    -2,    -2,    -3,    -2,     0,     1,    -1,    -4,    -3,    -2,    -1,     2,    -1,    -2,    -2,     2,     1,     0,    -1,    -4,    -1,    -4,    -1,     0,     0,     3,     2,     2,    -2,    -1,    -1,    -1,     0,    -3,    -3,    -2,     0,    -2,     0,     1,    -1,    -1,     0,     2,     1,     0,     1,     0,    -4,    -3,    -2,     0,     0,     0,     1,     1,     2,    -1,     0,    -1,    -1,    -2,    -2,    -4,    -2,    -4,    -1,    -3,    -2,    -3,    -1,    -2,     0,    -1,    -1,    -1,     0,     0,     2,    -2,    -3,     0,     2,     2,     2,     2,    -2,    -1,     1,    -2,    -4,    -3,    -3,    -2,    -3,    -3,    -3,    -1,     1,     0,     0,     0,     1,    -1,     0,    -3,    -5,    -4,    -3,    -3,    -3,    -5,    -5,    -5,    -3,    -2,    -6,    -6,    -6,    -7,    -5,    -4,    -3,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -5,    -2,    -2,    -4,    -4,    -5,    -3,    -3,    -3,    -4,    -3,    -5,    -5,    -3,    -4,    -3,    -1,    -2,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,     0,     0,     0,     0),
		    41 => (    1,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,     0,     1,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -1,     3,     4,     5,     5,     3,     3,     5,     4,    -3,    -4,    -3,     0,     0,     0,     0,     1,     0,     2,     4,     0,    -2,    -3,     2,     2,    -1,    -5,    -5,     0,     0,     1,     2,     5,     2,     2,     2,     4,     4,    -2,    -2,    -1,    -1,     1,     1,     1,     0,     0,     2,     0,     1,    -1,    -3,    -2,    -1,     1,    -1,    -3,    -4,     1,     3,     3,     1,     3,     1,     1,     2,    -2,    -2,    -1,    -3,    -3,    -2,    -1,     0,     2,     1,     0,     3,     1,    -3,    -2,    -2,    -1,    -1,    -4,    -2,    -1,     2,     3,     1,     0,    -1,    -1,     2,    -2,    -1,    -1,    -2,    -2,    -1,     0,     0,    -2,     0,     0,     1,    -2,    -3,    -2,    -2,    -3,    -3,    -1,     1,     1,     2,     3,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,     0,    -1,    -3,    -1,    -2,    -4,    -5,    -1,     2,     1,    -1,     0,     0,    -1,     3,     1,     0,     1,    -5,    -3,    -1,    -2,    -3,    -1,     0,     0,    -2,    -2,    -1,    -1,    -3,     0,    -2,    -5,    -2,    -2,     1,     6,     0,    -2,    -1,    -1,     1,     2,     0,    -1,    -1,    -3,     0,    -2,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,    -4,    -1,    -2,    -2,     0,     1,     3,     2,     1,    -2,    -2,    -1,     1,     2,     2,    -4,    -2,    -5,    -2,    -3,    -1,    -2,    -1,    -1,    -1,    -2,     1,     0,    -4,     0,    -3,    -4,    -2,     2,    -2,    -2,    -1,     0,     0,    -2,     0,     0,     0,     0,    -2,    -2,    -2,    -3,    -1,    -1,    -1,    -1,    -2,     2,     0,     1,     0,     0,    -2,    -2,     0,    -1,    -4,     1,     2,     0,     0,    -3,     0,     0,    -1,    -2,    -5,    -2,    -3,    -1,    -2,     0,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -3,     2,     0,     2,    -2,    -5,     0,     0,     1,    -4,    -2,    -4,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -2,    -1,     3,     1,     0,    -1,    -8,     0,     1,     0,    -2,    -6,    -4,    -2,    -3,    -2,    -4,    -3,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -3,    -4,     3,     2,     1,    -3,    -8,    -4,     2,     0,    -1,    -4,    -6,    -4,    -4,    -3,    -3,    -3,    -1,    -1,     1,     0,     0,     0,     1,     1,    -3,    -3,    -4,    -3,     3,     2,    -2,    -5,    -6,     1,     1,     0,     0,    -5,    -6,    -5,    -4,    -2,    -2,    -3,    -2,    -1,     0,    -2,     0,     0,     0,    -1,    -2,    -3,    -2,    -2,    -1,    -1,    -7,    -6,    -8,    -1,    -2,    -2,    -4,    -6,    -7,    -5,    -3,    -2,    -2,    -4,     1,    -2,    -3,    -1,     0,     0,     0,    -2,     0,     1,     4,    -1,    -2,    -2,    -1,    -5,    -6,    -2,     0,    -3,    -2,    -3,     0,     3,     1,     0,    -1,    -4,     0,    -5,    -1,    -2,     0,     0,     0,    -1,    -1,     3,     0,    -1,     1,    -1,     0,    -5,    -6,    -1,     0,    -1,     1,     0,     1,     2,     3,     0,    -1,    -1,     0,    -2,    -3,     0,     0,     0,     1,    -1,    -2,    -1,     0,     0,     1,     1,    -1,    -1,    -3,    -1,     0,     1,     3,     0,    -1,     2,     3,    -1,     0,     1,     0,    -2,    -3,    -2,     0,     0,     1,     3,     3,    -6,    -1,    -2,    -1,     5,     1,     0,     0,     2,     2,     1,     3,     1,     3,     3,     2,     1,     4,     2,     0,    -1,    -1,     1,     2,     2,    -1,     4,     4,     2,    -1,     2,     2,     2,     3,    -2,    -1,     2,    -1,     0,     1,    -1,     1,     0,     2,     3,     0,    -1,     1,     1,    -2,     0,     1,     1,    -2,     2,     1,     5,     4,     0,     1,     1,     0,     0,     0,     0,    -3,     0,     0,     0,     0,     0,     1,     2,     2,     3,     3,     3,     1,     0,     1,     0,     0,    -1,     0,     2,     4,    -2,    -3,     1,     0,    -2,     0,     0,     0,     1,     0,    -1,    -3,    -9,    -7,    -5,    -1,    -3,    -3,    -2,     1,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -2,    -1,     1,     1,    -1,     1,     0,     1,     0,    -3,    -4,    -3,    -4,    -3,     0,    -2,    -2,    -4,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     1,     0,     0,    -1,    -4,     0,     1,    -2,    -8,     0,    -1,    -2,    -3,    -2,    -2,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,    -1,     0,    -2,    -2,     0,     0,    -4,    -4,     1,     2,     2,    -2,    -1,     0,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -2,     0,     0,     0,     0,     1,     0,     1,    -1,     0,     0,     1),
		    42 => (   -1,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,    -1,     1,     1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,    -1,    -2,     1,     0,    -1,    -4,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,    -2,    -1,     0,     0,    -1,     0,     0,     3,     3,     0,     1,     2,     2,     3,     3,     1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -3,    -1,    -1,    -2,     1,     2,     4,     0,    -1,     0,    -1,    -1,     1,     3,    -2,     0,     0,     2,     0,    -2,    -1,    -1,     0,     0,     0,    -1,    -1,    -2,     0,    -1,    -1,     0,     3,     5,     2,     0,     3,    -1,    -1,     0,     2,     1,     1,    -1,    -3,    -2,    -1,    -2,    -3,    -2,    -4,    -2,     0,     0,    -1,     0,    -1,     0,     1,     1,     0,     1,     2,     4,     1,     3,     3,     2,     3,    -1,    -1,     2,     1,     0,    -3,    -2,    -2,    -1,    -5,    -2,     0,     0,     1,    -2,    -1,     2,     2,     3,     2,     1,     2,     1,     0,    -1,     1,     2,     2,     1,     3,     0,     1,     3,    -2,    -6,    -6,     0,    -4,    -1,     0,     0,     2,    -1,    -1,     1,     2,     3,     1,     0,    -1,    -1,     2,     2,     0,     2,     2,     1,     0,    -1,    -1,     1,    -3,    -3,     0,     3,    -7,    -3,    -2,     2,     2,    -1,     0,     1,     1,     0,    -1,     0,    -2,     1,    -1,    -1,    -1,    -2,     1,    -1,    -2,    -1,    -3,    -2,    -1,     4,     2,    -1,    -5,    -3,     0,    -3,     3,     1,     0,     0,     1,     0,     0,     1,     2,     0,    -2,    -2,    -3,    -1,    -1,    -1,    -3,    -3,    -1,     1,    -1,     2,     0,    -4,    -2,    -1,    -1,    -1,     3,     0,     1,     0,     0,     0,    -2,     0,     1,     1,     3,     0,    -1,     0,     0,     1,    -2,    -2,    -2,    -1,    -3,    -3,    -1,    -2,    -1,    -2,     0,    -2,    -1,    -2,     0,     1,     0,    -1,    -1,    -3,     0,     1,     2,    -2,     0,     1,     0,    -1,    -3,    -1,     1,     0,    -2,     1,    -1,     2,    -3,    -3,     0,    -1,    -4,    -1,     0,     0,     0,    -1,     2,     4,     2,     1,     2,    -2,     1,     0,    -1,    -1,     0,     3,    -1,     2,     3,     2,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     2,     2,     3,     1,     0,    -1,     0,     0,     0,    -1,     0,     1,     3,     3,     2,     2,     2,     1,    -1,    -2,     3,     0,     0,    -2,    -1,     0,    -3,    -3,     1,     4,     3,     1,    -2,    -1,    -2,    -2,    -3,    -1,    -1,     0,     4,     3,     2,     3,     4,     5,     4,     1,     2,     2,     1,    -1,     2,     1,    -2,    -1,     0,     1,     3,     1,    -2,     1,    -1,    -5,    -4,    -1,    -1,     1,     0,     3,     4,     3,     2,     3,     0,     1,     0,     2,     0,     0,     3,    -2,    -2,    -3,    -1,     2,     2,     2,     1,     1,    -2,    -3,    -3,     2,     0,     1,     4,     4,     4,     5,     3,     6,     2,     2,     3,     2,     0,     0,     3,    -1,    -3,    -1,    -2,    -1,     2,     4,     3,     2,     1,    -1,     0,     1,    -2,     0,     3,     5,     3,     1,     1,     1,    -1,    -2,     3,     2,     0,     0,     0,    -1,    -1,    -1,     0,     0,     1,     3,     5,     2,     0,    -1,    -2,    -1,     0,     3,     5,     6,     5,     2,     1,     1,     1,    -3,    -1,     3,     0,    -1,    -2,     0,    -1,     0,    -1,     1,     1,     3,     3,     1,     1,    -3,     0,     0,     0,     8,     8,     7,     3,     2,     2,     1,     1,    -3,     0,     2,     0,    -1,     1,     1,     0,    -2,    -3,     0,     2,     1,     2,     2,     2,    -1,    -2,     1,     6,     5,     6,     4,     2,     0,    -2,     0,    -1,    -1,    -1,     0,     0,     0,     2,     0,     3,    -1,    -3,     0,     0,    -1,    -1,     0,     0,     1,    -1,     4,     7,     6,     4,     5,     1,    -1,    -1,    -1,    -3,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -2,    -2,     0,    -2,    -1,     0,     3,     0,    -1,     4,     9,     6,     7,     3,     2,    -1,    -1,    -1,     0,     2,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     2,    -2,    -5,    -3,     0,     1,     3,     7,     9,     8,     6,     3,     0,     2,    -2,     0,     1,     1,    -2,     0,     0,     0,    -2,    -2,    -7,    -7,    -2,    -1,     0,    -4,    -4,    -2,    -2,     3,     4,     3,     7,     6,     5,     1,     0,     0,    -2,    -1,     1,     0,     1,     0,     0,     1,     0,    -1,    -3,    -4,     3,     1,    -1,    -2,     0,     3,     5,     6,     7,     6,     4,     2,     2,     1,    -1,    -1,    -4,     0,     1,     2,     1,     0,     0,     1,     0,     0,    -1,    -3,    -5,    -4,    -4,    -5,    -5,    -3,    -4,    -3,    -5,    -3,    -3,    -3,    -3,    -4,    -2,    -2,    -5,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,    -3,    -4,    -1,    -1,    -1,     0,    -1,     0),
		    43 => (    0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -2,    -4,    -5,    -6,    -2,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -4,    -4,    -1,     0,     0,     0,     0,     0,     1,     0,    -2,    -2,    -2,    -3,    -3,    -4,    -1,     0,     0,     0,     0,     0,     0,    -2,    -1,     1,     0,     1,     2,    -1,     0,     1,     4,     0,     0,     4,     4,     3,     1,    -2,     0,    -2,    -3,    -7,    -5,    -2,     0,     0,     0,     3,    -4,     1,     1,    -1,    -3,    -3,     1,     2,     3,    -1,     0,     0,     0,     1,     2,    -1,    -2,    -3,    -2,    -1,     3,    -3,    -7,    -6,    -2,     0,     0,     0,    -1,     1,    -1,     0,     1,     1,     0,     0,     0,     0,     0,     1,     0,     1,     2,    -1,    -4,     0,     2,    -1,    -2,     3,    -1,    -7,    -2,     0,     0,     1,    -3,    -1,    -3,     0,     3,     2,     0,     1,    -1,    -3,    -3,     0,     1,     2,     2,     3,     2,     2,     1,     3,     1,     1,     4,    -6,    -5,    -2,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     0,    -2,    -1,     0,     1,     1,     0,    -1,     2,     2,     1,    -1,     1,    -1,     5,     2,    -8,    -5,    -3,    -2,    -1,     1,     2,     1,     0,    -1,     1,    -1,    -1,     1,     0,     2,     2,    -2,    -3,    -1,     1,     1,     3,     0,    -2,     2,     2,     0,    -9,    -6,     0,     0,    -3,     0,    -1,     2,     0,    -2,    -3,    -3,     0,    -3,    -1,     6,     4,     2,     1,     2,     1,     0,     1,     2,     0,     4,     3,    -5,    -7,    -6,    -3,     0,    -3,     1,     1,    -2,    -2,    -4,    -4,    -5,    -5,    -6,    -1,     3,     5,     7,     2,    -2,    -1,    -2,    -1,     0,     1,     0,     1,    -5,    -3,    -5,    -3,     0,    -2,    -1,     3,     0,    -2,    -6,    -5,    -2,    -4,    -7,    -2,     1,     5,     3,     3,     1,     0,     0,    -2,    -1,    -2,    -2,    -5,   -12,    -6,    -4,    -1,     0,    -1,     0,     0,    -1,     0,    -2,    -4,    -1,    -7,    -1,    -3,     1,     3,     7,     4,    -1,     1,     2,    -2,     0,    -1,    -7,    -8,    -9,    -4,    -3,    -1,     0,    -1,    -7,    -2,    -2,    -2,    -1,    -2,    -1,    -3,    -3,    -2,     1,     2,     5,     2,     5,     1,     1,     1,     1,    -2,    -5,    -2,    -5,    -5,    -3,    -1,    -1,     2,     0,    -4,    -5,    -3,    -2,    -2,    -2,    -1,    -4,    -1,     0,     3,     2,     3,     1,     0,    -3,    -2,    -2,    -3,    -2,     0,    -4,    -5,    -3,    -1,     0,     1,     0,    -3,    -1,    -1,     1,     0,     1,    -4,    -4,     1,     4,     4,     3,     4,    -1,    -4,    -5,    -2,    -1,    -1,     2,     2,     2,    -4,     1,    -2,     0,     0,     1,     2,     0,    -1,     0,     0,     0,    -2,    -1,     2,     1,     1,     3,    -1,    -5,    -3,    -1,    -1,    -2,    -2,     3,     1,     2,    -7,    -4,    -2,     0,     1,     2,     2,     1,    -2,    -1,    -1,    -3,    -2,     0,     3,     0,     2,     0,    -3,    -4,    -2,    -2,    -1,    -3,    -1,     0,     0,     0,    -5,    -1,    -2,    -1,     1,     2,     3,     0,    -1,     1,     2,    -2,    -1,     2,     4,     0,     0,    -2,    -2,    -1,     0,    -2,     0,     1,     2,    -1,    -2,    -3,    -5,    -1,    -3,     0,    -2,     2,     5,     2,     3,    -2,     2,     0,     1,     3,     1,    -3,    -2,    -4,     1,     1,     2,     2,     0,     1,     1,    -2,    -1,    -2,    -4,    -4,    -3,     0,    -2,    -3,     1,     0,    -2,    -2,     1,     2,     1,     2,     1,    -3,    -1,    -1,     2,     2,     1,     0,    -1,    -1,     1,    -1,     0,    -2,    -3,    -1,     0,     0,    -1,    -2,     1,     0,    -4,     0,     2,     2,    -1,    -2,    -2,    -2,     0,    -1,     0,    -1,     0,     0,     0,    -2,    -1,     0,    -2,    -6,    -4,    -1,     0,     0,     0,    -1,     1,    -2,    -2,     3,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -1,    -1,     0,     0,    -4,    -5,    -7,    -1,     0,     0,     0,     1,     4,    -1,     0,     3,     1,     2,     1,     3,     2,    -2,     2,    -2,     0,     2,     0,     2,    -1,    -2,    -2,    -3,    -3,     3,     1,    -2,     0,     0,     0,     1,     4,    -1,     0,     1,     0,    -2,    -2,     0,     5,    -3,     0,     4,    -1,    -1,    -2,     0,     0,     0,    -1,    -2,    -2,    -3,    -3,    -1,     1,     0,     0,     0,    -2,    -2,    -2,    -3,     1,     1,     0,     4,     4,     7,     2,     0,    -2,     2,     0,     1,     2,    -3,    -5,    -6,    -7,    -3,    -1,    -1,     0,     0,     1,     0,    -2,    -4,    -2,    -2,    -1,     0,    -1,     2,     1,     2,     1,    -4,    -2,     0,     1,     1,    -2,    -2,    -4,    -5,    -3,     0,     0,    -1,     0,    -1,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,    -3,    -4,    -4,    -3,    -6,    -3,    -3,    -2,    -1,    -1,    -4,    -4,    -2,     0,     1,     0,     0,     0,     0),
		    44 => (    0,     0,     1,     1,    -1,     0,     1,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     1,     0,     1,     0,     0,     1,    -1,     0,    -1,    -1,    -1,     0,    -1,    -3,    -1,    -4,    -3,     0,    -2,    -2,     0,    -1,     0,    -2,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -4,    -2,    -3,    -2,    -2,    -1,    -4,     1,     0,    -2,    -5,    -3,    -2,    -2,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -4,    -6,    -3,    -4,    -3,    -4,    -2,     2,    -2,    -4,    -8,    -5,     0,    -1,     0,    -3,    -3,    -1,    -1,    -3,    -1,     0,    -1,     0,     1,    -1,     0,    -1,    -3,    -1,     1,     1,     0,    -1,     0,    -3,    -6,    -1,     1,    -5,    -7,    -7,    -6,    -3,    -1,     0,     0,     1,     2,     3,     1,    -2,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -3,    -6,    -4,     0,     4,    -1,    -2,    -1,    -3,   -12,    -6,     1,     3,     1,     0,     0,     0,     0,    -2,    -1,    -1,     0,     0,    -2,     2,     6,    -1,    -4,    -2,    -2,    -3,     1,     3,     1,    -2,    -2,    -9,    -9,    -4,     3,     2,     1,     0,     2,     3,    -6,     2,    -5,     0,    -4,     0,    -2,     1,     5,    -3,    -1,    -1,     0,     1,     2,     0,     2,    -1,    -5,   -10,   -10,    -1,     3,     1,    -1,     0,     1,    -1,    -1,     2,    -5,    -2,    -4,     1,    -1,     0,     1,    -2,     1,    -2,     0,    -2,     0,     2,     1,     1,    -5,   -12,    -4,     2,     2,     1,    -1,     2,    -2,     0,     3,     1,    -3,     0,    -3,     0,    -2,    -1,     1,    -2,    -1,    -1,     1,     0,     0,     3,     3,     2,    -6,    -6,     2,     3,     1,     2,     1,     1,     1,     3,    -3,    -3,    -2,     0,    -2,    -3,     1,     2,     3,     0,    -2,     0,     1,    -1,    -1,     0,     4,    -2,    -7,    -5,     1,     3,     3,     0,     0,     1,     2,     1,    -6,    -2,     0,    -1,    -1,    -2,    -4,    -2,     1,     3,    -1,     1,    -1,     1,     0,     3,    -1,    -5,    -7,    -4,    -2,     1,     1,    -3,     2,     0,    -1,     2,    -3,    -3,    -2,     0,     0,    -3,    -4,    -5,    -2,     1,     3,     2,    -2,    -1,     2,     3,     2,    -6,    -3,    -1,    -1,    -1,     2,     0,     3,     1,     2,    -3,    -3,    -6,    -3,     0,    -1,    -3,    -4,    -4,    -2,    -1,    -1,     1,     1,     2,     3,     1,     1,     0,     1,     1,     2,    -2,     2,     2,     1,     0,    -1,    -6,    -5,    -5,     0,     0,    -1,    -1,    -4,    -3,     0,     0,     0,    -1,     2,     0,     2,     0,    -1,     2,     1,     0,     0,    -1,     2,     1,    -1,    -2,    -1,    -3,    -3,    -4,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     2,     1,     2,     1,     0,     1,     1,     0,    -1,    -1,     0,     3,    -6,    -2,    -1,    -1,    -3,    -4,    -3,     0,     0,    -1,    -2,     1,     0,    -1,    -4,     0,     0,     0,     0,     0,    -1,     0,    -2,     0,    -1,    -1,    -1,    -1,    -4,    -2,    -1,    -2,    -4,    -5,    -5,    -1,     0,     0,    -2,     1,     3,     0,    -3,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,    -2,     1,    -1,    -3,    -5,     1,    -1,    -1,    -4,     0,    -1,    -1,    -2,     0,    -3,     4,     6,    -2,    -2,    -3,    -2,    -3,    -6,     0,    -2,     0,     1,     0,     1,    -3,     0,    -1,     0,     2,     1,     1,     0,     2,     0,    -1,     0,    -3,    -1,     3,     2,    -3,    -3,    -2,    -1,    -3,    -3,    -1,    -3,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,     1,     1,     1,     2,     1,    -1,    -1,     1,     0,    -1,    -4,    -4,    -5,    -4,    -2,    -3,     0,    -2,    -2,    -2,     0,    -1,    -1,     1,     0,    -2,    -2,    -4,    -4,    -2,    -1,    -4,    -6,    -1,     0,     0,     0,    -1,    -3,    -4,     5,     0,     1,     3,     4,    -1,     0,     0,     0,    -1,    -1,    -1,    -4,    -4,     0,     0,    -1,     1,     2,    -2,    -8,    -3,    -1,    -1,     1,     0,    -3,    -5,     3,     3,     2,     2,     0,     2,     0,     0,     0,    -2,    -1,     0,    -2,    -3,    -1,     0,     1,     0,     2,    -2,    -2,     1,     1,     0,     0,     0,    -3,    -4,    -8,     1,     2,     2,     1,     1,     0,     1,    -1,     1,     1,     2,    -2,    -2,    -1,    -1,     1,     1,     1,    -2,     0,     1,     0,     0,     0,     0,    -1,    -6,    -5,    -1,    -3,     0,     1,     1,    -1,     1,     0,     0,     2,     1,    -3,    -7,    -2,    -1,     2,     1,     2,    -2,     3,    -2,    -1,     1,    -1,    -1,     0,     0,    -4,    -3,     0,     0,    -2,     0,     1,     1,     2,     0,    -2,    -3,    -6,    -3,    -2,    -1,    -1,     2,     4,    -1,    -2,     0,     0,     0,     0,     0,    -3,     0,    -3,    -3,    -5,    -3,    -3,    -4,    -2,    -5,    -6,    -7,   -10,    -2,    -3,    -4,    -2,    -3,    -3,    -2,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -2,    -3,    -4,    -1,    -2,    -4,     0,    -3,    -4,    -2,    -2,     0,    -1,     0,     0,     0,     1,     0,     0),
		    45 => (    0,    -1,     0,     0,     0,    -1,     0,    -1,     1,    -1,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -3,    -2,    -3,    -3,    -3,    -2,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -3,    -1,    -2,    -1,    -2,    -3,    -3,    -3,    -1,    -2,    -2,    -2,    -2,    -3,    -2,     2,    -4,    -1,     0,    -1,     1,     0,    -1,     3,     6,    -1,    -2,    -3,    -1,     1,    -1,    -4,    -3,    -5,    -4,    -2,     1,     0,     0,     0,     0,     1,    -4,    -3,     0,     5,     4,     0,     0,     0,    -2,     5,     0,     0,    -3,    -2,    -2,    -1,     0,    -5,    -5,    -3,    -3,    -2,    -3,    -3,     0,     3,     0,     0,    -3,     0,     4,     3,     0,    -1,     0,     0,    -3,     5,    -1,    -1,    -2,    -3,    -3,    -1,     0,     0,    -4,    -2,    -1,    -1,    -2,    -1,    -1,     2,     0,    -1,    -2,    -1,    -2,     1,     0,    -1,     0,     0,    -3,    -1,    -2,    -1,    -2,    -3,    -2,     0,    -1,    -3,     0,     0,    -1,     0,     0,    -2,     0,    -1,    -1,    -2,     4,     3,     2,     4,     4,     0,     0,    -1,     0,    -1,    -1,    -2,    -2,    -2,     0,    -1,     0,     0,     1,     2,     2,     1,     2,     3,    -1,    -2,     0,     2,     1,     2,     1,     0,     5,     1,    -2,     0,    -3,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,     2,     0,    -1,     1,     1,     5,     5,     2,     4,     3,     1,    -1,     2,     2,     1,    -1,    -5,    -4,    -2,    -2,    -3,    -1,    -1,    -2,    -2,     0,     1,     0,     1,     0,     0,     1,    -1,    -3,     2,     1,     2,     3,     7,     5,     1,     1,     0,     0,    -2,    -3,    -3,     1,    -1,     0,     1,    -2,    -2,     0,     2,     0,     0,     1,     2,    -3,   -10,   -11,    -6,    -5,    -5,    -2,     0,     1,     1,     2,     0,     0,     0,     2,     1,     1,    -1,    -1,    -2,    -4,    -1,    -3,    -3,    -2,     0,    -1,     1,    -1,    -5,    -6,    -9,    -9,    -9,    -7,    -6,    -1,     0,    -1,     0,     0,     0,     3,     1,    -1,    -3,    -4,    -4,    -3,    -1,    -3,    -4,     0,     2,    -1,    -1,     1,     0,    -1,    -4,    -7,    -6,   -11,    -7,    -4,    -1,    -2,     0,    -1,     0,     4,     0,    -2,    -1,    -2,    -2,     0,    -1,     0,     2,     1,     1,     1,    -1,     1,     2,     3,     2,     2,     0,    -4,    -6,    -2,     0,    -2,     1,     0,    -1,     2,    -3,    -4,     0,    -2,    -3,    -1,     0,     1,    -1,     0,     1,     2,     2,    -2,     0,     1,     3,    -1,     0,     3,     1,    -2,    -1,    -2,     1,     0,    -2,     0,    -2,     0,     1,    -1,    -1,    -3,    -1,    -1,    -1,     2,     0,    -2,    -1,     0,    -1,    -1,     3,     0,    -1,     2,     4,     0,     0,     0,    -1,    -2,    -5,     0,     1,    -3,     3,     1,     0,    -5,    -4,    -4,    -3,    -1,     0,    -2,     2,     1,     0,     0,     4,     3,     0,    -2,     0,     2,    -1,    -1,    -1,    -2,    -6,    -2,     2,    -1,     3,     5,     2,     0,     0,    -3,    -6,    -2,    -3,    -2,     0,     0,     0,    -2,     2,     0,    -4,    -3,    -1,    -1,    -2,    -1,     0,     0,    -4,     0,     1,     1,     2,     4,     2,     0,     1,    -1,     0,    -2,     0,     0,     0,     0,    -2,    -2,    -2,    -1,    -2,    -5,    -3,    -1,    -4,    -3,     0,    -1,     4,    -4,    -1,    -1,     2,     3,     2,     3,     2,     3,     3,     2,     1,     0,    -1,    -2,     1,     1,    -1,    -2,    -2,    -3,    -2,    -1,    -2,    -2,     0,    -1,     3,    -5,    -4,     0,     0,    -2,     1,     1,     2,     1,     1,     0,     1,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,     0,    -2,     1,    -1,     0,    -3,    -2,    -2,     1,    -1,    -1,     1,     0,     1,     1,     1,    -1,    -2,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -5,     2,     2,     0,    -3,     0,    -3,    -2,    -1,    -1,     0,    -1,     1,     1,     0,     0,     0,    -2,     0,     1,     1,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     3,     4,     0,    -2,    -3,    -2,     0,     0,    -2,    -3,     0,    -1,     0,     2,     2,     0,     0,     1,     1,     0,    -2,    -1,    -1,    -1,     0,     0,    -2,     0,    -1,    -1,    -3,    -5,    -5,    -2,    -5,    -6,    -2,    -1,    -2,    -3,    -3,    -2,     0,     2,     2,     0,     1,     0,     1,    -3,    -1,     0,     0,     1,     0,     1,    -2,    -1,     0,    -1,    -3,    -1,    -6,    -5,     0,    -1,    -2,    -1,     0,    -1,     0,    -1,    -1,    -2,     1,     0,     1,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,    -2,    -1,    -2,    -1,    -1,    -1,    -1,     2,     5,     4,     4,     2,     0,     3,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -3,    -1,     0,     0,     0,     0),
		    46 => (    0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     2,     3,     4,     2,     1,     0,     1,     1,     0,     0,     0,     1,     1,     4,     1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     3,     4,     4,     2,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,     2,     2,     1,     1,     2,     2,     1,     0,     0,     0,     0,    -3,    -2,     0,     0,     2,     3,     1,     2,     0,    -3,    -3,    -1,     0,     0,     0,    -1,    -1,     1,     0,     2,     0,     2,     3,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     1,     0,     1,     1,    -2,    -2,     0,    -2,    -1,     2,     1,     0,    -1,     0,     0,     1,     0,     1,     1,     0,     1,     2,     0,     0,     0,    -1,     1,    -1,     0,     1,     1,    -1,    -3,     0,     0,    -1,     1,    -1,    -2,     1,     1,     0,     1,     0,     0,     1,     1,     0,     3,     2,     0,     0,     0,     0,    -1,     0,    -1,     1,     0,    -1,     1,     0,     0,    -2,    -2,    -3,    -3,     0,     1,     1,     2,     2,     2,     1,     0,    -2,     1,     1,     0,     0,     0,    -1,     0,    -1,    -2,    -2,     1,     0,     0,    -1,    -3,    -1,     1,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,     1,    -1,     0,     1,     0,     0,     0,    -2,    -1,     0,    -1,    -2,     1,     1,     0,    -3,    -2,    -1,    -1,    -2,     1,     1,    -1,    -1,    -3,    -1,    -4,    -3,    -2,    -2,    -1,    -3,     0,     0,     0,    -1,    -1,    -2,     0,     0,     2,     0,    -1,    -2,    -2,    -2,    -1,     1,     0,    -1,    -2,    -3,    -4,    -3,    -5,    -3,    -1,    -2,     0,    -1,     0,     0,     0,    -1,    -1,    -2,     0,    -1,     1,    -2,    -2,    -3,    -1,    -2,     0,     1,     0,    -3,    -3,    -2,    -3,    -2,    -3,    -3,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     1,     2,     0,     0,    -2,    -3,    -2,    -1,     0,     1,     0,    -3,    -3,    -3,     0,     0,     0,    -1,    -1,     0,    -2,    -1,     0,     0,     0,     0,     0,    -2,     1,     0,    -1,     0,    -1,    -3,    -1,    -1,     1,    -1,    -2,    -2,     1,     1,     0,     1,     1,     1,     1,     1,    -2,    -3,    -1,     0,     0,    -1,     0,    -1,     2,    -1,     1,     1,    -2,    -3,    -2,     1,     1,    -2,    -1,     0,     0,     1,     1,    -1,    -1,     0,     1,     2,    -2,    -2,     0,    -1,    -1,     0,     0,    -1,     3,    -1,     1,     1,    -2,    -2,     2,     1,    -1,    -2,     0,     0,     2,     2,     2,     0,    -2,    -1,     1,     2,    -1,    -1,    -1,     0,     1,    -1,    -1,     0,     1,     0,     0,     0,    -1,    -2,    -1,    -1,    -3,    -1,     1,     2,     2,     2,     3,     0,    -1,    -1,     2,     2,    -1,    -1,    -3,    -1,     0,    -1,    -1,     0,     1,    -1,    -2,     1,    -1,    -1,    -1,    -2,    -1,     1,     0,     1,     2,     0,    -2,     0,    -1,     0,     0,     0,    -1,    -1,    -2,     0,     0,    -1,     0,     0,    -2,     0,    -3,     1,     0,    -1,    -4,    -3,     0,     1,     0,     0,     0,     0,    -1,     2,     1,     0,    -1,     0,     0,    -1,    -3,     0,     0,    -1,     0,    -1,    -2,    -3,    -1,     1,     1,    -1,    -2,    -1,     1,     0,     1,     0,    -1,    -1,    -1,     2,     0,     0,    -2,    -1,     0,    -3,    -2,     0,    -1,     0,     0,     0,    -2,     0,     0,    -1,     0,    -2,     1,     0,    -1,     1,    -2,     0,    -1,     0,    -1,     1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -1,    -1,     0,    -1,     1,     0,    -2,    -1,     0,    -1,    -2,    -1,     0,     0,     2,     1,    -1,    -2,    -1,     1,    -1,     0,    -1,     1,     0,    -1,     0,    -1,    -2,     0,    -1,     1,     0,     0,    -2,    -2,    -1,    -1,    -1,    -1,     0,     1,     1,    -1,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,     0,     0,    -1,    -2,    -1,    -2,    -1,    -3,    -1,    -1,    -1,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     1,     1,     0,     1,     2,    -2,    -1,    -1,     1,    -1,    -2,    -3,    -2,    -2,    -1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,     0,     0,     0,    -3,    -3,    -1,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -2,     0,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0),
		    47 => (    0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,     1,     0,    -3,    -2,    -3,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -3,    -2,    -2,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,    -1,    -2,    -1,     0,    -3,    -3,    -2,    -1,     0,    -1,     0,    -2,    -1,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,    -2,    -2,    -2,    -3,    -1,    -2,    -3,    -3,    -3,    -2,    -2,    -2,    -2,    -1,     0,    -1,    -1,    -3,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -1,    -3,    -4,    -3,    -1,    -1,    -3,     0,     1,     0,    -2,    -5,    -5,    -4,    -5,    -6,    -6,    -4,    -3,    -3,    -3,    -1,     0,     1,     0,     0,     0,     1,    -2,    -4,    -5,    -6,    -5,    -7,    -6,    -2,     2,     2,     1,    -2,    -4,     1,     2,     0,     1,     5,     1,     3,    -3,    -1,    -3,    -1,    -1,     3,     2,     2,     1,    -1,     2,     0,    -2,    -6,    -6,    -5,    -4,    -1,    -1,    -3,     0,     0,     1,    -2,    -4,    -2,    -2,    -1,    -1,     0,    -2,    -1,    -2,     3,    -1,     0,     0,     0,     3,     3,    -2,    -5,    -5,    -5,    -2,    -4,    -4,    -5,    -3,    -2,     1,    -2,    -2,    -4,    -1,     2,     1,     0,    -5,    -2,    -1,     3,    -1,    -1,     0,     1,     4,     0,     1,    -1,    -4,    -1,    -2,    -4,     0,    -1,     0,     0,     0,    -2,    -2,     4,     2,     5,     3,     1,    -3,     0,    -1,     2,     1,    -1,    -4,    -1,     2,     0,    -2,    -1,     0,     0,     0,     2,     1,     0,    -1,     3,     2,     2,     0,     2,     2,     0,    -2,    -1,    -3,     1,     0,     1,     0,     0,     0,     1,    -1,     3,    -1,     0,     0,     4,     3,     2,     2,     0,    -2,    -1,     0,     1,     1,     1,     1,     1,    -1,    -2,    -1,     4,     0,     0,     1,     3,     2,     2,    -2,     2,     3,     0,     1,     3,     4,     1,    -2,    -2,     2,     3,     1,    -1,     0,    -1,     2,     0,     3,     2,     5,     5,     0,     1,     2,     3,     2,     1,     1,    -3,    -1,     0,     2,     1,     0,    -2,    -2,    -2,     1,    -1,    -1,     0,     3,     2,     2,    -4,     3,     3,     2,    -1,    -1,     2,     4,     3,     1,     5,     0,    -3,     1,     2,     2,    -1,    -5,    -6,    -2,    -2,    -1,    -2,     2,     1,     2,     1,     1,     1,     0,    -1,    -3,    -1,     0,    -1,     0,     4,    -3,     1,    -1,     2,     0,     3,     2,    -3,    -8,    -7,    -4,    -1,     0,     1,     0,     3,     2,     0,    -1,    -4,    -3,    -1,     0,     0,     0,    -1,     0,     2,     5,     0,     1,     1,     0,     0,    -2,   -10,   -11,    -2,    -1,     0,     0,     0,    -3,     1,     2,     2,     1,    -2,    -4,    -5,     0,    -2,     0,     0,     2,     0,     3,     0,    -1,    -1,     0,    -3,    -6,    -8,    -6,     0,    -1,     1,    -2,    -1,    -1,    -2,     3,     2,     1,    -2,    -3,    -4,     1,    -3,     1,     0,     2,    -4,     0,    -1,     0,     2,    -1,    -5,    -8,    -4,    -2,     0,     1,     0,    -3,     0,    -1,    -1,     3,     1,     0,    -3,    -3,     0,     1,     0,     0,     3,     0,    -4,    -1,     0,     2,     1,    -2,    -6,    -7,    -2,    -1,     3,     0,    -1,     0,     2,    -2,     1,    -1,    -2,    -1,    -3,    -3,     1,    -1,     0,     0,     1,     0,    -2,    -1,    -1,    -1,    -2,    -3,    -5,    -3,    -1,     1,     0,     1,    -1,    -3,     1,    -1,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,     1,     1,     0,    -3,    -3,    -2,    -4,    -5,    -3,    -2,     0,     1,     0,     0,     0,    -2,    -2,     0,     1,     1,     0,     1,    -1,    -3,     4,     0,    -1,     0,     0,     0,    -1,    -4,    -2,    -2,    -3,    -4,    -3,     0,    -1,     0,     1,     1,    -1,     1,    -1,    -2,     1,    -2,     3,    -1,     0,    -3,     1,     0,     0,     0,    -1,     0,    -1,    -3,     0,     1,    -4,    -2,    -1,    -2,     2,     1,     1,     0,     0,    -2,     0,     0,    -1,     0,     1,    -2,    -1,    -3,     1,     0,    -1,     0,     0,     0,     0,     1,     2,     0,    -2,     0,     0,     2,     0,     2,     1,    -3,     2,     0,    -1,     0,    -2,    -3,     2,     1,    -1,    -4,     1,    -2,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     1,     0,     0,     1,     3,     2,     0,     3,     1,     2,     0,    -1,     1,    -1,     1,     0,    -4,     1,    -1,     1,     0,     0,     0,     0,    -1,     0,    -2,     0,    -2,     0,     0,    -3,     0,     4,     3,    -1,    -1,     0,     1,    -2,    -2,     0,     1,     1,     1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     1,     2,    -1,     1,     2,     2,    -1,     0,     1,     2,    -1,    -2,     1,     3,    -3,    -1,     0,     4,     4,     3,    -1,     0,    -1,     0),
		    48 => (   -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -2,    -1,    -1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -3,     0,     0,     0,    -2,    -2,     0,    -1,     0,    -2,    -2,    -2,    -1,    -1,     0,     1,     0,    -1,    -1,    -1,     0,    -1,    -2,    -3,    -2,    -2,    -2,    -2,     1,     2,     1,     0,    -1,     0,    -1,     2,     1,     0,     0,     0,     4,     0,     1,    -1,     1,     0,     0,     1,    -1,    -3,    -4,    -3,    -3,    -1,     1,    -1,    -1,    -2,    -2,     0,    -2,    -1,    -1,    -2,     2,     5,     6,     1,    -4,    -4,    -1,     2,     0,     0,     0,    -1,    -1,    -3,    -2,    -1,    -1,     0,    -2,    -1,     0,     0,    -2,     0,    -5,    -4,    -3,    -3,     1,     3,     4,     2,    -2,    -3,    -1,     0,    -1,     0,     0,    -1,    -4,    -1,    -2,    -1,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,    -3,    -2,     0,     1,     0,    -1,    -1,    -3,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -3,     0,     0,     1,     0,    -2,     0,     3,     0,     0,     1,    -1,    -3,    -2,     1,     2,     0,    -2,    -1,     1,     1,     1,     1,     0,     0,    -2,    -2,    -4,    -3,    -3,    -1,     1,    -1,     1,    -1,    -2,     1,     3,     3,     0,    -2,     1,     1,     3,     0,    -1,    -2,    -1,     1,     0,     1,     1,    -1,     1,     0,    -2,    -4,    -5,    -2,    -1,    -1,    -1,     0,    -1,     0,     1,     0,    -1,    -1,    -1,    -1,     0,     1,    -1,    -3,    -3,     0,     1,     0,     0,    -1,     1,    -1,    -1,    -3,    -4,    -2,    -1,     1,     1,    -1,     2,     3,     0,    -1,    -1,    -1,    -3,     0,    -1,     0,     0,    -1,     2,    -1,     0,     1,    -1,     0,     1,     1,    -1,    -1,     0,    -1,    -4,    -1,     2,    -1,     0,     1,    -1,    -2,    -2,    -3,    -2,     0,    -1,     0,     0,    -2,    -2,    -1,     0,    -1,    -2,    -3,    -1,     1,     3,     1,    -2,    -3,    -3,     0,     1,    -1,    -1,     0,     0,    -2,     0,     0,    -1,    -2,    -1,     0,     0,    -2,    -2,    -3,    -1,    -1,     0,     0,     1,     1,     3,     2,     1,    -3,    -2,     0,    -1,    -5,    -1,    -2,    -1,     0,    -1,    -2,    -2,     0,     0,    -1,    -1,    -1,    -3,    -2,    -2,    -4,    -3,     1,    -2,    -1,     1,     1,     1,    -1,    -2,     1,    -3,    -3,    -4,    -3,    -1,    -2,    -2,    -3,    -1,    -4,    -2,    -1,     0,    -1,     1,     0,     0,    -3,    -3,    -2,    -2,    -4,    -1,    -1,     2,     2,     2,     1,     0,    -3,    -4,    -3,    -1,    -2,    -1,    -1,    -1,    -3,    -3,    -1,    -1,    -1,     2,     0,    -1,    -2,    -3,     0,    -2,    -2,    -1,    -2,     1,    -2,    -1,    -1,     0,    -3,    -1,    -2,     1,    -2,    -2,    -1,    -2,    -3,    -3,     0,    -1,    -2,     2,     0,    -2,    -3,    -3,    -5,    -5,    -1,     0,     1,     2,    -2,    -1,    -3,     0,     0,    -2,     1,     1,     3,    -1,    -2,     0,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -2,    -4,    -3,    -3,    -2,     0,     1,     3,    -1,     0,     1,    -1,     2,     1,     1,    -1,     0,     1,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -3,    -1,    -1,     0,     3,    -2,     0,     2,    -3,     3,     3,     1,    -1,    -1,     0,     1,    -2,    -1,    -2,    -1,     1,     1,    -1,    -1,    -2,    -1,    -4,    -3,    -2,     0,     2,     2,     2,    -1,    -2,     0,    -4,     3,    -2,     2,     1,     0,     0,     0,    -1,    -1,    -3,     0,    -1,     0,    -1,    -1,    -2,    -2,    -5,    -4,    -2,    -1,     1,     2,     1,    -2,    -1,     0,     0,     0,     0,     2,     0,     1,     1,     1,    -3,    -1,    -2,     0,    -1,     0,    -1,     0,    -1,    -2,    -6,    -5,    -4,    -3,     0,     0,    -1,     1,    -1,     0,    -1,    -3,    -1,     0,     0,     3,     1,    -2,    -2,     0,    -2,    -1,     0,     1,    -1,    -2,    -1,    -1,    -2,    -2,    -4,    -3,    -1,    -2,     0,    -1,     0,     1,     0,     1,    -2,     0,     3,     1,     2,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -4,    -4,    -4,    -2,     0,    -1,    -3,    -4,    -2,    -1,     2,    -2,     1,     0,     3,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,    -2,     0,    -2,    -2,    -1,    -4,    -3,    -3,    -2,    -3,    -2,    -2,     0,     3,     4,     2,     2,     1,     1,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -2,     0,    -1,    -2,    -1,    -1,    -2,    -4,    -2,    -2,    -3,    -4,    -3,    -2,    -1,    -1,    -4,    -4,    -2,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,    -1,     0,    -1,     1,     0,     1,     0),
		    49 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,     0,    -5,    -4,    -4,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,    -2,    -1,    -1,    -3,    -1,    -1,    -4,    -2,    -3,    -1,     0,    -1,    -2,    -1,    -1,    -2,     0,     1,     0,     0,     0,     1,     0,    -5,    -1,    -1,    -1,    -3,    -3,    -4,    -4,    -4,    -7,    -5,    -6,    -6,    -5,    -3,     1,    -3,    -3,    -2,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,    -2,    -4,    -5,    -4,    -3,    -5,    -4,    -7,    -8,    -2,    -5,    -3,    -2,     0,     2,    -8,    -4,    -6,    -3,    -1,    -1,    -3,    -3,    -1,     0,     0,    -1,    -2,     0,    -2,    -4,    -3,    -3,    -3,    -2,     1,    -1,     2,    -2,    -1,    -3,    -3,    -3,    -2,    -1,    -2,    -5,    -5,    -3,    -3,    -2,     0,     0,    -1,    -1,    -5,    -5,   -11,    -6,    -1,     0,     5,     1,     2,    -1,     4,     0,     0,     1,     2,     2,     0,     2,     1,    -3,    -3,    -5,    -5,    -3,    -2,     1,    -3,    -4,    -5,    -9,   -11,    -1,    -3,    -1,     1,     2,     2,     3,     1,    -1,     3,     0,     2,     1,     0,    -1,     0,    -2,    -5,    -5,    -4,    -3,    -1,    -5,    -3,    -3,    -3,    -5,     0,     0,    -3,     0,    -1,    -1,     0,     0,    -2,     0,    -2,     0,    -1,     1,    -1,     0,     2,    -2,    -2,    -3,    -5,    -4,    -2,    -1,    -2,     0,    -2,    -5,     0,    -1,     0,    -1,    -2,     0,     1,     0,    -1,    -2,     3,    -1,    -1,    -2,     1,     0,     2,     0,    -1,    -2,    -4,    -5,    -2,    -1,    -3,    -5,     0,     1,     1,    -2,    -2,    -1,     1,    -1,     1,     1,    -2,    -2,    -2,    -1,     1,    -1,     1,     2,     1,     1,    -1,    -2,     6,    -5,    -3,     0,    -8,     2,    -1,     3,    -1,    -1,    -1,     1,    -1,     3,     0,     0,     1,    -2,    -1,     0,     3,     1,     1,     2,     2,     4,    -2,     1,     6,    -4,    -4,    -1,    -2,     1,     1,     5,     1,     1,     2,     0,     3,     0,     2,    -3,    -4,     1,     0,     1,     3,     4,     4,     1,     3,     3,     5,    -5,    -9,    -6,    -1,     0,    -4,    -3,     1,     6,     5,     2,     4,     3,     2,     2,     0,     1,     1,     2,     2,     4,     0,     2,     3,     3,     2,     7,     1,    -8,    -5,    -3,     0,    -1,    -3,    -2,     1,     5,     4,     1,     2,     4,     1,     3,    -1,    -2,     1,    -1,     0,     3,     0,     2,     3,     0,     1,     7,     0,   -11,    -7,    -1,     0,    -1,     0,    -6,     1,     4,     0,    -2,     2,     5,     3,     0,    -3,    -2,     1,    -2,     2,     2,     4,     3,     3,    -1,    -3,     0,    -3,   -10,    -6,     2,    -1,     0,    -1,    -5,    -3,     1,    -3,     0,     0,    -1,    -3,     3,    -3,    -1,    -1,    -1,     0,    -1,     0,     0,    -2,    -1,    -5,    -1,    -2,    -8,    -4,    -1,    -3,     0,     0,    -6,     0,    -2,    -2,    -2,     1,     0,    -1,    -1,    -4,    -1,    -2,    -2,     1,     1,     1,    -2,    -3,    -3,    -2,    -2,    -2,    -7,     0,    -1,    -2,     3,     0,    -6,     1,    -2,    -4,    -2,    -1,     0,    -1,     1,    -1,    -2,    -4,     0,    -1,    -1,     0,     1,     0,    -3,     1,     0,    -5,   -12,    -1,    -3,    -2,     0,    -1,    -3,     4,    -2,    -4,    -4,    -4,    -3,    -3,    -3,    -2,    -3,    -7,    -1,     0,    -2,    -2,    -1,     1,     0,    -2,     2,    -3,    -5,    -1,    -2,    -1,     1,     0,    -6,     3,    -2,     3,    -2,    -8,    -6,    -4,    -5,    -1,    -4,    -4,     1,    -2,     1,     1,    -2,     1,    -3,    -2,    -1,    -1,     1,     2,    -1,     0,     0,     0,    -6,     4,     1,     4,    -2,    -3,    -4,    -3,    -5,    -4,    -4,     0,    -5,    -2,     1,    -2,    -3,    -2,    -4,    -1,    -2,    -4,    -2,     2,   -10,     0,     1,    -1,    -5,     3,    -3,    -1,     1,     3,     3,     0,     1,    -2,    -1,     0,     0,     1,    -1,    -2,    -3,    -4,    -2,    -1,    -1,    -4,     0,    -1,    -6,    -1,     0,     0,    -4,     3,    -1,    -2,    -2,     1,     0,    -2,     0,    -2,    -2,     0,     0,    -3,    -2,    -2,    -2,    -1,     0,     2,     2,    -1,     0,     0,    -1,     1,     0,     0,    -4,    -4,    -1,     2,    -3,     1,    -1,    -1,     1,     2,    -1,    -2,    -4,    -1,     1,    -3,     0,     1,    -2,     0,     3,     4,     0,    -1,    -2,     0,     0,     0,     3,    -3,     4,     2,    -5,    -6,    -2,    -1,    -4,    -3,     1,     0,     4,     0,     2,     3,     3,     2,     4,     5,     1,    -1,    -2,     0,    -2,     1,     0,     0,     0,     2,     3,     0,     1,     0,     1,     1,    -2,    -1,     3,     1,     4,     1,     2,     4,     6,     1,     4,     4,     2,     2,     2,     1,     1,     0,     0,     0,     0,     0,    -3,    -4,     1,     1,     2,     1,    -1,     1,     0,    -2,     3,     2,     1,    -5,    -2,     3,     0,    -3,     1,    -3,     0,     0,     0,     0),
		    50 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     1,     0,     0,     0,    -1,     1,     0,     1,     0,     0,     1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     2,    -1,    -1,    -1,    -1,    -2,    -2,    -4,    -4,    -4,    -2,    -3,    -2,    -2,    -1,     0,     1,     0,    -3,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     1,    -1,    -1,    -4,    -4,    -1,     0,     0,     2,     0,    -3,    -4,    -2,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     0,     0,    -1,    -4,     2,     0,     2,     3,     1,     2,    -1,     0,     0,    -3,    -1,     1,     1,     0,    -3,    -4,    -1,     0,    -1,     0,    -1,     0,     0,     0,     0,     1,     1,    -2,     0,    -1,    -4,    -1,     1,     2,     1,     2,     1,     0,     2,     0,     1,    -1,    -1,    -1,     0,    -1,    -2,    -3,    -2,    -3,     0,     0,    -2,    -1,     1,    -1,     0,    -2,    -2,    -1,     1,     1,     0,     0,     0,     1,     3,     1,     1,    -1,    -1,    -3,    -1,     4,     2,    -3,    -3,    -1,     0,    -1,    -2,    -1,    -1,     2,     1,     1,    -1,     1,     3,     1,     1,     0,     1,     0,     0,     2,     0,    -1,    -3,    -2,    -2,     2,     2,    -2,    -3,     1,     1,     0,     0,    -2,    -2,     0,     0,     0,     2,     2,    -1,     0,     3,     2,     2,    -1,     0,    -2,     0,    -2,     0,    -1,     1,     0,     1,    -2,    -3,    -1,     0,     0,     0,    -1,    -3,     3,    -2,     0,     0,     1,     0,     0,    -1,     0,     0,     0,    -2,    -3,     3,     3,     3,     1,     2,     0,     3,    -4,    -3,     0,     0,     0,     0,    -1,    -4,     0,     0,     0,     1,     1,     2,     0,    -4,    -2,     0,    -1,    -2,     1,     2,    -1,    -2,    -1,     3,     1,     3,    -3,    -2,     0,     0,     1,    -2,    -2,    -3,     0,     1,     0,     0,     1,     2,    -3,    -4,    -4,    -3,    -4,    -1,     0,     0,    -3,    -2,    -3,    -2,     1,     2,    -1,     0,    -1,     1,     0,     0,    -1,     0,    -2,     1,    -1,     0,    -1,    -2,    -1,    -3,    -2,    -2,    -3,    -2,    -1,    -2,     1,    -1,    -1,     0,    -4,     0,    -1,    -3,    -1,     0,     1,     0,     1,     3,     0,     0,     0,     3,     1,    -2,    -5,    -5,    -7,    -6,    -4,    -3,    -3,    -1,    -2,     0,     0,     1,    -2,     0,    -1,    -1,    -1,     0,     0,     0,    -2,    -2,     3,     2,     3,     1,     1,    -2,    -7,    -5,    -6,    -2,    -4,    -5,    -4,    -1,     0,    -2,     0,    -1,     2,     3,     0,    -2,     0,     1,     0,     0,    -4,     1,     3,     3,    -1,     0,     2,     2,    -4,    -8,    -5,    -2,    -2,    -3,    -3,    -2,     0,    -1,     1,     0,    -1,     1,     0,     0,    -2,     1,     0,     0,    -5,     2,     3,     0,     4,    -2,    -1,     1,    -2,    -2,    -4,     0,    -3,    -6,    -5,    -4,    -3,     1,     3,     1,     0,    -1,    -1,    -2,     0,     0,     0,    -1,    -1,     2,     2,     1,     0,    -1,    -1,     2,     3,     1,     1,    -1,    -6,    -8,    -4,    -6,    -3,    -1,    -1,    -1,     0,    -2,    -2,    -3,     0,     0,     0,    -1,     1,    -2,     2,     4,     2,     1,     1,    -1,    -1,     0,    -2,    -4,    -5,    -6,    -3,    -1,    -1,     3,     2,     1,     1,     1,    -2,    -2,    -1,     0,     0,     0,     1,     0,     2,    -1,     1,     1,    -1,    -1,    -1,     1,    -1,    -1,    -3,     0,     2,    -3,     0,     1,     2,     2,     0,     0,    -2,     0,    -1,     0,     0,     0,     1,     3,     4,    -2,     0,    -2,    -3,    -2,     1,     1,    -1,     0,     0,     1,     1,     1,     0,     1,     2,    -1,     0,     1,    -2,    -1,     0,     0,    -1,     0,     3,     4,     1,     3,     1,    -3,    -1,    -2,     0,    -2,    -1,     2,     2,    -2,     0,     0,     0,     0,     2,     3,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,     1,     2,     2,     3,     2,    -1,     1,    -1,     0,     0,     1,     1,     1,     1,     0,    -1,     0,    -1,     1,     1,    -2,     0,     0,     1,     0,    -1,     0,    -3,    -3,     1,    -1,    -2,     0,     0,     1,     0,     2,     0,    -1,     2,     0,     2,     0,     0,    -3,    -3,    -1,    -1,    -5,     0,    -1,     0,     0,    -1,     0,    -1,    -2,     0,     1,     1,    -1,     2,     3,     1,     1,     2,    -2,     1,    -1,     2,     1,     2,    -3,    -3,    -3,    -1,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -3,    -2,    -2,    -3,    -5,    -6,    -6,    -7,    -5,    -4,    -4,    -2,     0,    -1,     0,     1,     0,     0,    -1,     0,     0,    -1,    -1,    -2,    -1,     0,    -2,    -1,    -2,    -1,    -3,    -3,    -5,    -4,    -3,    -4,    -4,    -3,    -4,    -2,    -3,     1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -3,    -2,    -3,    -1,     1,     1,    -1),
		    51 => (   -1,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -4,    -3,    -2,     1,    -3,    -1,     4,     1,    -4,    -4,    -1,    -2,    -2,    -1,    -1,     1,     0,    -1,     0,     0,     6,     3,     0,    -3,    -2,    -1,    -1,    -2,    -3,    -5,    -3,     0,    -2,    -3,    -1,    -2,    -1,     4,     4,    -3,    -1,    -2,    -1,     0,     1,     0,     0,     0,     5,     5,     0,    -3,    -2,    -1,    -1,    -3,    -4,    -2,     0,     3,     2,     0,    -3,    -4,     2,     1,     1,    -1,    -1,    -1,     0,    -1,    -2,    -2,     0,     0,     5,     3,     1,     0,     0,    -2,    -6,    -6,    -1,     0,    -2,     1,     0,     0,     2,    -4,    -2,    -1,    -3,    -2,    -1,     0,    -1,    -1,    -2,    -2,     0,     0,    -2,     1,     0,    -1,    -2,     0,    -5,    -7,    -3,     0,     1,     3,     1,    -2,     0,    -4,    -1,    -4,    -4,    -1,     0,     0,     0,     0,    -2,    -2,     0,    -1,    -2,     1,     0,    -3,    -3,    -1,    -7,    -4,     0,     1,     2,     3,     1,    -1,    -2,    -3,    -1,    -7,    -3,    -2,     0,     0,     0,    -1,    -4,    -2,     0,    -1,    -2,     1,    -1,    -2,    -3,    -3,    -7,    -3,     0,     0,     1,     2,     4,     2,    -3,    -3,    -2,    -7,    -2,    -2,     1,     0,    -1,     0,    -2,    -1,     0,    -1,    -2,    -1,    -1,     0,    -2,    -1,    -4,     0,     1,    -1,    -3,     0,     4,     3,    -3,    -5,     0,     0,    -3,     0,     1,     0,    -2,    -1,    -2,    -3,     0,    -1,    -1,    -1,    -2,    -1,    -4,    -2,    -1,    -3,     3,     0,    -1,     2,     2,     0,    -1,    -4,    -3,     0,    -1,    -5,     0,     2,    -3,    -1,     1,     3,     0,     1,     0,    -1,    -1,    -2,    -4,    -2,    -4,    -3,    -1,     2,    -1,     0,     3,    -1,     0,    -2,    -4,    -1,     2,    -1,     2,     2,    -2,    -2,    -1,     5,     1,     0,    -5,     2,     0,     0,    -1,    -2,    -1,     3,     1,     0,     1,     0,     2,    -1,     0,    -4,    -5,    -2,     4,     0,     1,     2,    -3,     0,     0,     4,     0,     0,    -5,     0,     0,    -1,     0,     1,     3,     2,    -5,     1,     1,    -2,    -1,    -2,    -1,    -3,    -3,     1,     4,    -2,    -2,    -4,    -3,     3,     2,    -1,     0,     0,     0,     0,     0,    -2,     0,     2,    -1,    -2,    -4,    -3,     1,     0,    -1,    -2,     1,     0,     0,     0,     1,    -2,    -3,    -1,     0,    -1,     3,     1,     0,     0,     0,     2,     0,    -3,    -2,     0,    -1,    -2,    -2,     4,     2,     3,     1,    -3,     0,     0,     2,    -1,     3,    -1,    -3,    -1,    -3,    -2,     0,    -2,     0,     0,     1,    -2,     0,    -2,    -1,     0,    -1,    -2,    -1,     2,     1,     0,     1,    -2,    -2,    -1,     1,    -2,     0,    -1,    -2,    -2,     0,    -3,     0,    -1,     0,     1,     0,    -1,    -1,    -3,    -2,    -3,    -1,    -2,    -2,    -1,     1,     0,     1,    -1,    -2,    -2,     1,    -3,    -3,    -2,     1,     1,    -2,    -3,    -1,     1,     0,     0,    -1,    -1,    -2,     0,    -2,    -1,    -3,    -2,    -6,    -1,    -2,     4,     2,     0,     0,    -1,     2,    -4,     1,    -1,    -3,    -3,    -3,     0,     0,     3,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,     1,    -3,    -3,    -1,    -1,     2,     3,     2,     0,    -2,    -1,    -5,    -2,    -2,    -5,    -3,    -1,     2,     2,     3,     1,     1,     0,    -2,    -2,    -1,    -2,    -4,    -1,    -1,    -1,    -1,     3,     1,     1,     1,     0,    -1,    -1,    -2,     0,    -4,    -6,    -2,     0,    -1,     3,     0,     1,     1,     0,    -1,    -2,    -1,    -3,    -6,     0,     0,    -2,     0,     0,     0,    -1,     0,    -1,    -4,     3,    -1,     1,    -1,    -4,    -4,    -2,     1,    -1,     0,     1,     1,     1,     0,    -1,    -1,    -1,    -5,     0,     0,    -1,    -2,    -1,     0,     0,    -1,    -1,    -1,     1,     1,     2,     0,    -4,    -2,    -3,     2,     2,     0,     0,     0,    -1,    -2,    -1,     1,     2,    -2,     1,     4,     0,     2,    -1,     0,     0,     0,     1,     4,     3,     1,     2,    -1,    -1,    -2,    -2,    -1,     5,     0,     0,     0,     0,    -1,    -1,    -1,     3,     1,     0,     1,     3,     4,    -1,    -3,    -3,    -4,    -5,    -2,    -4,    -3,    -2,    -1,    -4,     0,    -2,     3,     3,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -8,    -6,    -5,    -4,    -1,    -5,    -5,    -5,    -4,    -5,    -8,    -3,    -2,    -2,     0,     0,    -1,     0,     0,    -1,     0,     0,    -2,    -4,    -3,    -2,    -2,    -2,    -2,    -2,    -4,    -4,    -4,    -4,    -3,    -3,    -1,    -2,     0,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1),
		    52 => (    0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,    -1,     1,     1,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     1,    -1,     1,     1,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     1,     1,     0,    -3,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,     1,    -1,    -1,     2,     4,     4,     2,     2,    -1,     0,    -2,    -5,    -3,     0,     1,     0,     1,    -1,     1,     2,     1,    -1,     0,     0,     0,    -1,    -4,    -3,    -3,    -1,    -2,     1,     1,    -1,    -1,    -1,     1,     2,    -1,     0,     0,    -1,     3,    -1,    -1,    -1,    -5,    -2,     1,    -1,     0,     0,     0,    -1,    -1,     3,    -1,     0,     0,     0,     1,    -1,     0,     2,     1,     0,     1,    -2,     1,    -2,    -1,     2,    -2,    -1,    -4,    -4,     2,    -3,    -2,     0,     0,     0,    -1,     0,    -4,    -4,    -5,    -3,     0,     3,     0,    -2,     2,     1,     1,    -2,     1,    -1,     0,     0,     1,     0,     2,    -4,     4,    -3,     0,     0,     0,     0,     4,     3,    -3,    -2,    -1,     1,     2,     2,     0,     0,     3,     1,     0,    -1,     1,     0,     0,    -1,    -3,    -1,    -1,     0,    -3,    -3,     0,     0,     0,    -1,     5,     4,     3,    -1,     1,    -1,     0,    -1,     1,     1,     2,     0,     2,     2,     2,     1,     2,    -1,    -2,     3,     0,    -3,    -3,    -2,    -2,    -2,     3,    -1,     4,     2,     2,    -3,    -1,    -1,     2,     0,    -1,    -1,    -2,    -1,     0,     2,     3,     0,     3,    -2,     0,     3,     3,    -7,    -4,    -3,    -2,     1,    -1,     1,     1,    -1,     1,    -2,    -2,    -1,     2,    -2,     0,     1,    -3,    -1,     1,     1,     1,    -1,     3,     0,    -2,    -2,     3,    -6,    -4,    -2,    -1,     0,     0,     0,     2,    -4,     4,     2,     0,    -1,     0,    -2,    -3,     0,     2,    -1,    -1,    -1,    -1,     0,     1,     2,     0,    -1,     3,    -1,    -1,     1,    -1,     0,    -2,    -1,     3,     0,     1,     2,     0,    -1,    -3,    -5,     0,    -2,    -3,    -4,    -3,     0,    -1,    -3,    -1,    -1,     0,    -1,     1,     0,     0,    -3,    -1,     0,     0,    -4,     0,     1,    -4,    -2,    -3,    -4,    -3,    -3,    -3,    -1,    -5,    -6,    -2,     0,    -1,    -3,    -1,    -2,    -1,    -1,    -2,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -5,    -5,    -8,    -5,    -4,    -5,    -6,    -3,    -3,    -1,    -1,    -3,    -2,    -3,    -2,    -3,     1,    -2,    -1,     2,     3,    -1,     0,    -2,    -2,    -1,    -3,    -6,    -6,    -6,   -10,    -6,    -3,    -3,    -1,    -2,     0,    -1,    -4,    -1,    -1,    -1,    -3,    -4,     0,    -5,     0,     0,     3,     2,     0,    -2,     0,    -1,    -6,    -3,    -3,    -4,     1,     0,    -2,     2,     0,     2,     1,    -3,     0,     0,    -4,    -4,    -4,    -2,    -5,    -2,     1,    -1,     4,     5,     0,     0,    -2,    -4,    -7,    -2,    -3,    -2,    -1,     1,     1,     1,    -2,     1,     1,    -1,    -2,    -1,    -2,    -4,    -3,    -1,     2,    -1,     2,     4,     5,     3,     0,     0,     0,    -3,    -2,    -3,     0,    -1,     0,     0,     2,     1,    -2,     4,     2,     0,    -1,    -1,    -1,    -3,    -2,    -1,    -1,    -1,    -3,     6,     4,     3,     0,     0,    -1,    -5,    -2,    -1,     2,     2,    -1,    -2,     0,     0,     1,     0,    -1,    -1,    -1,     2,    -2,    -2,    -3,     2,     2,     2,     5,     8,     0,     4,     0,    -1,     1,    -3,    -3,    -1,     2,     2,    -2,    -2,     1,     1,     0,     5,     4,     1,     2,     0,    -1,    -2,     0,     2,     1,     2,    -1,     2,     2,     4,     0,    -1,     2,     0,     0,    -2,     6,     2,     1,     2,     4,     3,     2,     6,     2,     2,     4,     0,    -1,    -1,     4,     4,     1,     1,     1,     3,     1,     0,     0,     1,     1,     3,     1,     1,     3,     2,    -1,     2,     1,     1,     0,     5,     4,     3,     2,     3,     1,     2,     2,     2,     3,     6,     3,     3,     3,    -1,     0,     0,     0,     0,     0,     3,     4,     2,     1,     3,     1,     1,     1,     0,     2,     1,    -1,    -3,     0,    -3,     1,     3,     5,     5,     4,     0,    -4,    -1,    -1,     0,     0,    -3,    -2,     1,     3,     2,     1,     3,     1,     4,     3,     2,     1,    -1,    -3,    -2,    -2,     0,     2,     3,     6,     4,     3,     0,    -2,     0,     0,     0,    -3,    -2,    -1,    -2,     0,     2,     4,    -1,     0,     0,     3,    -1,     2,     1,    -3,    -1,     0,     0,    -3,    -2,     0,     3,     7,     4,     2,     0,     0,     0,    -2,     0,    -3,    -6,     3,    -1,    -3,    -6,    -8,    -2,    -1,    -1,     3,     2,    -2,     1,    -4,    -6,    -1,     1,    -5,    -2,     1,     3,     2,     0,     0,     0,     0,     0,    -2,    -4,    -4,    -3,    -3,    -4,    -7,    -6,    -3,    -4,    -4,    -2,    -6,    -5,    -4,     0,    -2,    -2,    -1,     0,    -1,     0,    -1,     0,    -1,     1,    -1,     0,     0,     0,    -1,     0,     1,     0,    -2,    -3,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0),
		    53 => (    0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     1,     0,     0,     1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -3,     2,     3,     2,    -1,    -2,    -2,    -4,    -4,    -3,    -1,     0,    -2,    -2,    -3,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     1,     1,    -1,     2,     2,     1,     2,     0,    -2,     1,     2,     2,    -1,    -1,    -1,    -1,    -5,    -2,     0,     0,     0,     0,     1,     0,     0,    -1,     1,     1,     2,     1,    -1,    -1,    -2,    -3,    -3,     0,    -1,    -1,    -4,    -2,     0,    -2,    -2,     2,    -5,    -4,    -2,    -1,     0,     0,     0,     1,    -1,    -1,     2,     2,     4,     0,    -3,    -4,    -2,    -1,    -2,     0,    -1,     0,    -1,    -1,     1,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -1,     0,     1,     0,     1,     0,     0,     0,    -1,    -3,    -2,     2,    -1,     0,    -1,    -2,    -1,    -1,     0,     0,    -3,    -2,    -1,    -1,    -1,    -1,    -4,    -2,    -1,     1,     1,     2,    -2,    -6,    -2,     0,    -2,    -3,    -1,    -1,     0,    -1,     0,     0,     0,    -1,     1,     0,    -3,     1,    -2,     0,    -2,    -1,    -3,    -2,    -1,     0,    -1,     2,    -3,    -5,     0,    -2,    -3,    -1,     1,     1,    -1,     0,    -2,     0,    -1,     0,     0,     2,     1,     1,     3,     2,    -4,    -7,    -2,    -3,     0,     0,    -3,    -2,    -3,     0,     0,     2,     0,    -1,    -1,     1,     2,     3,     2,     2,    -1,    -2,    -1,    -2,    -1,     2,     1,     1,    -3,    -9,    -4,    -4,    -1,     0,    -3,    -1,     2,     1,     1,     4,     0,     5,     2,     3,     2,     0,     0,    -1,    -2,    -4,     0,     2,     2,     1,    -1,     2,    -1,    -8,    -1,    -3,     0,     0,    -3,    -1,     5,     4,     4,     1,     2,     1,     3,     1,    -2,    -5,    -5,    -4,     1,     1,     1,     2,     3,     4,     1,     1,     0,    -5,    -5,    -1,    -1,     0,    -3,    -3,     5,     3,     2,     0,     1,    -3,    -3,    -4,    -9,    -6,    -1,     2,     4,     1,     0,     2,     0,    -1,    -2,    -1,    -3,     0,     0,     0,     0,     0,    -2,    -6,     2,    -3,    -2,    -1,    -2,    -4,    -8,    -9,    -5,    -1,     1,     3,     1,     1,     0,    -2,    -2,    -2,    -1,    -4,    -3,     3,    -2,    -1,     0,    -1,     1,    -1,    -2,    -4,    -5,    -7,    -6,    -6,    -3,    -1,    -2,     1,     2,     1,     1,    -1,     1,    -3,    -2,    -3,    -2,    -5,    -1,     4,    -1,    -2,    -1,     0,     2,     1,     1,    -1,    -2,    -5,    -7,    -5,     0,     1,    -1,     2,     3,     5,     0,     2,    -1,    -1,     0,    -1,     0,    -2,    -1,     3,    -1,     3,     1,     0,     0,     2,     3,     1,    -2,    -3,    -2,    -4,    -3,    -3,    -6,    -1,     0,    -1,    -3,     2,     1,    -2,     0,     0,     4,    -1,    -3,     2,    -3,     1,     0,     0,     0,     1,     1,     0,     0,    -1,    -3,    -5,    -7,    -9,    -9,   -11,    -9,    -6,    -4,     2,    -1,    -3,     2,     2,     3,     1,    -2,    -1,    -4,    -1,     0,    -1,     0,     4,     1,     4,     0,    -2,     0,    -1,    -4,    -4,    -6,    -9,    -7,    -4,    -4,     0,     3,     2,     2,     1,    -1,     1,    -1,    -6,    -2,     0,    -1,     0,    -2,    -2,    -2,     1,     2,     0,     0,    -2,     1,    -1,    -2,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     1,     0,     3,     0,    -2,     1,    -1,    -1,     0,     0,    -2,     0,     1,     2,     2,     2,     1,     3,     2,     4,     2,     0,    -1,    -3,    -1,    -2,    -2,     0,     2,     0,     1,    -2,    -3,    -2,    -1,    -1,     0,     1,    -1,     0,    -1,     1,     1,     2,     3,     1,     0,     0,     0,    -1,     0,    -2,    -2,    -3,    -1,     1,     2,     0,    -1,    -2,    -3,    -1,    -1,     0,    -1,     0,    -2,     0,     0,    -1,    -2,    -2,     0,    -1,     1,     0,     1,     1,     1,    -1,     0,     0,     0,     2,     0,     1,    -3,    -3,    -3,    -1,    -1,     0,     0,     0,     2,     2,     3,     2,    -1,    -1,    -1,    -1,    -3,    -1,    -2,    -1,    -1,     2,     0,     2,     2,     0,     1,     1,    -3,    -3,     2,     2,     0,     0,     0,     0,     0,     2,     3,     0,    -2,    -1,     0,     2,     0,     1,     1,     0,     0,    -1,     2,     2,    -1,    -3,    -1,    -1,    -2,    -4,    -3,    -2,    -1,     0,     0,     0,     0,    -3,    -2,     1,     2,     1,    -1,    -1,    -4,    -4,    -3,    -6,    -4,     0,     0,    -3,    -3,    -3,    -2,    -2,    -2,    -3,     0,     0,     0,     0,     0,     0,     0,    -2,    -5,    -4,    -3,    -4,    -5,    -4,    -6,    -5,    -4,    -2,    -2,    -2,    -3,    -6,    -6,    -5,     0,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -3,    -2,    -3,     0,    -2,    -2,    -3,    -2,    -2,    -2,    -3,    -1,    -1,     0,     0,     0,     0,     1,     0),
		    54 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     0,     1,     1,     0,    -3,    -2,    -1,     0,    -1,     0,    -1,     1,     2,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     1,     0,     0,    -1,     0,     0,    -1,    -4,     0,    -2,    -3,    -4,    -1,    -1,    -1,    -1,    -3,    -2,    -3,    -5,    -2,    -1,    -1,    -3,    -2,     0,    -1,     0,    -2,     0,     0,     0,     0,    -1,    -2,    -3,    -1,    -2,    -3,    -1,    -1,    -1,    -1,     0,    -1,    -2,     0,     0,     2,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,     2,     4,     2,    -2,    -5,    -6,    -4,    -3,    -3,    -5,    -6,    -6,    -4,    -2,    -1,     0,     5,     4,     2,    -5,    -1,    -1,     0,    -1,     1,    -2,     0,    -2,     1,     5,     2,    -3,    -6,    -4,    -2,     6,     3,     2,    -1,    -6,    -7,    -3,    -2,     0,     2,     1,    -2,    -1,    -1,     0,     0,    -1,    -2,     2,     3,    -1,     2,     2,    -2,    -7,    -8,    -1,     1,     1,     3,     3,     1,    -6,   -11,   -10,    -1,     3,     4,     2,    -5,     1,    -4,     0,    -2,     0,    -2,     1,     2,     1,     2,     0,    -1,    -4,    -2,    -4,     0,     3,     3,     2,     2,    -8,   -11,    -5,     1,     5,     5,     1,    -6,     0,    -4,    -1,    -2,     0,    -3,     0,     3,     2,     2,    -1,    -1,    -3,    -4,    -5,     0,     2,     4,    -2,    -6,   -10,    -5,    -1,     3,     2,    -1,     0,    -2,     1,    -3,     0,    -1,    -1,    -3,     1,     0,     2,     4,     0,    -2,    -3,    -5,    -2,     0,     3,     2,    -1,    -5,    -5,    -2,     2,     2,    -1,     1,    -1,    -1,     1,    -3,     0,    -1,    -3,    -3,    -1,     0,     1,     0,    -3,     1,    -1,    -4,     1,     0,     3,     1,    -1,    -3,    -3,     0,     1,     0,     0,    -2,     0,     1,    -1,    -2,    -1,     0,    -3,    -2,    -2,     1,    -1,    -1,     0,     2,     0,     1,     1,    -3,     0,     0,    -2,    -3,    -2,    -1,     0,     0,     1,     0,    -2,     0,    -2,    -4,     0,     0,    -2,    -7,    -2,     1,    -1,     0,     1,     1,     2,    -3,     1,     1,     0,    -2,    -2,    -2,    -3,     0,     1,     1,     0,    -3,    -1,    -2,    -5,    -4,     0,     1,    -2,    -4,    -3,     0,     0,     1,     0,     1,     4,     0,    -3,     2,    -3,    -2,     1,     0,    -1,     2,     0,     0,     0,    -1,    -3,    -4,    -5,     0,     0,     0,    -2,    -4,    -1,     0,     2,     0,     0,     1,     2,     0,     0,     2,     1,    -1,     0,     2,    -1,     0,     1,     1,     2,    -2,     0,    -3,    -1,     0,     0,     0,     0,    -4,     0,     1,     1,     3,     2,     2,     2,     1,     1,     0,     1,    -1,    -2,     0,     0,     1,    -1,    -1,     0,     0,    -2,    -2,    -1,     1,     1,     0,    -1,    -3,    -2,     1,     3,     4,     2,     0,    -2,    -1,     0,     0,     0,     3,     1,     0,    -1,     0,     1,    -1,    -3,    -2,    -1,    -1,    -4,    -1,     0,     0,    -1,    -2,    -1,     0,     1,     0,     2,    -1,     0,    -1,     0,     0,     2,     1,     1,    -1,    -1,    -2,    -1,    -1,     0,    -2,    -3,    -3,    -2,    -1,    -2,     0,     0,     3,     2,    -1,    -2,    -2,    -2,     1,    -4,    -4,    -2,     0,     2,    -1,    -1,    -2,    -1,    -3,    -4,    -2,    -2,    -3,    -1,    -2,    -1,    -2,    -1,    -1,    -2,     4,     1,    -6,    -4,    -2,    -1,    -1,    -6,    -3,    -2,    -3,     0,    -1,    -1,    -1,     1,    -2,    -3,    -4,    -3,    -3,     0,    -2,    -1,    -1,     0,     0,     0,    -2,     0,    -2,    -2,    -2,    -3,     1,    -3,     0,     0,    -3,     3,     0,    -2,     0,     2,    -2,    -6,     0,    -1,    -1,     2,    -3,    -1,     0,     0,     0,    -1,    -5,    -3,     0,    -3,    -4,     1,     1,     0,     1,    -1,    -5,     0,    -2,    -1,    -1,     1,    -1,    -4,     0,    -1,     1,     0,    -3,    -2,     0,     0,     0,     0,    -3,    -3,     1,    -1,     1,     2,    -2,    -1,     0,    -1,    -3,    -1,    -2,     1,    -2,     0,     3,    -1,     0,     1,    -1,     2,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -4,    -1,     1,     1,     0,     4,     2,     1,    -3,    -2,    -3,    -3,    -2,     0,     1,     2,     0,    -1,     0,     1,     2,     0,     0,     0,    -1,     0,     0,    -4,    -3,     1,     1,     1,     1,     0,     3,     2,    -2,    -1,     0,    -5,     0,     1,     1,     3,     0,     2,     1,     0,     3,     0,     0,     0,     0,    -1,     0,    -2,    -5,     1,     0,     0,     0,     2,     2,    -5,    -7,    -2,     0,    -4,     1,    -2,    -4,     0,     0,     2,     0,    -1,    -1,     0,     0,     0,     0,     0,    -3,    -1,    -3,    -3,    -1,    -2,    -3,    -4,    -3,    -3,    -4,    -1,     0,    -1,     1,    -3,    -4,    -4,    -5,    -4,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,    -3,    -2,    -2,    -2,    -4,     0,    -2,    -3,    -3,    -2,    -3,    -2,    -3,     0,     0,     0,     0,     0),
		    55 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -2,    -1,    -1,    -2,    -3,    -3,    -3,    -2,    -3,    -4,    -4,    -1,     0,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -2,    -2,    -3,    -5,    -4,    -5,    -6,    -8,    -4,     1,     2,     2,     1,    -1,     0,    -3,    -3,    -1,    -3,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -3,    -6,    -4,    -8,     2,     3,     0,     1,     0,    -2,    -4,    -3,     0,     2,     4,     0,     3,     0,    -3,    -1,     2,     5,     0,     0,    -1,    -2,     0,    -3,    -1,     0,     1,     0,    -1,     1,     0,     1,    -2,    -1,    -2,    -3,    -2,     2,    -3,    -3,     0,    -2,    -1,     5,     3,     1,    -2,     0,     0,    -2,     0,    -3,    -1,    -2,     0,    -2,     0,     0,     4,     3,    -1,     1,     3,     0,    -2,    -6,    -1,     0,     0,     0,     2,     0,     3,     1,     0,     1,     0,     0,    -4,    -4,    -2,     0,     2,     1,     0,     0,     3,     4,     1,     0,    -2,    -2,    -3,    -3,     0,    -1,    -1,     1,     4,     4,     5,     0,     1,     0,    -2,     0,    -6,    -5,    -2,     2,     4,     3,     3,     3,     1,    -1,     0,     2,     0,     2,     1,    -3,    -1,     1,     0,     0,     0,     1,     1,    -1,     2,    -1,    -2,    -5,    -8,    -4,     2,     0,    -3,    -1,     1,     1,     0,     0,     0,     2,     2,     0,     2,    -3,    -5,    -1,    -1,     0,     0,     5,     2,    -4,     1,     0,     0,    -3,    -6,    -2,     2,     1,    -3,     1,    -2,     0,     4,     3,     4,     5,     3,     0,    -1,    -5,    -6,    -6,    -3,     1,     0,     3,     3,    -2,    -2,     0,     0,    -4,    -9,     3,     4,     2,     1,    -2,    -1,     2,     3,     6,     4,     4,     4,     0,    -6,    -3,    -4,    -4,    -2,    -8,    -7,     2,     4,     3,    -2,     0,    -1,     0,    -2,     1,     2,     1,    -1,    -1,    -1,     0,     1,     3,     3,     1,     3,     1,    -1,    -2,    -5,    -3,    -2,    -8,    -9,     0,     0,     1,     1,     0,     0,    -1,    -1,     2,     1,     0,     0,     0,     0,     0,    -3,     1,     0,    -1,     1,    -2,    -2,     0,    -1,    -3,    -1,    -6,    -4,    -9,    -4,     3,    -4,     0,     0,    -2,     0,     0,     2,    -1,     0,     0,     0,     0,     1,     0,     0,    -1,     1,    -1,    -3,     0,     1,     0,     0,    -1,    -5,    -7,    -5,     0,    -3,     1,    -1,    -1,     0,    -4,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,    -2,     1,    -2,     2,     0,    -2,     1,     2,    -1,     0,     4,     0,    -4,    -2,    -1,     0,     0,    -2,    -1,     1,     0,     0,    -1,    -4,    -3,     1,     0,     0,    -2,     0,     0,    -1,    -1,     0,    -2,    -2,    -5,     0,     4,     2,    -4,    -3,    -4,     0,    -1,    -4,     4,     0,     1,    -5,    -8,    -4,    -4,    -2,     3,     0,    -1,    -1,    -2,    -1,    -2,     0,     1,    -1,    -2,     0,     2,    -1,    -8,    -4,    -4,     0,    -1,    -7,     7,     1,     0,    -2,    -7,    -5,    -4,    -2,     0,    -3,    -2,    -2,    -1,     1,     2,     1,     3,     0,     0,     1,     1,    -4,    -8,    -6,    -6,    -1,     1,    -4,     7,     6,     4,     0,    -4,    -5,    -8,    -1,    -3,    -2,    -3,     0,     0,     1,     2,    -1,    -1,     1,     2,     2,     3,     0,    -1,    -7,    -2,     0,    -2,     3,     0,     5,     5,     1,    -3,    -1,    -4,    -2,    -2,    -1,     0,     0,     2,    -1,     1,     4,     0,     4,     0,     3,     4,     4,     2,    -4,    -5,    -1,    -2,     3,    -1,     2,     3,     0,     0,     0,    -1,    -3,     0,     0,     2,    -1,    -1,     2,     3,     0,    -2,     2,    -1,     5,     2,     2,     4,    -4,     0,     0,    -1,    -3,    -6,     0,     2,    -1,    -2,     2,     2,     0,    -1,    -1,     0,     1,     3,     3,     1,     3,     3,     1,     3,     0,     3,     1,     5,     2,    -1,    -1,     0,    -5,    -2,    -4,    -3,    -2,     0,     1,     1,     2,    -1,     0,     1,    -1,     0,     1,     0,     1,     2,    -2,     0,     0,     6,     6,     7,     4,     0,     0,     0,     1,     1,    -2,    -1,     0,    -1,    -3,     0,    -1,     0,    -1,     1,     1,    -1,     1,     1,     2,     2,    -1,     1,    -2,     4,     4,     5,     3,     0,     1,     0,    -3,    -1,    -3,    -2,    -2,     1,     2,     4,     3,     3,    -1,    -2,    -3,     1,    -1,     3,     2,     3,     1,    -2,     1,     0,     5,    -3,    -2,     0,     1,     0,     0,     2,    -5,    -6,    -2,    -1,     1,    -2,    -3,    -3,     0,    -2,    -4,     0,     3,     5,     4,     3,     1,     3,     5,     4,     4,    -2,    -1,     0,     1,     0,    -1,    -1,    -2,    -4,    -6,    -5,    -2,     0,     1,     1,     0,    -1,    -5,     2,    -1,     1,     1,     5,     1,     0,    -1,    -2,    -1,     0,     1,     0,     0,     1,     1,     0,    -1,    -1,     0,    -1,    -1,    -1,     1,     1,     1,     0,    -6,    -5,    -1,    -2,    -1,    -3,    -3,    -4,    -2,     0,     0,     0,     0,     0),
		    56 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     1,    -1,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     1,     2,     3,     2,     1,     1,     0,     2,     0,    -1,    -1,     0,     0,     1,     4,     2,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     2,     0,     1,     3,     3,     2,     2,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,     2,     2,     3,     2,     3,     1,     1,     0,     0,     0,    -1,    -3,    -3,    -1,     2,     2,     1,     1,     2,     0,    -2,    -3,    -6,    -3,    -1,     0,    -2,     1,     3,     2,     1,     1,     3,     2,     0,     0,     0,     1,     0,    -3,    -4,     3,     3,     2,     0,    -1,     1,     0,    -3,    -4,    -6,    -4,     0,    -1,    -2,    -4,     0,     0,    -1,    -3,     0,     3,     2,     4,     4,     0,     1,    -2,    -3,     5,     3,     1,     1,     1,     0,     0,    -2,    -2,    -4,    -2,     1,    -1,     1,    -2,    -2,    -2,    -1,    -1,     1,     2,     2,     4,     3,     0,     0,     1,    -1,     4,     1,     2,     1,     4,     2,    -2,    -4,    -4,    -5,    -1,    -1,    -4,    -2,     0,    -3,    -2,     0,    -1,     0,     1,    -2,     1,     5,     0,     0,     0,    -1,     4,     2,    -1,     2,     2,     2,    -1,    -4,    -5,    -3,     0,    -3,    -4,     0,     0,    -1,    -1,    -2,    -2,    -3,    -3,    -1,     2,     4,     0,     0,     0,    -1,     3,     1,    -1,     2,     0,     0,    -3,    -5,    -5,     0,     0,    -4,    -1,     2,     1,     1,     2,     1,    -2,    -1,    -1,    -1,     2,    -3,     0,     0,    -1,    -3,     2,     1,    -1,     2,    -1,    -2,    -5,    -6,    -5,    -2,    -1,    -2,     1,     3,     0,     1,     2,     0,    -1,     0,    -1,    -3,    -1,    -1,     0,     0,    -1,    -3,     3,     2,     1,     4,     0,    -3,    -4,    -5,    -4,    -1,     0,     1,     1,     2,    -2,    -1,    -1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,    -1,     2,     2,     2,     1,     0,    -2,    -3,    -4,    -2,     0,     1,     0,    -1,    -4,    -3,    -1,    -2,     0,     1,     2,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,     1,     4,     0,     1,     0,    -2,    -3,    -4,    -1,     4,     1,     1,     1,    -2,    -2,    -2,    -1,     1,     2,     2,     2,     0,     0,    -3,     1,     1,     0,    -1,     1,     1,    -1,     0,     1,    -2,    -2,    -5,     0,     2,    -1,    -2,     0,     0,    -2,    -2,    -1,     1,     1,     2,     2,     0,     0,    -1,     0,     0,     0,    -2,     0,     1,    -1,     1,     0,     0,    -3,    -2,     2,     3,    -4,    -3,     0,     0,    -1,    -1,    -2,    -1,     0,     1,     1,     0,    -1,    -1,    -1,     0,     0,    -1,     2,     1,    -1,     0,     0,     0,    -2,     0,     0,     1,    -2,    -1,     0,    -1,     0,    -2,    -2,     0,     1,     2,     1,     0,     0,    -4,     0,     0,    -1,     0,     2,     0,    -2,    -1,    -2,    -1,    -1,    -1,     2,     0,     1,     3,     0,     0,     2,    -3,    -1,     0,     2,     1,     0,     1,     0,    -2,     0,     0,     0,     2,     0,     0,    -1,    -1,    -1,     0,     1,     0,    -1,     2,     0,     1,     3,     0,     1,     0,    -2,     0,     0,     1,     0,     0,    -1,    -2,     0,     0,     0,     0,    -1,     1,    -2,    -2,    -2,     0,     0,     1,    -1,     1,    -1,     1,     1,     0,     2,     1,     0,    -1,     1,     2,     0,     0,     0,    -1,    -1,    -1,    -1,     2,     0,     0,    -3,    -3,    -3,     0,     0,     0,    -1,     0,     1,     2,     0,     0,     2,     3,     2,     1,     0,    -2,    -1,     1,    -3,     0,     0,    -1,     0,    -1,    -1,    -2,    -1,    -4,    -3,    -1,     1,    -1,    -1,     1,     1,     2,     1,     3,     2,    -2,     0,    -1,    -4,    -2,    -1,     1,    -1,     0,    -1,     0,     0,    -1,     0,    -2,     0,    -2,    -1,     0,     0,     0,     0,     2,     1,     1,     1,    -1,    -2,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,    -2,     0,    -1,    -2,    -1,     0,     0,    -1,    -2,     0,     2,    -1,     1,    -1,    -1,    -3,     0,     0,    -2,    -3,    -3,    -3,    -1,     0,     1,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,    -2,     0,    -3,    -2,     1,    -2,    -4,    -2,    -1,    -1,     0,    -2,    -2,    -2,     0,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,    -2,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -2,    -1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0),
		    57 => (    0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,    -2,    -5,    -6,    -7,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -4,    -4,    -6,    -5,    -3,    -2,    -1,    -3,    -3,    -1,    -2,     0,    -3,    -3,    -2,    -2,    -2,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -4,    -7,    -7,    -6,    -4,    -6,    -9,    -9,    -6,    -6,    -5,    -4,    -2,    -2,    -4,    -2,    -3,    -9,    -6,    -3,    -1,     0,    -1,     0,     0,     0,    -3,    -3,    -5,    -6,    -9,   -10,   -12,   -12,    -2,    -1,    -1,    -2,    -3,    -7,    -9,    -8,    -5,    -4,    -3,    -6,    -8,    -8,    -4,    -1,     0,     1,     0,     0,    -3,    -5,    -2,    -4,    -3,    -1,     2,    -2,     1,     3,     2,     0,    -1,    -2,    -5,    -6,    -8,    -8,    -5,    -5,   -11,    -8,    -7,    -1,     0,     0,     0,    -2,    -2,    -1,     2,     1,     1,     0,     1,     3,     3,     0,     1,    -3,    -1,     1,    -2,     0,    -3,    -4,    -2,    -4,    -4,    -5,    -5,    -3,    -2,     0,     2,    -2,     1,    -1,     4,     3,     3,     2,     3,     3,     0,     1,     2,     2,     0,     2,     2,     3,     2,    -1,    -1,    -1,    -2,    -4,    -8,    -5,    -3,    -2,     1,     0,     2,     0,     4,     0,     1,     1,    -1,     2,     2,    -3,    -3,    -2,     1,     2,     1,     2,     2,     2,     2,    -1,     0,    -4,    -5,    -5,    -2,     0,     2,     2,     2,     2,     0,    -1,     0,     0,    -1,     0,     2,    -1,    -1,    -3,     0,     1,     3,     3,     1,     0,     2,     1,     2,    -4,    -1,     5,     6,     0,     3,     0,    -1,     1,    -3,     0,    -2,     1,     1,     0,     1,    -2,    -3,     0,     0,     2,     2,     3,     2,     2,    -1,     2,    -1,    -1,     2,     4,     5,     0,     0,     0,    -1,     2,     2,    -2,    -1,     0,     2,     1,    -2,    -1,     2,    -1,     0,     2,     1,     3,     2,    -2,     0,     3,     2,    -1,    -4,     0,     3,     0,     2,     2,     0,     3,     4,     0,    -2,     2,    -1,    -3,    -1,    -1,    -1,    -1,     3,     2,     3,     1,     0,     0,     1,     0,     1,     0,     2,     4,     6,     0,     1,     3,     0,     3,     3,    -1,    -1,     1,     0,     0,     0,    -2,     0,    -2,     1,     0,     0,     0,     0,    -1,    -1,     3,     1,     3,     3,    -1,    -2,     0,     1,     1,     0,     0,     2,    -2,     1,     1,    -1,     0,    -1,     0,    -2,    -1,     0,    -1,     2,     0,     1,    -1,    -1,     1,    -1,    -1,    -6,    -6,    -1,     1,     0,    -1,     0,    -1,    -2,     0,     1,     1,     1,     2,     1,    -1,     0,     1,     2,    -1,     0,     1,     1,     0,     0,    -2,    -4,    -5,    -6,    -1,    -4,     0,     0,    -1,    -3,     1,     2,    -2,    -2,    -1,     1,     1,     0,     1,     3,     2,     5,     1,     1,     0,    -1,    -2,    -1,    -1,    -1,    -2,    -6,    -4,    -4,    -1,    -1,    -2,    -4,     1,     1,     0,    -2,    -2,    -4,    -1,    -2,     2,     3,     2,     2,     0,    -1,    -2,    -2,    -1,    -1,     0,     0,     3,    -3,    -2,    -4,     1,     0,     1,    -7,     0,    -1,    -3,    -2,    -2,    -2,    -2,     0,     1,     1,     1,    -1,    -4,     0,     0,    -2,     3,     3,     1,     3,     1,    -5,     1,    -3,     1,     1,     0,    -3,    -2,     0,    -1,    -3,     0,    -2,    -2,    -1,     1,     2,    -1,    -4,     0,     0,    -1,     0,     1,     3,    -1,    -3,     2,    -5,    -5,    -2,     0,     0,    -1,    -2,    -6,    -4,    -3,    -2,    -4,    -2,    -4,    -4,    -2,     1,     1,    -2,    -1,     0,    -5,     0,     0,     1,    -2,    -5,    -2,    -5,    -4,     0,     0,     0,    -2,    -4,    -5,    -1,    -1,    -1,    -2,    -4,    -1,    -1,    -1,     1,    -1,    -1,     1,     0,    -4,    -2,    -2,     3,    -2,    -5,    -7,    -2,    -1,     0,    -1,    -1,    -3,    -4,     0,     1,     0,    -1,     2,     0,    -1,    -1,     1,    -2,     0,     0,     3,     0,    -1,     1,     3,     0,    -3,   -12,    -6,    -1,    -2,     0,     0,    -1,    -2,    -4,     1,     1,     1,     1,     3,     1,     0,     1,     3,     2,     4,     1,     2,     2,     0,     0,     2,     0,    -3,   -10,    -6,    -3,    -5,     0,     0,     0,     2,    -1,     4,     4,     4,     4,     3,     0,     2,     3,     3,     6,     6,     0,     4,     3,     1,     2,     2,     1,    -1,    -7,    -4,    -4,    -3,     0,     0,     0,     0,     2,     2,     2,     2,     2,     2,     3,     5,     4,     3,     3,     1,    -2,     5,     2,     2,     2,     0,     3,     3,    -1,    -1,    -3,    -2,     0,     0,     0,     0,    -2,    -2,    -3,     0,     2,     2,     3,     4,     4,     3,    -3,    -5,    -1,     2,     0,     1,     3,     2,     3,     4,     1,    -2,     0,     0,     0,     0,     0,     0,     0,     1,     1,    -1,    -1,     0,     2,     3,     1,     0,    -4,    -1,     1,    -2,     2,     1,     1,     1,     3,     1,     4,     0,     0,     0,     0),
		    58 => (    0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,    -2,    -1,    -1,    -1,    -2,    -2,    -2,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -4,    -4,    -5,    -3,     0,     0,    -2,    -2,    -3,     1,     0,    -2,    -2,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -4,    -7,     1,     2,     2,     0,    -2,    -2,    -2,     2,    -2,    -3,     1,    -2,    -1,    -2,     2,     3,     0,    -1,    -2,     1,     0,    -2,    -2,    -5,    -4,    -4,    -2,     3,     6,     5,     4,     2,    -1,     0,     2,     2,     2,     4,    -1,    -2,    -3,    -4,    -2,    -3,    -4,     0,     2,    -1,     0,     0,    -3,    -4,    -3,    -5,     0,     6,     2,     3,     2,     3,     4,     2,     0,     1,     2,     4,     0,     4,     0,     1,     1,    -1,    -2,    -1,    -3,    -1,     0,    -1,    -5,    -4,    -4,    -2,    -2,     3,    -1,     0,     2,     0,     0,     1,     0,     1,     0,    -1,     1,     1,     2,     0,     0,     2,    -1,    -2,    -1,    -1,     0,    -3,    -4,    -5,    -4,    -3,     0,     0,    -1,     0,    -1,     3,     0,     1,    -2,     2,     1,     0,    -1,     1,    -1,    -1,    -1,     5,     3,    -5,    -3,     1,     1,    -2,    -4,     0,     0,     0,    -1,     3,     1,     1,     1,     0,    -1,     1,     0,     0,    -1,     0,     2,     4,    -2,     3,     3,     4,     5,    -3,     4,     4,     0,    -1,    -5,     1,     2,    -1,     0,     2,     1,     0,    -2,     0,     0,     0,     1,    -1,    -1,     1,     1,     0,     3,     3,     3,     2,     1,    -1,     4,    -5,     0,     0,    -6,    -4,     5,     2,    -2,     2,     2,     1,     2,     1,     1,    -1,     2,    -4,    -3,     0,    -1,     0,     1,     3,     1,     3,     2,    -4,     2,    -2,     0,    -1,    -3,     0,     5,     4,     1,     3,     1,     0,     1,     0,    -1,    -1,     1,    -4,    -3,    -2,     0,     0,     1,     2,     2,     3,     3,     1,     5,    -1,     0,     0,    -4,     1,     5,     8,     0,     0,     3,     1,     0,    -2,    -3,    -2,     0,    -2,     0,     0,    -2,    -1,     2,     2,     4,     0,     2,    -2,     2,    -4,     1,     0,    -2,     0,     2,     5,     2,     1,     2,     0,     0,    -1,    -1,    -1,    -1,     1,     0,    -3,    -2,    -1,     2,     1,     4,     0,    -2,    -3,     2,     1,     0,    -1,    -1,    -3,    -4,     1,     3,    -4,     2,    -5,    -3,    -1,    -2,    -2,     0,     0,    -1,    -3,     0,    -3,    -4,     1,     0,    -1,    -3,    -1,    -2,    -1,     0,     0,    -2,     2,    -7,    -2,    -2,    -3,     1,    -3,    -1,    -1,    -4,     0,     1,    -2,    -2,     0,    -3,    -1,    -2,    -3,    -1,    -4,    -5,    -1,    -6,    -3,     0,    -1,    -1,     2,    -7,    -3,    -4,    -6,    -3,     0,    -4,    -3,     0,     2,     0,    -1,    -3,    -5,    -2,     0,    -3,    -4,    -2,    -1,    -2,    -2,    -6,    -3,     0,    -1,    -1,    -3,    -2,    -4,    -4,    -4,    -1,    -2,    -2,    -4,    -1,    -1,    -2,    -4,    -2,    -2,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -6,    -3,    -5,    -1,    -1,    -2,    -6,     0,    -4,     0,     1,     1,    -1,    -1,    -2,     1,     0,    -2,    -7,     0,     1,     0,     1,    -1,    -1,     0,     0,     0,    -6,    -2,    -3,     0,     0,    -5,    -6,    -1,    -4,    -2,     1,     4,     1,     1,    -1,    -2,    -2,    -4,    -3,    -1,     3,     0,     1,     1,    -2,     1,     3,     4,    -8,    -6,    -4,     0,     0,    -2,    -5,    -4,     1,     2,     0,     3,    -1,     3,     0,     2,     0,    -3,    -1,     3,     2,     0,     0,     2,     3,     2,     6,     1,    -9,    -6,     0,    -2,    -2,    -2,    -3,    -3,     1,     4,     1,     3,     4,     2,     2,     1,     2,     2,     5,     0,     3,    -4,     2,     0,     0,     5,     4,    -2,    -7,    -4,     0,    -2,    -2,    -1,    -2,     2,     4,     2,     4,     3,     3,     5,     5,     2,     3,     6,     6,     1,     1,     1,    -1,     0,     0,     4,     2,    -2,     0,    -4,     0,    -1,     0,    -1,    -1,     4,     0,     2,    -1,     2,     2,     0,     1,     4,     4,     4,     4,     4,     3,     4,     5,     1,    -1,     5,     3,    -1,     0,    -4,     0,     0,     0,    -2,    -3,    -2,    -2,    -1,    -1,     1,     3,     1,     0,     3,     1,     2,     3,     5,    -1,     0,    -1,     1,    -3,     1,     1,    -3,    -6,    -3,     0,     1,     0,    -2,     0,    -7,    -6,     0,     0,    -2,    -4,    -2,    -2,    -2,    -1,     2,     2,    -1,    -1,     1,    -1,    -4,    -4,    -4,    -2,    -2,    -2,    -1,     0,     0,     0,     0,    -2,    -3,    -6,    -5,    -1,     1,     0,    -3,    -2,     1,     1,    -5,   -10,    -5,    -3,    -2,    -7,    -6,    -3,    -3,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,    -2,     0,    -1,    -2,    -4,    -5,    -4,    -2,    -3,    -2,    -2,     0,     0,    -1,     0,     0,    -1,     0,     0),
		    59 => (    0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     1,     0,    -1,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     1,    -1,     0,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,    -2,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -2,    -2,    -1,    -2,    -1,    -3,    -2,    -2,     0,     0,     1,     0,    -2,    -2,    -1,    -1,     0,    -1,     0,     1,     1,     0,     0,     0,     0,    -1,    -3,    -1,    -1,     0,    -1,     0,    -4,    -5,    -4,    -3,    -3,    -3,    -1,    -3,    -4,     0,    -1,     0,     0,    -3,    -2,    -1,    -1,     0,     0,     0,    -1,     0,    -1,    -2,    -5,    -2,    -2,     0,     1,     0,     1,     0,    -1,    -4,    -5,    -3,    -1,    -1,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,    -2,    -3,    -2,    -4,    -1,     2,     0,     3,     3,     2,     0,    -1,     2,    -1,    -6,    -6,    -3,     0,     0,     0,     0,     0,     0,    -2,    -1,     0,    -1,     0,    -1,    -3,    -5,    -4,     0,    -2,     1,     3,     0,     1,    -1,    -4,    -3,    -3,    -7,    -9,    -3,     1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,     2,     0,    -3,     3,    -1,     2,     0,     0,     1,    -1,     0,    -1,    -3,    -3,    -2,     1,    -2,    -5,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -2,     1,     0,    -2,     2,     2,     1,     2,     3,    -1,    -2,     1,     0,    -3,    -4,     2,     2,    -2,    -3,    -2,    -3,    -1,    -2,    -3,    -1,    -1,     0,    -1,    -1,     1,    -1,    -3,     3,     1,     1,     0,     0,    -5,    -5,     1,     3,    -1,     2,     0,     0,    -2,    -3,    -3,    -3,    -2,    -2,    -2,     0,    -2,     0,    -3,    -1,     2,    -1,    -4,     1,     3,     2,     1,    -1,    -1,     2,     6,     0,    -1,    -1,     2,    -1,     0,    -5,    -5,    -3,    -3,    -1,    -2,     0,    -2,     0,    -1,    -1,     2,    -1,     1,     1,    -1,     0,     2,     1,     0,     2,     4,    -2,    -3,    -1,     2,     0,     0,    -2,    -3,    -4,    -3,    -2,    -2,    -2,    -2,     0,    -1,    -1,    -2,    -2,     0,     5,     1,    -3,     0,     1,    -1,     0,    -1,    -1,    -1,     0,     0,    -2,     1,    -2,    -3,    -3,    -2,    -1,    -1,    -2,     0,    -1,     0,    -1,    -1,    -2,    -1,     4,     0,    -1,    -1,     3,     0,    -2,    -1,     1,     1,    -1,     0,     0,     0,    -2,    -3,    -4,    -4,    -2,    -3,     0,     0,    -1,     0,    -1,    -1,     2,    -2,    -2,     0,    -1,    -2,     1,     1,    -1,    -4,    -2,     1,     1,     0,    -1,    -1,    -6,    -5,    -3,    -3,    -1,    -1,     0,    -2,     0,     0,    -2,     0,     0,    -1,    -5,    -1,     1,    -2,     1,     6,     2,     1,     0,    -3,    -2,    -2,    -1,    -2,    -7,    -3,    -2,    -1,    -1,    -1,     0,    -3,     0,     0,    -2,     0,     0,    -2,    -4,    -5,     0,    -4,    -1,     2,     3,     2,     0,     0,    -3,    -3,    -2,    -2,    -5,    -3,    -1,    -2,    -3,     2,    -2,    -1,    -1,     0,    -2,     0,     0,     0,    -1,    -3,    -4,    -4,    -4,    -2,     2,    -1,    -1,    -1,    -1,     0,    -3,    -1,    -2,    -3,     0,    -1,    -3,     0,    -2,    -1,    -1,     0,    -2,     0,     0,    -1,    -1,     0,    -1,    -1,    -3,    -5,    -5,    -5,    -3,     2,     1,     0,    -2,    -2,    -3,    -4,    -2,     0,    -2,     2,    -2,    -1,     0,    -1,     0,    -1,     0,     0,     0,    -2,     0,    -2,    -3,    -5,    -6,    -4,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -2,     0,     1,    -2,     0,     0,    -1,     0,    -1,     0,     2,    -1,    -1,     0,     0,     1,    -1,    -2,    -1,     1,    -2,     0,     0,     0,    -3,    -1,    -2,    -1,    -1,     1,     2,    -3,    -1,     0,     0,    -1,     2,     0,     1,     1,     1,     1,     2,    -1,     1,     2,     1,     1,     1,     0,     1,    -1,    -3,    -2,    -3,    -1,     0,     1,    -1,     0,     0,     0,     0,    -1,     1,    -1,    -1,     1,     0,     1,    -1,     1,    -1,     0,     0,     0,     2,     0,     1,     2,    -1,    -1,    -2,     0,     1,     1,     1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,    -1,     2,    -2,    -4,    -3,    -1,     1,     2,     1,     1,     2,     1,     0,     0,     1,     1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,     1,    -2,    -3,    -2,     1,    -3,    -2,     1,     2,     1,    -3,    -3,    -3,    -2,    -1,    -1,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     2,    -1,    -3,     2,     0,     3,     1,     1,     6,     2,    -3,     1,     0,    -1,     1,     1,     0,     0,    -1,    -1,     0,     0,     0,     0,    -1,     1,     1,     1,    -2,    -1,     1,     0,    -2,    -2,     5,     4,     0,    -1,     2,     1,    -2,    -1,     0,     0,     0,     1,     0),
		    60 => (    0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,    -2,    -3,    -1,     0,     1,    -4,     3,     4,     4,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     4,     4,    -1,    -2,     1,    -1,    -2,    -4,    -3,    -4,    -8,    -4,    -2,     0,    -3,    -2,    -2,    -2,    -2,    -6,    -2,    -3,    -1,     0,     1,     0,     0,     0,     4,     1,    -4,    -4,    -4,    -4,    -3,    -2,    -5,    -6,    -3,    -4,    -4,     1,     2,     0,    -3,    -3,    -4,    -6,    -3,    -2,    -3,    -5,     1,     0,     0,     0,    -1,    -1,    -8,    -3,    -3,     0,     3,     0,     1,    -4,     0,    -1,     1,     3,     2,     0,     0,    -3,    -3,    -1,    -2,    -5,    -9,    -4,     0,     0,    -1,    -2,    -1,    -2,    -4,     2,    -1,     1,     5,     3,     3,     1,     0,     2,     2,     2,     2,     2,     0,     0,    -1,    -2,    -2,    -5,    -8,    -2,    -1,     0,     0,    -3,     0,    -5,     1,     3,     3,     3,     2,     3,     2,     0,     0,     2,    -2,     1,    -1,    -2,     1,    -1,    -3,     0,    -6,    -3,    -9,    -3,    -1,     0,    -1,    -2,    -3,    -3,     0,     3,     3,    -1,     1,    -1,     1,     1,     1,    -3,    -3,    -1,    -1,    -1,    -3,    -1,    -3,    -1,     0,    -3,    -2,    -5,     1,     6,    -4,     0,    -4,    -4,     0,     0,    -3,     1,     1,    -1,    -3,     0,    -1,    -5,     0,    -1,     2,     0,    -1,    -2,     1,     0,     2,    -4,    -8,    -4,    -1,    -1,    -1,     2,     0,    -1,     1,    -3,    -1,    -1,     1,    -1,     1,     2,     1,     1,     2,     2,     2,     1,     1,     1,    -1,     0,     2,    -1,    -5,    -1,    -1,    -1,    -1,     3,     1,     0,    -2,    -1,    -2,     0,     2,    -1,    -1,     0,     2,     6,     4,     4,     5,    -1,     2,     1,    -2,     1,     2,     0,    -3,    -4,     0,     0,     6,    -4,     0,    -1,    -4,    -1,    -2,    -2,    -1,    -2,     0,     2,     7,     3,     3,     8,     6,     5,     3,     2,     1,     1,     1,     4,    -4,    -4,     0,     0,     0,    -4,    -1,     2,    -4,    -3,    -4,    -3,    -1,    -1,     0,     4,     5,     4,     4,     3,     3,     3,     2,    -1,     0,     0,     1,     2,    -2,    -3,    -2,     0,     1,     0,    -2,     3,    -1,     0,    -2,    -1,    -2,    -2,     1,     1,     0,     0,     1,     0,    -1,    -1,    -1,    -1,     1,     1,     3,     1,     2,    -5,    -2,     0,     0,    -1,    -5,    -2,    -1,    -2,    -1,     0,    -1,    -2,     0,    -1,    -1,    -5,    -5,    -6,    -2,     1,    -1,     2,     4,     5,     3,     4,     4,    -5,    -1,     0,     0,    -3,    -4,    -1,    -2,    -3,     1,     0,    -3,    -3,    -2,    -3,    -3,    -7,    -4,    -3,    -1,    -2,     0,     3,     2,     0,     2,     3,     4,    -5,    -4,    -1,     0,    -2,    -2,     2,    -1,    -3,     1,    -1,    -2,     0,    -2,    -3,    -4,    -4,    -1,    -3,    -3,    -1,     2,     2,    -1,    -2,    -3,     0,    -1,    -7,    -2,     0,     0,    -2,     0,     1,     1,    -2,     1,    -1,     1,     1,     2,     1,     3,    -2,    -2,    -3,    -1,    -1,     2,     0,    -4,    -1,    -1,    -1,    -4,    -4,     1,     0,     0,    -2,    -1,     2,     2,     2,    -1,     1,     2,     3,     1,     0,    -2,    -3,    -1,    -1,     1,     1,     1,    -3,    -2,    -1,     2,    -4,    -4,    -3,    -2,     0,     1,    -1,    -1,     0,     3,     2,     4,     3,     1,     0,     1,     3,    -1,    -2,     0,     0,     0,     0,     3,    -1,    -2,    -1,     2,     0,    -7,    -1,    -1,     0,     1,    -3,    -2,     4,     2,     2,     3,     2,     4,     0,     1,     4,     1,     0,     2,     0,     1,     0,     1,    -3,    -3,    -2,    -1,    -2,    -8,     1,     0,     0,    -1,    -3,    -2,     0,     0,     3,     4,     4,     3,     2,     1,     2,     0,    -1,     2,     1,     0,     1,     1,    -1,    -2,     0,     0,    -4,    -4,     8,     0,     0,     0,    -2,    -2,    -5,    -3,    -1,     4,     3,     1,     4,     2,    -1,    -1,     1,     3,     2,     1,    -1,    -1,    -3,    -3,    -1,     0,    -3,    -2,     5,     1,     0,     0,    -2,    -4,    -1,    -3,    -3,     0,     3,     2,     2,    -2,     2,    -1,     1,     1,     1,     3,    -1,    -3,    -5,    -4,    -4,    -1,    -3,    -4,    -4,    -1,     1,     0,    -1,    -2,     1,     2,    -3,    -2,    -2,    -1,    -2,    -6,    -4,    -3,    -3,     2,    -1,     0,    -2,    -5,    -3,    -5,    -4,    -3,    -3,    -1,     0,     0,     0,     0,    -1,    -1,    -5,    -3,    -5,    -8,    -5,    -5,    -5,    -3,    -5,    -3,    -3,    -4,    -9,    -8,    -8,    -9,    -6,    -7,    -5,    -2,     0,     0,     1,     1,     0,     0,     0,     0,    -2,    -5,    -7,    -3,    -3,    -5,    -3,    -4,    -3,    -3,    -4,    -6,    -5,    -5,    -5,    -6,    -5,    -6,    -4,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,     0,     0,     0,    -4,    -1,    -1,     0,     0,    -2,    -2,    -1,    -3,    -1,    -2,     0,     0,    -1,     1),
		    61 => (    0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -2,    -5,    -5,    -2,    -1,     0,     1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,     5,     3,     1,    -1,     0,     2,     1,     1,    -1,     0,    -4,   -10,    -8,    -6,    -4,    -4,    -2,     0,     0,    -1,     6,     1,     0,    -2,     0,     1,     1,    -1,     4,     4,     2,    -1,    -2,    -1,    -4,    -2,    -3,    -4,    -6,    -7,     3,     2,     2,     2,     1,     1,     0,     1,     2,    -2,    -3,    -4,    -3,    -3,     0,    -1,     3,     5,     3,     1,    -1,    -2,    -7,    -5,    -7,    -7,    -7,    -4,     0,     2,    -1,    -2,    -4,    -2,    -1,     1,     3,     0,    -2,    -4,    -4,    -3,     0,     0,    -3,     2,     4,    -2,     3,     5,    -3,    -7,    -8,    -7,    -4,    -1,     0,    -1,    -1,     0,    -2,    -1,     2,     0,     0,    -1,    -3,    -3,    -2,    -2,    -1,    -4,    -4,    -1,    -3,     3,     3,     4,    -5,    -5,   -11,    -6,    -3,    -2,     0,     0,     2,     1,     0,     2,     3,     0,    -2,    -1,    -4,    -3,    -2,    -2,     0,    -3,    -4,     1,    -3,     2,     3,     1,    -3,    -4,    -5,    -6,    -6,    -3,     0,     2,     2,     1,     1,     1,     1,     0,    -2,    -3,    -5,    -2,    -4,    -1,     0,     0,    -3,     1,    -2,    -2,     3,     4,     2,     1,    -1,    -6,    -2,    -5,     0,     3,     5,     1,     2,     0,    -1,    -2,    -2,    -1,    -3,    -1,     0,    -1,     0,     1,    -4,    -1,    -2,    -3,     0,     3,    -1,    -1,     2,    -1,    -2,    -4,     0,     1,     2,     1,    -1,    -2,    -5,    -6,     0,    -1,    -3,     0,     0,     4,     0,     0,    -1,     2,     0,     3,     2,    -4,    -6,    -2,     1,    -1,    -6,     0,     1,     1,     1,     0,    -2,    -5,    -2,    -1,     0,    -1,    -1,     0,     0,     3,     0,     0,    -2,     3,    -1,     4,     3,    -1,    -2,     0,    -1,    -2,    -2,     1,     2,     1,     1,     2,    -3,    -4,    -1,     3,    -1,    -2,    -3,     2,     0,     3,     0,     0,    -1,     2,     1,     1,     3,     1,     2,     2,    -1,    -3,    -2,     0,     3,     0,     1,     3,    -5,    -8,    -4,     3,    -2,    -2,    -3,     0,     0,     1,     0,     0,     2,     1,     4,    -2,    -2,    -6,     2,     0,     1,    -2,    -2,     1,     1,    -1,     2,    -1,     0,    -4,    -3,     4,     2,     0,    -1,     3,     4,     0,     0,     0,     0,     4,     2,    -5,     0,    -1,     2,     0,    -1,     1,     0,     1,    -2,    -2,     3,     2,    -6,    -6,    -2,     1,     0,    -2,    -3,     2,     2,    -1,     0,     1,     2,    -1,     0,     0,     0,    -4,     0,     0,    -4,     1,    -2,     2,    -1,    -1,     3,     0,    -3,    -6,    -3,     2,     0,     2,     2,     1,     0,    -1,    -1,     0,     0,    -4,     1,     0,     1,    -1,    -2,    -2,    -3,     2,     0,     1,    -1,    -2,    -1,    -5,    -4,    -3,    -2,     1,    -1,     0,     1,     2,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -5,    -4,    -4,    -1,     0,    -1,     1,     0,     1,    -1,    -2,    -4,    -4,    -3,    -4,    -4,     1,     0,     2,     1,     2,     0,     2,    -1,     0,     2,     1,     0,    -4,    -1,    -2,    -1,     2,     0,     1,    -1,     2,     0,     0,    -3,    -2,    -1,    -4,    -3,     0,    -2,     2,     3,     3,     1,     2,     0,     0,     2,     0,     2,    -1,    -1,    -2,     0,    -2,     0,     0,    -1,     1,     2,    -1,     0,    -4,     0,    -1,     2,    -1,    -1,     1,     4,     4,     0,     0,     2,     3,     2,     2,     1,     3,    -2,     0,     0,    -1,     1,    -2,     0,     0,     0,     0,    -2,    -5,     0,     2,     4,     1,     0,     2,     4,     2,     0,     0,     2,     3,     2,     2,    -1,     1,     0,    -3,    -3,    -1,    -2,    -2,     0,     0,     2,     4,     2,     0,     4,     2,     0,    -1,     1,     3,     0,    -1,     1,     0,     1,     1,     0,     0,    -1,    -1,     2,     3,     4,     5,     0,    -1,    -1,     1,     1,     5,     2,     3,     2,     0,    -4,    -4,    -1,    -1,     1,     3,     5,    -1,     0,     0,     0,    -1,    -5,    -4,    -4,    -1,     0,     4,    -2,    -1,    -1,     0,     0,     3,    -1,     0,    -1,     1,     0,     2,     0,    -2,    -1,     2,     1,     0,     0,     0,     1,    -1,    -2,    -2,    -2,    -6,     0,     3,    -8,    -7,     0,    -1,     2,    -1,    -4,    -7,    -4,    -2,    -3,    -2,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -5,    -6,    -5,    -6,    -2,    -3,    -5,    -5,    -3,    -1,     2,    -3,     0,    -1,    -1,    -1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -3,    -2,     0,     0,    -2,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1),
		    62 => (    0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     1,     0,     0,     0,     0,    -2,     2,     1,     0,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,     1,    -1,     1,     5,     3,     6,     2,    -1,    -1,    -2,    -3,    -8,    -6,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -2,    -2,     1,     3,     0,    -1,     2,    -1,     1,    -1,     0,     0,     1,     3,     0,    -4,    -3,    -4,    -2,     2,     0,     0,     0,     0,     0,     1,     0,    -1,     1,     1,     2,     5,     5,    -1,     0,     3,     3,     2,     5,     3,     3,     0,     1,     0,    -2,     1,     1,     1,    -3,    -4,    -1,    -2,    -1,     0,     0,     1,     0,    -1,    -2,    -2,     3,    -1,    -2,     1,     0,     2,     1,     0,     2,     2,     0,     0,    -1,    -3,     2,     4,     1,    -2,    -2,    -2,    -1,     0,     0,     2,     1,    -1,    -4,     1,     1,    -1,     0,    -1,    -1,     0,    -1,     2,     0,     0,    -2,     1,    -3,     0,     2,     5,     1,    -2,    -3,    -1,    -1,     0,     0,     0,     3,     0,    -1,    -4,     0,     2,    -1,     1,     0,     1,     1,     3,     2,     0,    -1,    -2,    -3,     1,     0,     2,    -4,    -3,    -4,    -1,    -1,    -2,     1,     1,     0,     3,    -2,    -3,    -1,     1,     0,     2,     2,    -1,    -2,    -2,     1,     1,     0,    -1,     0,     0,     0,     1,     0,    -2,    -2,    -3,    -1,     0,    -1,     5,    -1,     2,     3,    -3,     0,     0,     0,     0,    -2,     0,    -6,    -9,    -1,     1,     1,     0,    -1,     0,     0,     0,     2,    -4,    -2,     1,    -1,     0,    -1,     3,     1,    -1,     0,    -1,     3,     1,    -2,    -2,    -2,    -5,    -7,    -3,    -3,     0,     0,    -2,     0,    -2,     1,    -4,     2,    -2,    -1,     2,    -1,     0,     0,    -1,     2,     2,    -1,     0,    -1,    -1,    -5,    -4,    -7,    -8,    -8,    -2,    -1,     0,    -2,    -3,    -2,    -1,    -1,    -2,     3,     0,     0,    -2,     0,     0,     0,    -2,    -1,     0,    -1,    -2,    -7,    -5,    -6,    -6,    -5,    -6,    -2,     0,    -2,     2,     0,    -3,    -2,     0,     0,    -2,     2,     0,     1,     3,    -1,     0,     0,     2,     0,    -1,    -4,    -6,    -9,   -10,    -9,    -5,    -4,    -2,     3,    -1,    -2,     1,     0,    -1,    -4,    -3,    -1,    -3,     1,    -1,     0,     3,     0,     0,    -1,    -1,     0,     0,    -4,    -5,    -7,    -7,    -5,    -1,    -1,     0,     1,    -2,    -2,     0,    -1,    -3,    -2,    -3,    -1,     0,    -1,    -1,     0,     2,     2,     0,    -1,     0,    -1,    -4,    -3,    -1,    -3,    -1,     2,     3,     2,    -1,     1,    -1,    -2,     0,    -2,    -3,    -2,    -4,     0,     0,    -1,    -1,     2,     2,     4,    -1,     0,     0,    -2,    -4,    -2,     0,    -3,    -2,     1,     1,     1,     0,     0,     1,    -4,    -1,    -3,    -5,    -3,    -4,    -1,     0,     0,    -1,     5,     2,     2,     0,     0,     0,     0,    -3,    -1,    -3,    -2,    -1,     0,     0,     1,     2,     1,    -1,    -1,    -2,    -4,    -6,    -3,     0,     0,    -3,    -3,    -2,     2,    -1,     2,     1,     0,    -1,     1,     3,    -1,    -1,    -1,     3,     2,     1,     1,     4,    -1,    -1,    -5,    -4,    -3,    -1,    -1,     0,     1,     0,    -2,    -2,     6,    -2,     4,     0,     0,     1,     3,     3,     0,     0,     2,     4,    -1,     2,     2,     4,     2,    -3,    -2,    -3,    -4,    -1,     0,     0,     0,    -3,    -4,     2,     2,     3,     4,     0,     0,     3,     3,     3,     3,    -3,     1,     0,     0,     1,     2,     3,     1,     0,     2,     0,     3,    -3,     1,     1,     1,     0,    -1,     2,     2,     3,     1,     0,     1,     4,     3,     2,     2,    -2,    -1,    -1,     1,     1,     0,     2,    -1,     0,     1,     2,    -2,     0,     3,     1,     2,     2,     2,     6,     7,     2,     0,     0,     0,     3,     3,     1,     0,    -1,     0,     1,    -1,     2,     1,     1,     0,     2,     2,     0,    -5,    -1,     2,     2,    -1,     1,    -2,     0,     1,    -3,    -1,     0,     0,    -1,     1,    -2,     1,     0,     1,     3,     0,    -1,     2,     0,    -1,     1,     3,     1,    -3,     2,     1,     0,     2,     2,     3,     2,     1,    -2,     0,     0,     0,    -2,    -1,    -2,    -4,    -6,    -9,    -6,    -2,     0,     1,     1,     1,     5,     0,    -2,     1,     3,     3,    -2,     2,     7,     4,     4,     1,     2,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -3,    -6,    -6,    -1,     0,    -1,     0,     3,     4,     2,     5,    -1,    -5,     0,     1,     1,     0,     2,     2,     2,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,    -2,    -1,     0,    -2,     0,    -3,    -3,    -2,    -6,    -4,    -3,    -1,     0,     0,    -2,     0,    -1,     0,     0,     0,     1,     1,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,     0,     0,     0,     0,     0,     1),
		    63 => (    0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -1,    -3,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -5,    -4,     2,     2,    -2,    -3,    -4,     0,    -2,    -1,    -1,    -1,    -3,    -2,    -2,    -2,    -1,     0,     0,     1,     1,     1,     0,    -1,     0,     1,     1,     3,     3,     0,    -1,     2,     2,     2,     4,     1,    -2,    -1,    -2,    -2,     1,     0,    -5,    -8,    -4,    -3,     0,     0,     0,    -1,    -2,     2,    -4,     0,     4,     2,     1,    -2,    -1,    -1,     1,     2,     3,     0,     0,    -4,    -3,    -1,    -2,     1,     1,   -10,    -9,    -5,    -4,     1,     0,     0,    -1,     0,    -2,    -1,     2,     0,    -2,    -3,    -1,     2,     3,     0,     1,    -1,     1,     1,     0,     1,     1,     5,     2,     3,     2,    -8,    -2,     0,     0,     0,     2,     1,     2,    -1,     1,     3,    -4,     0,     1,     3,     1,     1,    -2,    -2,    -1,     1,     1,     0,     4,     4,     0,    -1,     2,    -6,    -4,    -1,     0,     1,     0,     2,     6,     2,     4,     1,     0,     0,     1,     3,     2,     0,     2,     2,    -3,    -1,     0,     3,     0,     1,    -3,    -1,     1,    -5,    -7,    -2,    -1,     0,     0,     1,     2,     1,    -1,    -2,     1,     0,     0,     1,     0,    -2,     2,     1,     1,    -2,     2,     4,     2,     3,    -2,    -1,    -1,    -7,    -7,    -1,     0,    -2,    -1,    -1,     2,     1,     0,    -1,     0,    -1,    -2,     0,     0,     1,     2,     1,     3,     2,     1,     1,    -1,    -2,    -1,    -2,    -8,    -9,    -8,    -3,     0,    -3,    -2,    -2,    -1,    -2,    -3,     0,    -1,     0,    -1,     0,     2,     2,    -2,     0,     1,     4,     1,    -4,    -1,    -6,    -3,    -1,    -6,    -4,    -6,    -3,     0,    -3,    -3,     0,    -1,    -1,    -1,     1,     0,    -2,     0,     1,     0,    -1,    -2,    -2,     0,     6,     2,     0,    -1,    -3,    -3,    -3,    -8,   -10,    -6,    -1,     0,    -2,    -4,     0,    -1,     0,    -1,    -2,    -1,     0,     0,     1,     3,     0,    -1,    -1,     2,     3,     3,     3,     2,    -1,    -1,    -1,   -10,    -5,    -3,     0,     0,    -1,    -3,     0,    -3,    -2,    -2,     0,     0,    -3,    -1,     0,     2,    -1,    -1,    -2,     4,     3,     1,     3,     2,     1,    -2,    -1,    -1,    -6,    -5,    -2,    -1,     1,     0,    -1,    -3,     0,     0,     0,    -1,    -2,     0,     1,     1,    -1,    -2,    -1,     1,     4,     3,     5,     2,     3,    -1,     0,     2,    -7,    -4,    -1,     0,     1,     0,     0,    -1,     4,     4,     0,     0,    -1,    -2,     0,    -2,     0,    -2,    -1,     1,     2,     1,     3,     2,     1,     1,     1,     3,    -4,    -2,    -1,     0,     1,     0,     1,     0,     1,     4,     2,    -1,     0,     0,     0,     1,    -2,    -2,    -2,     2,     4,     2,     1,     3,     3,    -1,    -2,     0,    -6,    -7,    -2,     0,     0,     0,     3,    -1,    -1,     4,     4,    -2,    -1,     0,     0,     1,    -1,    -4,     0,     3,     2,    -1,    -2,     0,     0,    -1,    -1,    -7,    -6,    -3,    -1,    -2,     1,     1,     3,     0,    -1,     3,     1,     0,     1,     2,     1,     0,    -4,    -1,     2,     2,     0,    -2,     0,     1,     1,    -1,    -3,    -6,    -6,    -1,    -2,     0,    -3,    -1,     0,     3,     3,     2,     3,     1,     1,     2,     0,    -4,    -5,    -2,     0,    -4,    -4,    -1,    -1,     0,    -2,     2,     0,    -4,    -6,    -6,    -3,     0,    -1,    -2,    -1,     1,     4,     2,     3,    -1,     1,     1,     2,    -4,    -4,    -2,    -2,    -4,    -5,    -3,    -1,    -2,    -4,     3,     0,    -1,    -4,    -1,    -1,     0,     0,     1,     0,    -1,     1,     2,     0,    -1,     0,     2,     4,     1,    -3,     0,     0,     0,    -2,     0,     1,    -1,     0,     1,     0,    -3,    -5,    -2,     0,    -1,    -1,     2,     0,    -1,     1,     2,    -1,     1,    -1,     4,     5,     3,    -3,    -1,     3,     0,     1,     2,    -1,     0,     0,     3,    -1,    -6,    -4,    -3,     0,     0,     1,     1,     1,     0,     0,    -1,     1,     1,     2,     4,     5,     1,     3,     2,     3,     2,     1,     2,     0,    -1,     1,    -1,    -2,    -3,    -4,    -5,     0,     0,     0,    -1,     3,     0,    -1,     0,     3,     4,     4,     4,     0,     1,     1,     2,     2,     4,     1,    -1,    -2,     0,     1,    -1,     0,    -5,    -4,    -2,    -1,     0,     0,     0,    -2,    -2,     3,     3,     3,     3,     4,     2,    -1,     1,     0,     2,     2,     3,     3,     2,     2,     3,     0,    -3,    -8,    -5,    -2,    -1,     0,    -1,     1,     0,    -2,    -4,     3,     2,     2,    -3,    -3,     1,     1,    -1,    -3,    -3,    -2,     1,     1,    -1,    -1,    -1,    -3,    -3,    -2,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -3,    -3,    -1,    -3,    -3,    -2,     0,    -1,    -2,    -2,    -2,    -1,    -1,     0,     0,     0,     0,     0),
		    64 => (    0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -2,    -2,    -1,    -2,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -3,    -2,    -3,    -5,    -4,    -5,    -3,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -4,    -6,    -3,     0,    -1,    -4,    -3,     0,     0,    -1,     3,     1,    -2,    -1,    -2,     0,     1,     0,     1,     0,     0,     0,    -1,    -1,    -2,     0,     0,    -1,    -1,    -2,     0,    -1,    -2,    -2,    -2,    -2,    -1,    -2,     0,     1,    -2,    -1,     1,     4,     2,     1,    -2,    -1,     0,     1,     0,    -1,    -1,    -2,    -1,    -2,     1,     0,     2,    -4,    -7,    -9,    -7,    -2,     3,     2,    -4,    -4,    -2,    -3,    -1,     3,     0,     2,    -2,    -1,     1,     0,    -1,    -3,    -2,    -1,     2,     1,     1,     3,    -3,    -7,    -8,   -12,    -8,    -1,     1,     3,    -1,    -5,    -2,     0,     2,     3,    -1,    -3,     1,    -2,    -1,    -3,     0,    -2,    -2,     0,     0,     0,     3,     4,     1,    -4,   -10,   -13,    -4,     2,     2,     2,    -5,    -1,     1,     3,     7,     2,    -4,    -4,    -1,    -4,    -2,    -2,    -1,    -3,    -3,    -1,     1,     0,     1,     4,     2,    -3,   -12,    -9,    -2,     1,     3,     0,    -4,    -3,     1,     2,     1,     2,    -5,    -1,    -3,    -3,     0,    -1,     0,    -3,    -2,    -1,    -2,     2,     3,     3,     2,    -1,    -4,    -3,    -1,     0,     1,    -1,    -1,     0,     0,     0,     0,     3,    -2,    -1,    -2,    -1,     0,     1,     0,    -4,     0,     0,    -1,     1,     2,     4,     3,     0,    -4,    -5,    -1,     2,     1,     0,     0,    -1,    -2,    -2,    -2,     0,     2,     1,    -1,    -2,     0,    -1,    -1,    -2,     1,     1,     1,     0,     3,     4,     2,    -2,    -4,    -4,    -3,    -1,    -1,     0,    -2,    -1,     0,    -1,     0,    -1,    -1,     2,    -1,    -4,     1,    -1,     1,    -5,    -2,     0,     2,    -1,     1,     3,     1,     0,     0,     1,    -1,     1,     0,     0,     0,     1,     2,     0,     0,    -4,    -3,    -1,    -2,    -3,     0,     0,    -1,    -3,    -3,    -2,     2,     1,    -1,     3,     1,     0,     0,     2,     1,     2,     0,     1,     2,     4,    -1,     1,     1,    -5,    -5,     0,    -2,     0,    -1,     1,    -4,    -1,     0,    -1,    -2,     1,    -2,    -2,     0,    -1,     0,    -1,     1,     3,     1,     2,     2,     0,     1,     2,    -2,    -5,    -4,     1,     4,     0,     0,     0,     2,     0,     3,     0,     3,     0,     3,    -2,    -1,    -2,    -3,     0,    -1,     2,     1,     0,    -1,     0,    -4,    -1,     1,     2,    -3,     1,     5,     1,     0,     0,    -2,     2,    -1,    -3,    -2,     2,     0,     1,    -1,    -1,    -1,    -1,    -2,     1,    -1,     0,     0,    -2,    -5,     0,     1,     0,     4,     4,     1,    -1,     1,     0,    -1,     0,     0,    -2,    -2,     1,     1,     0,    -1,    -2,    -2,    -1,    -3,     1,     0,    -1,     0,    -3,    -2,     2,    -1,     1,     2,     5,     4,    -1,     0,     0,    -1,     0,     0,    -3,    -2,     0,     0,     0,    -2,    -4,    -4,    -1,    -2,     1,    -2,    -1,     1,    -1,    -1,     0,    -1,     0,    -2,    -1,     0,    -1,     1,    -1,    -2,     1,    -1,    -2,    -1,     1,    -1,    -1,    -2,    -4,    -3,     0,    -1,     2,     0,    -2,     3,    -1,    -3,    -1,     0,    -1,    -2,    -2,     0,    -1,     1,     0,     0,    -2,    -2,    -2,    -2,     2,    -1,    -1,    -3,    -1,    -4,    -2,    -1,     0,     1,     0,     0,     1,     0,     1,     1,     0,    -1,    -4,     0,     0,     0,     0,    -2,    -2,     0,     0,    -1,     2,     1,    -1,    -2,    -6,    -3,    -1,     3,     1,    -1,    -1,     0,     1,     0,     0,    -1,     2,     0,    -4,    -2,     0,     0,     0,     0,    -1,    -2,     0,     1,     0,     1,    -2,    -3,    -4,    -3,    -1,     1,     1,    -1,    -3,    -1,     3,     0,     1,     1,     4,    -2,    -2,     1,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     0,    -1,     0,    -1,    -5,    -1,     1,     1,     0,    -1,    -3,     1,     2,    -2,     3,     0,    -2,    -4,     1,     0,     0,     0,     0,     0,     0,    -2,    -1,    -1,    -2,     1,    -1,    -2,    -2,    -1,    -1,     1,     2,     0,     0,     1,     1,     1,     1,     3,    -2,    -4,     0,    -1,     1,     0,     1,     0,     0,    -1,     0,    -1,    -1,     1,    -1,    -2,    -2,     0,     2,    -3,    -2,    -2,     1,     1,     1,     3,     1,    -1,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,    -2,    -1,    -1,    -7,    -8,    -7,    -4,    -1,    -2,    -4,    -5,    -5,    -6,     0,    -2,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -3,    -2,    -2,    -2,    -1,    -3,    -4,    -3,    -2,    -3,    -3,    -3,     0,     0,     0,     0,     1),
		    65 => (    0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,    -1,    -3,    -3,    -3,    -4,    -2,    -2,     2,     0,     1,     3,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -1,    -1,    -2,    -2,     1,    -1,    -2,    -1,    -1,     1,    -2,     2,     2,     2,     4,     4,     3,    -3,    -2,     1,     4,     0,     0,     0,    -1,    -1,    -1,    -1,    -4,    -2,    -3,     2,     2,     0,     0,    -4,    -2,    -1,    -4,    -1,     2,    -2,    -2,     1,     0,    -1,     0,     3,     2,    -2,     0,     0,    -2,    -2,    -1,    -2,    -7,    -7,    -2,     3,     1,     0,     1,     3,    -1,    -7,    -3,    -2,    -3,    -1,     3,     2,     2,    -2,    -2,     2,     3,    -1,     0,    -1,     3,    -1,    -2,    -5,    -6,    -7,    -3,    -1,     2,    -1,     3,     3,     0,    -2,    -2,     0,    -1,     1,     3,     1,     3,     0,     0,     5,     6,     2,     1,    -1,     3,    -3,    -2,    -2,    -6,    -6,    -3,     2,     0,     0,     3,     2,    -2,     2,     3,     3,     3,     4,     4,     1,     3,     0,    -1,     2,     6,     0,     0,    -1,    -2,    -2,    -1,    -6,    -5,    -3,     0,    -1,    -2,    -1,     0,    -2,     0,     2,     3,     3,     6,     4,     3,    -1,     1,     2,     0,    -1,     3,     2,     0,     0,    -4,    -4,    -4,    -4,    -2,    -2,    -3,     0,    -1,    -1,    -2,    -1,    -3,    -3,    -2,     3,     1,     0,    -3,    -2,     0,    -1,    -1,     2,     0,     3,     1,    -1,     0,    -1,     1,    -2,    -1,    -4,    -2,     1,    -2,     0,     0,    -2,    -4,    -9,   -10,    -8,    -6,    -8,    -7,    -3,    -3,    -7,    -3,     0,     3,     4,     0,     0,     0,    -1,     4,     0,    -4,    -3,    -2,     0,     0,    -1,     0,    -1,    -2,    -6,    -8,   -11,   -10,    -9,   -10,    -6,    -5,    -6,    -4,    -2,     1,     3,     0,     0,     0,     1,     2,    -2,    -4,    -1,    -1,    -1,     1,     0,     0,     3,     1,     0,    -2,    -4,    -3,    -4,    -5,    -7,    -7,    -5,    -4,    -2,     0,    -2,     0,    -1,     0,     2,     1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     2,     2,     1,    -2,    -2,    -2,    -2,    -1,    -5,    -9,    -5,    -4,    -1,     0,    -2,     0,    -1,    -1,     3,     1,    -2,    -1,     1,     1,     1,     0,     1,     1,     0,    -1,     1,    -2,    -1,    -2,     0,     3,    -1,    -2,    -2,    -2,    -1,     0,     0,     1,    -1,    -3,    -2,     1,     0,     2,    -2,    -1,     2,     0,     0,     1,    -2,    -1,    -1,     1,    -1,     0,    -1,     1,     3,    -1,    -1,     1,     0,    -1,    -2,     0,    -1,    -2,    -2,    -1,     0,    -2,    -3,     0,     0,     1,     2,     0,     2,     0,    -2,     0,     1,    -3,     0,    -1,    -1,    -3,    -4,     0,    -2,    -3,    -2,     0,    -1,    -2,     0,     0,    -3,    -3,    -1,    -2,    -1,     2,     2,     1,     2,    -1,    -1,    -1,    -1,    -1,     0,     1,    -2,    -3,    -5,    -1,    -2,    -1,    -3,     0,    -1,    -2,     1,     1,     0,    -4,    -6,    -4,    -5,    -3,     2,    -1,    -1,    -3,    -3,     2,     1,     1,     0,     3,    -2,    -2,     0,     1,    -1,    -3,    -2,     1,     0,    -2,    -3,     4,     0,     0,    -3,    -3,    -7,    -6,    -7,    -3,     0,    -2,    -4,     0,     2,     1,    -1,     2,    -2,    -2,     2,     2,    -1,     0,    -1,     0,    -1,    -1,    -1,     1,     2,     1,     0,    -1,    -4,    -1,    -3,    -5,    -1,    -1,     1,    -2,     1,     1,     2,     2,    -1,     0,     1,     0,    -1,    -1,     0,     0,     0,    -3,     0,     3,     2,     0,     0,     0,     1,     1,     0,     0,     2,     1,     0,    -1,    -1,     1,     3,     1,    -2,     2,     1,    -1,    -1,    -2,     0,     1,     0,    -3,     3,     1,    -2,    -1,    -2,     1,     4,     3,     2,     1,    -2,     1,    -1,    -1,     1,     0,     0,     1,     0,     0,     4,     0,    -1,     0,    -1,     0,     0,     1,     4,     4,     2,     2,     0,     1,    -2,     1,     2,     1,     0,    -1,     0,    -2,    -1,    -1,     0,     1,     0,     1,     4,    -1,    -2,     0,     0,     1,     0,    -2,     1,    -1,    -1,     0,     0,    -1,     0,     1,    -1,    -1,     0,     0,     0,    -2,    -1,     2,    -1,    -2,     1,     5,     1,     2,    -3,    -2,     0,    -1,    -1,    -1,     5,    -3,    -4,    -1,    -2,    -3,     0,    -2,    -2,     0,     3,    -1,    -1,    -6,     1,     1,     1,     2,     4,     6,     3,     2,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -3,    -1,     2,     3,     1,    -5,    -6,    -5,    -5,    -3,     1,    -2,     2,     1,    -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,     1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -2,    -1,     0,     0,     1,     0),
		    66 => (    0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     0,     2,     3,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     1,     1,     0,     3,     0,     1,     3,    -1,    -1,    -1,     1,     2,     3,     3,     2,     2,     2,     0,     1,     0,     0,     0,    -1,     0,    -1,     1,     2,     1,     0,     1,     2,     2,     2,     1,     2,     2,    -1,     2,     2,     3,     4,     3,     2,     6,     4,     3,     2,     0,     0,     1,     0,    -3,     2,     0,     3,     4,     4,     5,     5,     6,     6,     8,     5,     7,     5,     1,     1,     1,     0,    -2,    -2,    -2,     0,     2,    -5,    -4,     0,     0,     0,    -3,     0,     2,     3,     3,     5,     2,     5,     5,     2,     4,     1,     5,     4,     1,     2,     1,     3,     3,     2,    -1,    -1,    -2,    -3,    -1,     4,    -1,     0,    -1,    -3,     4,     2,     3,     3,     2,     2,     4,     1,    -2,     2,     4,     2,     1,     3,     0,    -1,     1,    -3,     0,     0,     4,     2,     3,     1,     0,     0,     0,     0,     3,     1,     4,     2,    -1,     1,    -1,    -2,     1,     1,     1,     0,     0,     0,    -4,     1,     0,    -2,    -2,    -2,    -1,     1,     3,     4,     0,    -1,     0,    -1,     3,     2,     1,     1,     0,    -1,    -2,    -1,    -3,    -4,     1,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     1,     0,     3,     3,     0,    -1,    -2,    -7,     4,     1,     1,    -1,     0,     2,    -2,    -2,    -1,    -2,     0,    -3,    -5,    -2,    -1,     0,     1,     1,    -1,    -2,    -2,    -5,     0,    -4,     0,    -1,    -2,    -4,     3,    -1,    -2,    -1,     0,    -1,    -2,    -2,    -3,    -4,     0,     0,    -2,    -5,    -1,    -1,     0,     3,     0,    -1,    -4,    -6,    -4,    -4,     0,    -1,    -3,    -2,     1,     0,    -2,    -2,    -1,    -1,    -1,    -3,    -4,    -2,     0,    -2,    -4,    -3,    -4,    -3,     0,     0,    -3,    -3,    -4,    -5,    -4,    -4,     0,    -1,     0,    -4,     1,     1,     0,    -1,    -2,    -1,    -2,    -3,     0,     0,    -1,    -3,    -2,    -2,    -2,    -1,    -1,     0,    -3,    -1,    -2,    -4,    -4,    -3,     1,    -1,    -2,    -4,    -1,     1,     3,     1,    -1,     1,     0,     0,    -1,     2,    -2,    -1,    -3,    -2,    -3,    -2,     2,     1,    -2,     2,     3,     0,    -6,    -3,     0,     0,    -1,    -3,    -1,     1,     0,    -2,    -1,     3,     3,     2,     2,     1,     1,     1,    -1,    -4,    -1,     2,     2,     2,    -1,     2,     1,    -2,    -6,     0,     0,     0,    -1,    -3,    -5,     1,    -2,    -3,     1,     1,     3,     3,     3,     2,     1,    -2,     0,    -2,     1,     1,     1,     1,     1,    -2,    -1,     3,    -5,    -1,     0,     0,    -2,    -2,    -5,    -2,    -2,    -1,    -2,    -1,     1,     2,     0,     4,     3,    -2,    -2,    -4,     0,     2,     0,     1,    -3,     0,     0,     3,    -2,    -6,     0,     0,    -3,    -2,    -1,     1,     1,     1,    -1,     2,     2,     1,    -1,    -2,    -1,    -1,    -1,    -2,     3,     3,    -1,    -1,     1,     0,    -1,     2,    -3,    -5,    -1,     0,    -3,    -3,    -2,     3,     0,     1,    -1,    -2,    -1,    -1,    -1,    -2,     0,     1,     1,     2,     2,     2,     2,    -1,    -1,    -1,    -1,     2,    -3,    -7,     0,     0,    -3,    -5,    -1,     0,    -2,     0,     0,     1,     2,    -4,     0,     0,     0,    -2,     0,     2,     5,     4,     0,    -2,     0,     1,     1,     3,     0,    -3,     0,     0,    -4,    -4,     1,     2,     1,    -1,     0,     0,     4,     4,     2,     1,     1,     1,     0,     3,     0,     4,     0,     0,    -1,    -2,    -3,     1,    -2,     0,     0,     0,    -4,    -5,     0,     0,     0,     2,     1,     1,     3,     4,     3,    -2,     1,     1,     1,     2,     2,     2,     2,     0,     0,    -4,    -5,    -1,    -1,     0,     0,    -1,    -4,    -5,    -4,    -4,    -1,     3,     4,     0,     2,     0,     5,     2,     1,     1,     4,     3,     2,     1,     1,    -1,    -1,    -4,    -2,     0,     0,    -1,     0,     0,    -3,    -4,    -7,    -8,   -11,     0,     0,     2,     1,     1,     0,     0,     0,     3,     3,     5,     3,     0,     1,     1,    -3,    -3,    -7,    -2,    -1,    -1,     0,     1,     1,    -4,    -5,    -6,    -5,    -1,    -1,     0,    -2,     1,     3,    -1,     1,     3,     0,    -2,     1,     0,     0,     2,    -4,    -5,    -5,    -3,    -4,     1,    -1,     0,     0,    -1,    -2,    -2,    -3,    -5,    -7,   -10,    -7,    -8,    -4,    -4,    -3,     1,     1,     2,     4,    -7,    -1,    -3,    -3,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -2,     1,     2,    -1,    -1,    -2,    -3,    -3,    -2,    -5,    -4,    -1,    -2,    -2,    -2,     1,     0,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,    -1,     0,    -1,    -1,     1,    -1,    -1,     0,     0,     0,     1,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,    -1,     0,     0,     0),
		    67 => (    0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     1,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,    -1,     1,     0,    -2,    -4,    -2,    -2,    -2,     1,     0,    -1,    -1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -3,    -2,    -1,    -2,    -2,    -4,    -4,    -3,    -3,    -2,    -2,    -1,     0,    -1,     1,    -1,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,    -2,     0,    -3,    -3,    -4,    -5,    -7,     0,     1,     0,    -1,    -3,    -7,    -5,    -4,    -4,    -3,     0,    -2,    -3,    -3,    -2,    -1,     0,     0,     0,     0,    -2,    -2,    -1,    -5,     0,     5,     1,    -1,     0,     2,    -1,     2,     0,     1,     0,     4,     0,    -3,    -1,    -1,    -2,    -4,    -1,    -1,     0,     0,     0,     2,    -1,    -1,    -1,    -3,     1,     2,     3,     2,    -1,    -1,    -1,    -1,     1,     1,     0,     2,     1,    -5,    -2,     0,    -2,    -3,    -2,    -2,    -1,     0,     1,     2,     0,     1,     0,     1,     1,     2,     1,     0,    -1,    -2,    -3,    -3,     0,     2,     2,     2,     3,     5,     1,    -2,    -2,    -3,    -2,    -2,    -1,    -3,     1,     5,     0,     2,     1,     1,     3,     3,     0,    -1,    -1,    -1,    -2,     0,     3,     1,     1,     1,     1,     3,     2,     0,    -4,    -3,    -1,    -1,    -1,     1,     1,     1,     2,     2,    -3,    -1,     0,     1,     0,     1,    -2,    -1,     1,     0,    -1,     1,     3,    -1,    -1,     1,    -2,    -1,    -3,    -2,     0,    -2,     1,     1,     0,    -1,     1,     3,    -1,    -1,     1,    -1,     1,     1,    -2,    -4,     1,     0,     1,     0,    -1,     0,     1,    -1,    -3,    -1,    -2,    -2,     0,    -2,     0,     1,     1,     0,    -2,     0,     0,    -1,     2,     1,    -1,     0,     0,    -4,    -3,     0,     4,     0,     0,     0,     0,    -3,    -2,    -2,    -5,    -3,    -3,    -2,     1,     0,     0,    -2,    -1,    -2,    -1,    -2,     2,     0,    -3,    -2,    -5,    -5,    -3,    -2,     2,    -1,    -3,    -1,    -4,    -3,    -2,    -5,    -5,    -5,    -1,    -1,     0,     0,     2,     2,    -1,    -1,    -1,    -2,     0,     0,    -2,    -3,    -4,    -9,    -6,    -3,    -1,    -2,     0,    -1,    -4,    -3,    -3,    -4,    -6,    -5,    -1,    -3,    -1,     0,     2,     1,     2,     0,     2,    -3,    -2,    -3,    -5,    -9,    -7,    -5,    -3,    -3,     0,    -2,     1,     2,     1,    -1,     1,    -3,    -4,    -1,    -1,    -2,    -1,     0,     0,     0,     2,     1,    -1,    -2,    -6,    -4,    -3,    -5,     0,    -1,    -1,    -3,     0,     0,     2,     3,     1,     2,     1,    -1,     0,     0,     1,    -1,    -1,     0,     0,     0,    -2,    -1,     0,    -4,    -2,     3,    -1,    -1,     3,     1,     0,    -1,     3,     1,     0,     2,    -1,     0,    -3,    -2,    -1,    -1,    -4,    -2,    -1,     1,     0,    -2,    -2,    -2,    -4,    -2,    -2,    -1,     0,    -3,     0,    -1,     0,    -1,     1,     1,     2,     1,     0,    -4,    -5,    -4,    -3,    -1,    -6,    -3,    -4,     1,     0,     1,    -2,    -2,    -1,    -2,     0,    -1,     1,     0,     0,    -3,     2,     1,     3,     0,     4,    -2,     1,     2,     0,    -3,    -4,    -2,    -5,     0,    -3,     0,     0,     0,     0,    -1,    -4,    -2,    -2,     1,    -1,    -1,    -3,    -1,    -1,     3,     4,    -2,    -2,    -1,     1,     2,     2,    -1,     0,     1,    -2,    -2,    -2,     0,     2,    -1,     0,    -1,    -3,    -3,     0,     1,     1,    -1,    -6,    -2,    -1,     1,     1,    -2,    -3,    -1,    -1,     2,     0,    -2,    -5,    -3,    -1,    -3,     0,    -1,     0,    -1,    -1,    -1,    -4,    -5,    -4,     1,    -1,    -2,    -3,    -1,     0,     2,     1,     3,    -4,    -2,    -2,    -1,     0,    -2,    -6,    -3,    -3,     0,     0,    -1,     0,    -1,     0,    -1,    -3,    -4,    -4,    -2,    -3,    -2,    -3,    -2,     2,     1,     2,     1,     1,    -2,    -1,    -2,    -5,    -8,    -6,    -3,    -2,    -3,     0,     0,     1,    -1,    -2,    -4,    -4,    -4,    -6,    -5,    -7,    -5,    -4,    -2,    -1,    -1,     0,    -1,    -4,    -6,    -4,    -4,    -4,    -4,    -3,     1,    -2,    -3,    -1,    -1,    -1,     0,     0,    -2,    -4,    -5,    -5,    -8,    -7,    -5,    -4,    -1,     0,     1,     3,    -1,    -1,    -5,    -3,     0,    -1,     0,    -2,    -2,    -2,     0,     0,     0,     0,    -3,     0,     0,    -2,    -3,    -4,    -4,    -6,    -4,     1,    -2,    -2,    -1,     3,     0,     1,     0,     2,     2,     2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     2,     1,     1,    -2,    -1,     2,     2,     1,     1,     0,     1,     7,     6,     4,     1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     3,     3,     2,     2,     2,     1,     3,     2,     4,     6,     4,     2,     0,    -1,     1,     0,    -1,     0,    -1),
		    68 => (    0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     1,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -3,    -2,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -1,     0,     0,     1,    -1,    -1,     0,     1,     1,     0,     0,    -1,     0,     1,     0,     0,    -1,    -1,    -1,    -2,    -2,     0,     0,     0,     2,     2,    -1,     0,    -3,    -3,    -1,     1,     0,     1,    -1,    -1,     0,    -1,     0,     0,     0,    -1,    -1,     0,    -1,    -3,    -3,     0,     0,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -1,     1,     0,    -1,    -1,     0,    -1,    -3,     0,     0,     0,     1,     0,    -1,    -2,    -3,    -1,    -3,    -2,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,     1,     3,     1,     1,     0,    -1,    -1,    -2,     0,     0,     1,     1,     1,     1,     0,     1,    -2,    -1,     1,     0,     1,     0,     0,    -1,     0,    -1,     0,     2,     4,     4,     1,     0,    -2,    -2,    -1,     1,     0,     1,     0,    -2,    -2,    -1,    -1,    -1,     0,     0,     1,    -1,    -1,     0,    -1,     0,     0,    -2,    -2,     2,     3,     4,     1,    -1,    -3,    -2,     1,    -2,    -2,    -1,    -2,    -3,    -3,    -1,    -1,     1,     2,     2,     0,     0,     0,     2,    -1,    -1,     0,    -1,    -2,     1,     1,     3,     2,     1,    -2,     0,     1,     0,     0,    -1,    -1,    -2,    -1,     0,    -1,     0,     1,     0,    -1,    -1,     0,    -2,    -1,    -1,     0,     0,    -3,    -1,    -1,     0,     2,     3,     2,     3,     2,     1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,     0,    -1,    -1,     0,    -1,    -1,    -1,     0,    -2,     0,     0,    -2,    -4,    -3,    -1,     0,    -1,     1,     1,     2,     0,     0,    -3,    -3,     0,     0,    -1,     0,    -2,    -2,     1,     0,    -1,    -1,    -2,    -2,    -3,     0,    -1,    -3,    -4,    -2,    -2,    -2,    -2,    -2,    -2,    -1,     0,     0,    -1,     1,     1,     0,    -2,    -1,    -3,    -2,     0,     0,    -1,    -2,    -3,    -2,     1,    -1,    -1,     1,    -4,    -2,    -1,    -2,    -3,    -3,    -4,    -2,    -3,    -2,     0,    -1,    -2,    -2,     0,     0,    -1,    -2,    -1,     0,     0,    -2,    -1,    -4,     0,     0,     1,    -1,     1,     0,    -1,    -2,    -3,    -2,    -2,    -2,    -1,    -1,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -2,    -1,    -1,    -2,     1,    -2,    -2,     0,    -1,     0,     1,     0,    -1,    -2,    -1,    -1,    -2,     0,     1,     0,    -1,    -3,    -3,     1,     1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -2,    -1,     1,     0,     0,     2,    -1,    -1,    -1,    -1,    -2,    -2,     2,     2,     0,    -2,    -2,    -3,    -2,     1,     0,    -1,    -1,     1,     1,    -2,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,     1,     0,     1,     0,    -3,    -2,    -2,     2,     1,    -1,    -2,    -1,     2,    -1,    -1,     0,     0,    -2,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -3,     0,     1,     2,     0,     0,    -2,    -2,    -2,     0,     2,     1,    -1,     0,     1,     1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -2,     0,     1,     2,     1,    -2,    -3,    -2,    -3,    -1,     1,     0,     0,     0,     2,     1,    -1,     0,    -2,     0,    -1,    -1,     0,    -2,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     1,     1,     0,    -1,    -1,    -2,     0,     1,     0,     0,     0,     2,     0,    -1,    -1,    -1,     0,    -2,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,     0,     0,    -1,    -1,    -1,    -1,    -2,     1,     0,     0,     0,     1,     1,    -1,    -2,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,    -2,    -1,     1,    -1,     0,     1,     0,    -1,     0,     1,     2,     1,    -1,     0,     0,    -3,     0,     0,     1,    -1,     0,     0,    -1,    -1,     1,    -1,     0,     0,    -2,    -2,    -2,     1,     1,     2,    -1,    -3,    -2,     0,    -2,    -2,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,     2,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -2,    -2,    -1,    -2,    -2,    -1,     0,     0,    -3,    -3,     0,    -2,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,     0,     0,     0,    -1,     0,     0,     0,    -1,     0),
		    69 => (    0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -3,    -1,    -3,    -3,    -3,    -2,     0,     0,     0,    -2,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -3,     0,     0,    -3,    -3,    -1,    -2,    -2,     0,     0,    -7,    -4,    -4,    -2,    -4,    -3,    -5,    -6,    -4,    -4,    -2,    -1,     1,     0,     0,     0,     0,    -3,    -4,    -3,    -2,    -4,    -8,   -10,   -13,   -12,    -8,   -10,   -10,   -10,   -14,   -12,    -4,    -5,    -8,    -7,    -6,    -3,    -3,    -2,     1,     0,     1,     0,    -2,    -3,    -4,    -6,    -8,    -5,    -6,    -7,    -4,    -1,     0,    -1,    -2,    -2,    -2,    -4,    -7,   -14,    -9,    -7,    -7,    -4,    -3,    -5,    -4,     0,     0,     0,    -2,    -2,    -2,    -3,    -3,    -2,    -5,     1,     1,     0,     2,     4,     1,     2,     3,     3,     0,    -2,    -4,    -2,    -8,    -3,    -5,    -5,    -4,    -1,     0,     1,    -2,    -5,    -4,    -5,    -3,    -2,     0,     3,     3,    -1,    -1,     4,     2,     4,     6,     4,     1,     1,    -1,     0,    -1,     1,     0,    -2,    -4,    -5,     0,    -2,    -3,    -5,    -3,    -5,    -1,    -1,    -1,     1,     1,    -1,     2,     5,     4,     4,     7,     4,     0,     1,     2,     0,     1,     1,     0,     0,    -4,    -4,    -3,    -4,    -3,    -4,    -4,     0,     1,    -1,     0,     1,     0,     0,     3,     3,     4,     6,     5,     3,     3,     4,     0,     2,     1,     2,     2,     0,    -4,    -2,    -1,    -3,    -4,    -4,     3,     1,     3,     1,     1,     3,     1,    -1,     1,     4,     3,     2,     2,     1,     1,     1,     3,     0,     0,    -1,    -1,    -4,    -5,    -4,     0,    -2,    -6,    -3,     3,     3,     0,     0,     0,     0,     0,     0,     2,     1,     1,    -3,     0,    -2,     0,     0,     1,    -3,    -2,    -1,    -3,     2,    -6,    -2,     0,    -9,     0,    -2,     1,     3,     1,    -1,    -3,    -1,    -1,    -2,     0,    -3,    -3,    -3,     0,     1,    -2,    -1,     2,    -1,    -4,    -3,    -3,     0,    -5,    -2,     0,    -1,    -1,    -2,     2,     1,     1,    -1,    -3,    -3,    -1,     0,    -3,    -3,    -2,    -3,    -1,     1,    -2,    -3,     1,    -2,    -2,     0,    -4,    -7,    -4,    -3,    -1,    -2,    -3,    -2,     1,    -1,     1,     1,     0,    -2,     0,    -2,     0,    -1,    -2,    -3,     1,     0,    -1,    -1,    -2,     0,    -2,    -2,    -2,    -5,    -3,    -1,    -1,    -2,    -2,     0,     1,    -1,     0,     1,     0,     0,     0,    -1,     2,    -3,    -2,     1,     0,     0,     1,     1,     0,    -2,    -3,    -6,    -2,    -6,    -3,     0,     0,     0,    -4,    -2,     1,     0,     1,     0,     2,     1,    -2,    -3,    -2,    -1,     1,     1,     2,     1,     2,     3,     4,     1,     1,    -4,    -2,    -6,    -1,    -4,     0,    -1,    -3,    -2,     0,     2,     2,    -1,     1,     0,    -1,    -3,    -3,    -1,     3,     2,     0,     3,    -1,     2,     3,     1,     0,    -3,    -1,    -7,    -4,    -4,     0,     0,    -4,     0,    -3,     1,    -2,    -1,     0,     1,    -1,    -2,    -1,    -1,     2,     1,     0,     1,    -2,     0,     1,    -1,    -6,    -7,    -2,    -8,    -5,    -3,     1,     0,    -5,     4,    -2,    -2,     0,     0,    -4,    -2,    -2,    -3,    -4,    -1,    -2,    -1,     2,     1,    -4,     1,     0,    -3,    -2,    -2,    -3,    -7,    -4,    -2,     0,    -1,    -4,     2,     0,    -2,    -3,    -1,    -4,    -2,     0,    -1,    -1,    -2,     0,    -2,     1,    -1,    -1,     0,     0,    -3,     0,     2,    -1,    -4,    -3,    -1,     0,    -1,    -8,     1,    -3,     1,     0,    -5,    -1,    -2,    -1,    -2,    -3,    -2,    -2,    -2,     1,     0,    -2,     1,    -2,    -3,     0,     4,     4,     2,    -2,     0,     1,     0,    -7,     1,    -1,     1,     1,    -1,    -2,    -3,     1,    -1,    -2,    -2,     0,    -1,     3,     2,    -1,    -2,    -4,    -1,     1,     3,     3,     0,    -6,     0,     0,     0,    -5,     2,    -2,     0,    -1,    -2,     0,    -2,     0,    -3,     1,    -1,     2,     0,     3,     3,     0,    -2,    -1,     1,     4,     4,     3,    -5,    -5,     0,     0,     0,    -1,     1,    -2,     0,     1,     4,     2,     0,    -1,     0,     0,     1,     3,     3,     2,     1,     1,     0,    -1,     0,     1,     3,     5,    -2,    -3,     0,    -1,     0,    -2,    -3,    -1,     2,     4,     6,     3,     2,     1,     2,     1,     1,    -3,    -2,    -2,     1,     5,     3,     3,     1,    -2,     1,     1,    -2,     0,     0,     0,     0,     2,    -3,    -1,     2,     4,     5,     3,     3,     0,     1,    -1,    -2,     2,    -1,     0,     4,     3,     1,     3,    -1,     0,    -2,     0,     0,    -1,     0,     0,     0,     0,     2,     0,     1,     3,     5,    -1,     1,     0,    -2,     1,    -1,     3,     3,     1,     0,     2,    -1,     5,     1,    -1,     3,     1,     0,     1,     0,     0,     0,     0,     0,     0,    -2,     1,     1,     1,     0,     1,     2,     2,     1,     2,     1,     2,    -3,     0,     1,    -2,    -4,    -3,    -2,     0,     0,     1,    -1),
		    70 => (    0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -2,    -1,     1,    -1,    -2,    -1,    -1,     0,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     1,    -1,    -1,     0,     1,    -1,    -1,    -1,    -5,    -3,    -2,     0,     2,     1,    -3,    -1,     0,     0,     0,    -1,    -3,    -3,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,    -1,    -4,    -1,     0,    -2,    -1,    -1,     3,     3,     4,     2,     1,    -3,    -4,    -1,     1,    -3,    -4,    -2,    -1,    -1,    -2,    -1,     0,     0,     0,    -1,     0,    -1,    -3,    -1,     0,     0,     0,     0,     1,     4,     1,     1,     2,    -1,    -4,    -3,     2,    -2,    -4,     0,     1,     0,    -3,    -2,    -2,     1,    -1,     0,    -1,     1,     1,     2,     1,     2,     0,     0,     4,     1,    -1,     0,     0,     2,     2,    -2,     0,    -1,    -1,     0,    -1,    -1,    -4,    -2,    -1,     0,     0,    -1,    -2,     0,     2,     2,     2,     1,     2,     0,     2,     0,     1,     3,     2,     3,     1,     1,     1,     2,     1,    -2,    -1,    -1,    -1,    -2,    -2,     1,     0,     2,    -2,     2,     0,     1,    -1,     0,     2,     2,    -1,    -1,     2,     2,    -1,    -2,    -2,     2,     0,     1,     2,     0,     0,    -2,    -1,    -4,    -2,     1,     0,     3,     0,    -1,    -1,    -3,    -2,     2,     2,     3,     0,    -1,     2,     0,     0,    -1,     0,    -1,     3,    -1,    -1,    -1,    -1,    -3,    -2,    -3,     1,     0,     0,     3,     1,    -2,     0,    -2,    -2,     1,     1,     0,     0,     0,    -3,    -1,     2,     0,    -1,    -2,    -2,    -3,    -2,    -1,     2,    -1,    -1,    -2,     0,     0,     3,     0,    -2,    -2,     0,    -1,    -2,     0,    -1,     1,    -2,    -5,    -7,    -5,    -1,    -2,    -2,    -2,    -3,    -1,    -1,    -1,    -1,     1,    -1,    -1,    -1,     0,     0,     0,    -1,    -2,    -3,    -1,    -3,    -1,     0,    -2,     0,    -6,    -7,    -8,    -4,     2,    -1,    -2,    -1,     0,     0,     0,    -1,    -3,    -2,    -2,    -1,     0,     1,     1,     2,    -1,     0,     0,    -2,    -1,     1,     1,     0,    -4,    -7,    -3,    -2,     0,     1,    -1,    -1,     1,     2,    -1,    -1,    -3,    -2,    -3,    -1,     0,     0,    -1,     2,     1,     0,    -1,    -1,    -2,     2,     4,     0,    -4,    -3,    -2,    -3,    -3,     0,     1,     0,     0,     2,     1,    -1,    -2,     0,    -3,    -1,     0,     0,    -1,     1,     2,     1,    -4,    -1,     1,     3,     5,     0,    -2,    -4,    -1,    -3,    -6,     0,     0,    -1,     2,     1,     2,    -2,    -2,     2,    -2,    -2,     0,     0,     0,     1,     1,    -2,    -3,    -2,     0,     1,     2,     2,    -3,    -2,    -2,    -2,    -7,     0,    -1,    -1,     2,    -1,     1,    -1,    -3,    -1,    -5,    -1,     0,    -1,    -1,     1,     1,    -1,    -3,    -1,     0,     1,     2,     1,    -1,    -4,    -5,    -9,    -4,     0,    -2,    -1,     1,    -1,     0,     0,    -1,    -2,    -4,     0,     0,     0,    -1,     0,     0,    -2,    -3,    -2,    -2,     1,     3,     1,    -1,    -3,    -7,    -8,    -5,    -3,     3,     0,     2,    -1,     0,     0,    -2,    -2,    -3,    -1,     0,     1,    -1,    -1,    -1,    -1,    -3,    -2,    -1,     3,     1,    -1,     1,    -2,    -3,    -2,    -1,    -1,     0,     0,     1,     0,    -2,     0,     0,    -5,    -1,     0,     0,     0,     0,    -1,     1,     2,    -3,    -2,    -2,     0,     1,     3,    -2,    -1,     3,     0,    -1,    -1,     0,    -2,     0,     1,    -2,     1,     0,    -4,     1,     1,     0,     0,     0,    -1,    -1,     0,    -5,    -1,    -2,    -1,     0,     2,     2,     2,     2,     2,    -2,    -2,    -1,     0,     2,     0,     0,     1,     1,     0,     1,     2,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -1,     2,     0,     1,     2,     0,     1,    -1,     0,     1,     2,     1,     1,     1,    -1,     0,     1,     1,     0,     0,     0,    -2,     0,    -1,    -3,    -4,    -1,     2,    -1,    -1,    -1,     2,     1,     3,     4,     4,     1,    -2,    -2,    -1,    -1,    -2,     1,    -2,    -1,     0,     0,     0,    -1,     0,     2,    -1,    -2,    -2,    -3,    -1,    -1,    -1,    -1,    -1,    -2,     0,     0,     1,     0,    -2,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,    -1,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,     0,    -5,    -3,    -4,    -2,    -3,    -3,    -2,    -2,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,     0,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -2,    -2,    -4,    -4,    -1,    -3,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     1,    -1,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0),
		    71 => (    0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     2,     1,     1,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -2,    -1,    -1,    -3,    -2,    -2,     0,     3,     0,    -1,    -1,    -2,    -5,    -3,    -2,    -1,    -1,     0,     0,     0,     0,     3,     0,     0,    -1,    -1,     0,    -2,    -3,    -3,    -4,     0,     0,    -4,    -1,     2,     2,     2,     2,     2,     3,    -1,     0,    -1,     0,     0,     1,     0,     0,     3,     3,     1,     1,     0,     0,     1,     0,     1,     0,     0,     1,    -2,    -3,     0,     1,     2,     3,    -1,     2,    -1,     0,    -1,    -2,    -3,    -1,     1,     0,     2,     0,     1,     1,     0,    -1,    -2,    -1,    -1,     0,     2,     0,     2,     2,     1,    -3,     0,     2,     1,     1,     1,     1,    -1,    -2,    -1,    -1,     0,     0,    -2,    -2,    -1,     1,     0,     0,    -5,    -8,    -3,     0,    -1,    -1,    -1,    -1,     0,    -3,     2,     0,     0,     2,     1,     1,     0,     0,    -1,    -1,     0,     0,    -2,    -2,    -3,     1,     1,    -3,    -5,    -2,     0,    -2,    -1,    -2,     0,    -3,    -2,    -1,     1,     1,     1,     3,     1,    -1,    -1,     0,    -3,    -1,     0,    -1,    -3,    -2,    -3,    -1,     3,     1,    -4,    -2,     0,    -1,     2,     2,     0,    -1,    -2,    -2,    -3,    -4,     0,     2,     2,    -1,    -2,     0,    -3,     0,     0,     0,    -2,    -3,    -2,     0,     0,     2,     1,     0,    -3,    -1,    -1,     1,     0,     0,    -2,    -2,    -4,    -5,    -2,    -1,     1,     2,    -1,     3,     2,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -3,    -1,     2,    -1,    -3,    -1,     0,     3,     1,    -2,    -1,     0,    -3,    -1,    -3,    -4,     2,     2,    -1,     3,     2,     2,     0,     0,    -1,    -1,    -1,    -2,    -3,    -2,    -3,    -4,    -3,     0,     1,     0,    -1,    -3,    -2,     0,    -3,    -2,    -1,    -2,     2,     2,    -1,     2,     1,     4,     1,     1,    -1,    -1,     0,     0,     0,     0,    -3,    -1,    -1,     0,     2,     2,    -1,    -1,     0,     3,    -3,    -3,    -1,    -1,    -2,    -1,     0,     3,     4,     5,     0,     0,     0,     0,     0,     1,     1,     1,     2,     2,    -1,    -1,    -1,    -3,     0,    -1,     1,     1,    -5,    -4,    -3,    -3,    -3,    -4,    -3,     4,     3,     0,     1,     0,     0,     1,    -1,     1,     2,    -1,     5,     4,     1,    -3,    -4,    -3,     1,    -1,     2,     0,    -2,    -4,    -1,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -2,     1,     2,     4,     0,    -1,    -1,     0,    -1,     0,     1,     0,    -1,    -3,    -3,    -3,    -2,    -2,    -3,     0,     0,    -1,     0,     0,     0,    -2,     0,     1,    -2,     0,     2,     1,     1,    -3,     0,    -1,     1,    -3,     0,    -1,    -2,    -5,    -3,    -5,    -3,    -2,     0,    -3,    -2,    -1,     1,     0,     0,    -2,     0,     1,    -1,    -3,    -1,    -2,    -3,    -6,     1,     2,     1,     0,     0,    -2,    -5,    -4,    -2,    -3,    -2,    -1,    -1,    -2,    -2,    -3,     1,     0,    -1,     0,    -3,    -2,    -4,    -4,    -4,    -7,    -6,    -6,    -3,    -1,     3,     0,     0,    -1,    -4,    -2,    -2,    -2,    -2,    -2,    -3,    -1,    -2,    -1,     0,     0,     0,    -2,    -2,    -5,    -2,    -4,    -1,    -4,    -4,    -6,    -4,    -3,     3,     2,     0,    -1,    -2,    -1,    -2,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     1,     2,    -1,     1,    -1,    -2,     1,     1,     0,     1,    -3,     3,     2,     2,     1,     4,     1,     2,    -2,    -3,     0,     1,    -2,    -1,     0,     1,     0,    -1,     2,     3,     2,     3,     2,     0,    -1,     0,    -1,    -3,    -2,     1,     1,     3,     0,     3,     1,     3,     1,    -4,    -2,    -1,     0,    -2,     0,     1,     1,    -4,    -2,     4,     5,     3,     2,     1,    -2,    -3,    -2,     0,    -1,    -1,     5,     2,    -1,     1,     0,     1,     0,    -2,    -2,    -2,     0,     0,     0,     0,     1,    -1,    -2,     1,     0,     2,    -3,    -4,    -2,    -4,    -3,     1,     0,     0,     1,     0,     0,     1,    -1,     0,    -2,     0,    -1,    -1,    -3,     3,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -2,     2,     2,     0,    -1,    -4,    -4,     1,    -1,     1,    -2,    -6,    -3,    -2,    -3,    -2,    -3,     4,     4,     1,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -3,    -6,    -3,    -4,    -3,    -6,    -4,    -3,    -5,    -1,    -1,    -1,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,     0,     0,    -4,    -3,     1,     1,     3,    -4,    -1,    -1,     0,    -1,     0,     0,     1,     0,     1,     1,     0,     0,     0,     0,     1,     1,     0,     0,    -1,     1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0),
		    72 => (    0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -1,     1,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -3,    -2,    -3,    -3,    -2,    -3,    -2,    -2,    -1,    -2,    -2,    -5,    -4,    -1,    -1,    -1,     1,     0,     0,     0,     0,     0,    -1,    -1,    -2,     0,     0,    -3,    -1,     3,     3,     0,    -1,    -5,    -4,    -7,    -5,    -1,     0,    -1,    -6,    -2,    -2,    -1,     1,     1,     0,     1,     0,     0,    -1,    -2,    -1,     1,     0,     0,     1,     1,     2,     0,    -3,    -6,    -5,    -5,    -5,    -4,    -5,    -4,    -5,    -3,    -2,    -1,     0,     0,     1,     0,     0,    -1,    -2,     0,     0,    -1,     2,     1,     0,    -1,     2,     0,    -2,    -5,    -5,    -4,    -5,    -3,    -4,    -4,    -3,    -3,    -2,    -2,     0,     0,    -2,    -1,    -1,     0,    -1,     0,     1,    -2,     3,     3,     3,     0,     2,    -2,     1,     0,    -2,     0,    -5,    -5,    -4,    -2,    -1,    -3,    -4,    -1,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     1,     3,     2,     1,     2,     2,     0,    -1,    -1,     2,     0,    -2,    -3,    -3,    -3,    -1,    -1,    -3,    -3,    -2,    -3,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,     0,    -2,    -1,     0,     1,    -3,     0,    -1,    -1,    -2,    -2,    -3,    -1,    -3,    -3,    -3,    -4,    -4,    -5,    -4,    -2,    -2,    -1,    -2,     4,    -1,     0,    -3,    -1,     1,    -1,     0,    -1,     1,    -1,    -2,     2,     2,     0,    -1,    -1,    -2,    -3,    -5,    -5,    -4,    -4,    -5,    -2,    -3,    -1,    -1,    -2,    -1,     1,    -4,    -1,     0,    -1,     0,     0,     1,     0,     1,     0,     5,     1,    -1,    -2,    -3,    -3,    -3,    -3,    -6,    -2,     4,    -4,    -1,    -2,     0,    -1,    -1,    -1,    -5,     2,     0,     0,     0,    -2,    -2,    -1,     1,    -1,     1,     3,     2,    -2,    -3,    -2,    -2,    -3,    -3,     1,     2,    -2,    -3,    -2,     0,     0,    -4,    -1,    -2,    -1,    -1,    -1,    -2,     0,     1,     4,    -2,    -3,    -1,     1,     0,    -1,    -1,    -3,    -3,    -5,    -3,     0,    -1,    -3,    -5,    -1,     0,    -1,    -4,    -1,     0,     1,    -3,    -5,    -1,    -2,    -2,    -2,     0,     0,    -1,    -1,     1,    -1,     0,    -3,    -3,    -1,     1,    -4,    -1,    -1,    -2,     0,     0,    -1,    -3,     0,    -1,    -1,    -4,    -5,    -1,    -2,    -4,    -2,    -1,     0,    -2,     1,     0,     1,    -2,    -2,     1,     3,     4,     1,    -1,    -1,     3,     2,     0,     0,    -1,    -1,    -3,     0,    -4,    -3,    -1,    -3,    -1,    -1,     0,     1,     1,     1,     1,     0,    -2,     0,     1,     3,     2,     0,    -1,     0,     5,     2,     0,    -1,     3,    -2,    -1,     0,    -1,    -2,    -1,     0,     1,     0,     2,     3,     1,     2,     0,    -1,    -1,     0,     2,     0,    -2,    -3,     0,     1,     1,     3,     0,     0,     3,    -1,     2,    -2,     0,    -1,    -4,    -1,     1,     2,     0,     2,     1,     1,     3,     2,     0,     1,     0,     1,     1,     1,     1,     2,    -1,     3,    -1,     0,     4,     1,     2,    -1,     2,     0,    -1,     0,     2,     2,     0,     0,     2,     2,     2,     2,     2,     3,     2,     3,    -1,     1,     0,    -1,    -3,     3,     0,     0,     2,     2,     1,     1,     3,     0,    -2,     1,     2,     2,    -1,     1,    -1,     2,     1,     0,     2,     1,     1,     2,     2,     2,     4,     2,    -2,     2,     0,    -2,     0,     3,     0,     2,     1,     1,     0,     3,     1,    -1,    -2,    -1,    -1,     2,     0,     0,    -1,    -2,    -2,     0,     2,     4,     2,     1,     2,     4,     0,    -1,     1,     3,     0,    -1,     0,    -1,     1,     0,     0,     0,    -1,     0,     1,     0,    -3,    -4,    -4,    -4,    -3,    -1,    -2,    -1,    -1,    -3,     2,     0,     1,     0,     0,     1,     1,     1,     4,     0,     0,     0,     2,    -2,     1,    -1,    -2,    -2,    -6,    -9,    -1,    -2,    -3,    -4,    -4,    -5,    -5,    -3,    -2,     0,     1,     0,     0,     0,     0,     1,     1,    -2,    -2,    -2,    -3,    -1,    -1,    -2,    -2,    -5,    -8,    -8,    -2,    -1,    -3,    -5,    -6,    -4,    -4,    -4,    -6,     0,     0,    -1,     1,    -1,    -1,    -1,    -1,    -3,     0,     0,    -4,    -4,    -7,    -6,    -8,    -7,    -8,    -7,    -5,    -5,    -5,    -5,    -5,    -7,    -5,    -3,    -5,     1,     0,     0,    -2,    -1,    -6,    -2,    -4,    -1,     0,    -3,     0,    -2,   -11,    -8,    -7,    -6,    -7,    -7,    -6,    -6,    -6,    -6,    -5,    -5,     1,     2,     2,     0,     0,     0,     0,     0,    -2,    -1,     0,    -1,    -4,    -6,    -6,    -4,    -6,    -6,    -4,    -5,    -5,    -4,    -3,    -5,    -5,    -4,    -1,    -1,     0,     1,     1,     0,     0,     0,    -1,     0,     0,    -2,    -3,    -3,    -5,    -6,    -4,    -1,    -2,    -2,    -3,    -1,    -2,    -2,    -1,    -4,    -2,    -1,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,    -1,     0,     1,     1,     0,     0),
		    73 => (    1,     0,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -5,    -5,    -5,    -1,    -1,     0,    -1,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     1,     0,    -1,    -3,    -2,    -3,    -4,    -4,    -4,    -2,    -1,    -1,    -1,    -1,    -2,    -3,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,    -4,    -3,    -6,     1,     2,    -1,    -1,     2,     1,     0,     0,     0,     0,    -1,     2,     4,    -3,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -5,    -5,    -2,     2,     2,    -2,    -1,    -1,     0,    -2,    -1,    -2,     0,    -2,    -1,    -2,    -2,    -6,    -2,     0,     0,     0,     1,     1,     0,    -2,     1,    -1,    -1,     1,     3,     1,     0,     1,    -1,     1,     1,    -2,    -1,    -3,     0,     0,    -2,     0,    -1,    -3,    -4,    -1,     1,     1,     0,     0,     1,    -6,    -5,    -2,     1,     0,     0,    -3,     1,     4,     0,    -2,    -2,    -1,     0,    -1,    -1,    -2,    -1,    -3,    -4,    -3,    -3,     0,     0,     0,     0,    -1,     0,    -4,    -3,     0,     1,     1,    -1,    -1,     2,     2,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,     0,    -2,    -7,    -2,    -5,     1,    -1,    -1,     0,    -1,    -2,    -2,    -1,     1,     0,     1,     1,     3,     2,    -1,    -1,    -2,     1,     2,    -1,     0,     1,    -1,     1,     1,    -6,    -2,    -3,    -2,     0,    -1,     0,    -1,    -1,    -2,    -1,    -2,     1,     0,     1,     3,     2,    -3,    -3,    -1,    -2,    -1,    -2,     1,     3,    -2,     1,     0,    -6,    -5,    -4,    -2,     0,    -2,     0,     1,     3,     2,     1,     0,     3,     0,    -3,    -3,   -11,    -4,    -2,    -2,    -2,    -1,    -2,     1,     2,     3,     0,     2,    -5,    -3,    -2,     0,     0,    -1,     5,     1,     4,     2,     0,    -4,    -3,    -5,    -5,    -8,    -6,    -1,     0,    -1,    -1,    -2,    -1,     0,     1,     2,     2,     2,    -3,     1,    -2,     0,     0,    -2,    -2,    -3,    -3,    -3,    -2,    -8,    -8,    -6,    -3,    -2,     0,     3,     3,    -2,     0,     0,    -1,     0,     0,    -1,    -1,     0,    -3,    -2,    -3,    -1,     0,     1,     2,    -1,    -2,    -7,    -6,    -7,    -1,     2,     1,    -1,     0,     2,     0,     1,    -1,     2,     0,    -2,    -3,    -2,    -2,     0,    -2,    -5,    -3,    -1,    -1,     0,     0,    -1,    -3,    -7,    -9,     3,     3,     0,     1,     1,     3,     3,     2,     1,     0,     0,     0,    -1,    -4,    -2,    -4,    -2,    -2,    -3,     3,    -1,     0,     1,     1,    -1,    -1,    -2,    -1,    -1,     2,     2,     2,     3,     2,     2,     2,    -1,     0,    -1,     0,    -2,    -4,    -3,    -3,     0,    -1,    -2,    -1,    -1,     0,     0,     1,     1,    -3,    -3,    -2,    -2,    -1,     1,     4,     1,     4,     3,     1,    -3,    -2,     0,    -1,     0,    -4,    -3,    -2,    -1,    -5,    -2,    -1,     0,    -1,    -1,     0,     1,    -3,    -5,    -6,    -2,    -3,     0,     1,     2,     3,     0,     0,    -1,    -1,    -3,     1,     0,     1,    -2,    -2,    -4,    -5,    -1,    -1,     0,    -1,    -2,     0,     0,    -5,    -4,    -5,    -5,    -6,    -4,    -5,    -2,    -4,    -1,    -3,    -1,     2,     1,     3,     0,    -2,     1,    -2,    -4,    -5,     0,    -2,    -1,     0,    -1,     1,     3,    -1,     0,    -5,    -8,    -8,   -12,   -16,   -12,    -9,    -3,     0,    -2,     0,     2,     3,     2,     1,    -1,    -2,    -6,    -4,    -3,    -1,     1,    -1,    -1,     2,     5,     3,     0,     0,    -3,    -1,    -2,    -3,    -4,    -3,    -2,     0,     1,     0,     0,     2,     0,     1,    -1,    -2,    -4,    -3,    -1,    -1,     1,     0,     0,     1,     3,     5,     5,     4,     2,     2,     1,     3,     1,    -1,     1,     1,     1,     1,     0,    -1,     0,    -2,    -1,    -3,    -2,    -3,    -2,     0,     0,     0,     1,     1,    -1,     4,     4,     3,     3,     1,    -1,     1,     0,     2,     4,     0,     2,    -4,     1,     0,    -2,     2,     0,    -1,    -1,    -3,    -2,     0,     1,     0,     0,     1,     2,     5,    -1,     2,     2,     0,     0,     2,     2,     1,     2,     0,    -1,    -1,     1,    -6,    -2,     1,     2,     2,     2,    -4,    -1,    -2,     0,     0,     0,     1,    -2,     0,     7,     4,     4,     2,     2,     0,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -7,    -1,    -2,    -4,    -2,    -5,    -3,    -2,    -2,     1,     0,     1,     0,    -2,    -4,     0,     0,    -1,    -1,    -3,     0,     0,    -1,     1,     0,    -3,     0,     1,     1,    -2,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,    -1,     0,     0,     0,    -4,    -3,    -3,    -2,    -2,    -2,    -2,     0,     0,    -1,    -3,    -2,     0,    -2,     0,    -1,     0,     0,     0),
		    74 => (    0,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     1,     0,    -2,     0,     0,    -1,     0,    -1,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     1,     1,    -2,    -2,    -1,    -2,    -4,    -2,    -5,    -3,     1,    -7,    -6,    -4,    -1,     0,    -3,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -3,    -4,    -3,    -1,    -4,    -2,    -2,    -6,    -8,    -6,    -1,     1,    -2,    -3,    -3,    -4,    -5,    -5,    -3,    -4,    -4,    -1,    -3,     0,    -1,    -1,     0,    -2,    -5,    -8,    -3,    -3,     0,    -5,    -6,    -4,    -5,    -9,    -3,     1,    -1,    -2,    -3,    -5,    -2,    -1,    -3,    -2,    -4,    -5,    -2,     0,     0,     0,     0,    -1,    -7,    -1,     0,     0,     1,     0,    -4,    -3,    -3,    -1,     2,     2,     1,     1,     2,     3,     0,    -1,     1,     5,     0,    -1,    -1,    -5,    -1,     0,     0,    -2,    -3,     1,     1,     1,     4,     2,     2,     2,    -1,     2,     3,     4,     1,     0,     3,     1,     4,    -1,     2,     2,     4,     4,     2,    -4,     0,     0,     0,    -1,    -1,     3,     2,     1,     4,     4,     4,     2,     1,     1,     4,     5,     6,     4,     1,    -2,     0,     2,     0,     0,     4,     5,     1,     1,    -3,     0,    -3,    -2,     1,     3,     1,     3,     4,     2,     9,     6,     8,     4,     5,     5,     4,     2,     3,     1,     3,     1,    -1,    -1,     0,     2,    -2,     5,    -4,    -3,    -3,     3,     1,     2,     0,     4,     2,     0,     8,     4,     5,     1,    -1,     0,     1,    -2,    -2,    -1,    -1,     1,     1,    -4,    -1,     0,     1,     2,    -4,     0,    -1,     3,    -2,     0,    -2,    -3,    -1,    -1,     0,     1,    -3,    -1,     1,    -1,     1,    -2,     1,    -1,    -1,    -1,    -1,    -4,     0,    -1,    -2,    -2,    -2,     0,    -2,     1,    -1,    -1,    -3,    -5,    -2,    -2,     1,    -1,    -4,     0,    -3,    -3,    -1,    -1,     0,    -3,     0,    -4,    -2,    -1,    -3,    -5,    -2,     0,    -3,     1,    -3,     1,    -2,    -3,    -2,     2,    -4,     1,    -2,    -3,    -1,     0,    -1,    -2,    -1,     0,     2,    -3,    -2,    -7,    -3,    -2,    -4,    -7,    -2,    -3,    -5,     0,     1,     0,    -2,    -4,    -1,     0,    -3,     0,     0,    -2,     1,     4,     2,    -4,     0,     1,     2,    -1,    -2,     0,     2,    -1,    -3,     1,     3,    -2,    -4,     0,    -1,    -4,    -3,    -4,     0,     0,     4,     2,    -2,     1,     4,     5,     0,     1,     1,     0,     2,     2,    -1,     0,    -2,    -2,    -1,     0,     2,    -1,    -1,    -1,     2,    -6,    -4,     0,     0,     0,     6,     3,     2,     3,     2,     1,    -1,    -1,     0,     1,     1,    -1,    -1,    -3,    -3,    -1,    -1,     0,     2,    -3,     0,    -1,     1,     3,     1,     3,     0,     2,     3,     3,     2,     1,     1,     3,     2,     1,     0,     1,     3,    -1,    -1,     0,     0,     3,     2,    -1,     0,    -2,    -3,     0,     0,    -4,     1,    -2,    -2,    -1,    -1,     0,     0,     2,     2,     0,     0,     1,     0,     1,     1,     1,     1,     3,     2,     2,     0,     1,     1,    -2,    -1,     0,     0,    -2,    -3,     0,     0,    -2,     3,     0,    -1,    -3,    -1,     0,    -2,    -1,    -2,     2,    -1,    -1,     1,     0,     2,     1,     4,     1,    -5,    -1,    -2,    -3,    -1,    -1,     0,     0,     2,     1,     0,    -3,    -1,    -3,    -2,     1,    -2,     0,    -2,    -2,    -4,    -1,     3,     5,     3,     2,     4,     2,    -1,    -2,    -3,     0,    -2,    -3,     7,    -2,    -1,    -2,    -3,    -1,    -3,    -4,    -4,     0,     0,     1,     2,     1,    -4,     0,     2,     2,     1,     2,     0,     1,     0,    -1,    -3,     0,    -1,    -2,     2,    -2,    -3,    -4,    -4,    -2,     2,     0,     0,     0,    -1,     0,     1,     2,    -1,     3,     2,     4,     2,     1,    -1,    -4,    -4,    -2,     0,    -1,     0,    -3,     2,     2,    -2,    -2,    -2,     1,     1,     0,     1,    -3,    -1,    -1,     2,     2,     2,    -1,     3,     7,     5,     6,     2,    -1,    -6,    -4,     0,    -1,    -1,    -1,    -3,    -7,    -4,     0,     1,     3,    -1,     4,     0,    -1,     0,    -3,    -2,     3,     3,     0,     5,     6,     7,     4,     3,     0,     0,    -1,    -1,     1,     0,     0,    -5,    -6,   -12,     2,     3,     5,     3,     6,     4,     2,     0,    -1,    -2,     1,     0,     2,     6,     6,     2,    -2,     2,     0,     4,    -1,     0,     0,     0,     0,    -2,    -6,    -1,     5,     5,     1,     4,     1,     4,    -1,     0,     0,    -4,    -2,    -2,     3,     5,     0,    -2,    -1,     0,    -3,     3,    -3,     0,     0,     0,    -2,     0,     5,     7,     2,    -2,    -1,     1,     3,     2,    -2,     1,    -3,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     1,    -1,    -3,    -2,     1,     0,    -1,     0,    -4,     8,     7,     4,    -1,    -3,    -4,    -8,    -2,    -2,    -2,    -1,    -6,    -6,    -4,    -1,     0,    -5,    -9,    -8,    -2,     0,    -1,     1,     0,     0,    -1,     0,     0,    -1,     0,    -3,    -3,    -2,    -2,    -3,    -4,    -3,    -1,    -2,    -1,    -5,    -7,    -6,    -3,    -4,    -2,    -3,     0,     1,     0,     0,     0),
		    75 => (    0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -2,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -4,    -4,    -2,    -2,    -6,    -1,     1,     1,    -1,     2,     3,     0,     0,     1,    -2,     0,     1,     0,     0,     0,    -1,     1,     2,    -3,    -3,    -3,    -2,    -1,    -1,    -2,     0,     1,     2,     2,     2,     0,    -2,    -2,     1,     2,     1,     2,     1,     1,     1,     1,     0,     0,     0,     1,     0,     0,     2,     2,     1,     2,     0,    -3,    -2,     0,     1,     2,     3,     0,     0,    -2,    -1,     0,     1,     2,     1,     2,    -1,    -2,    -1,     0,     0,     0,    -2,     0,     2,     1,     2,     0,    -1,    -2,    -3,    -1,     0,    -1,     0,     0,     0,     3,     2,     0,     2,     2,     2,     1,    -1,    -2,     0,    -1,    -3,    -2,     1,     2,     3,     1,     0,     0,     0,    -2,    -2,    -1,     0,     0,    -1,    -1,     1,     3,     3,     2,     2,     1,     2,     2,     1,     1,     0,     0,     0,    -2,     1,     4,     1,     1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -2,     0,    -1,    -1,     0,     1,    -1,     2,     2,     4,     2,     2,     2,    -1,    -2,    -2,    -3,     1,     0,     0,     0,    -1,     0,     0,     2,     1,     1,     0,    -2,    -2,    -3,     1,     1,    -1,     0,     3,     4,     2,     3,     2,     1,     0,    -1,    -4,    -3,     0,     1,     0,     0,    -1,    -1,     1,     2,     3,     2,    -1,    -1,    -3,    -2,    -1,     0,     1,     3,     4,     4,     3,     1,     2,     1,     0,     0,    -1,    -5,     0,     0,     0,     1,    -1,     0,     0,     3,     4,     0,     2,     0,    -3,    -1,     0,     2,     3,     5,     5,     4,     3,     2,     0,    -2,     0,    -1,     0,    -3,     1,     0,     1,     1,     2,    -1,    -1,     3,     2,     0,     2,    -2,    -2,    -4,     3,     3,     5,     2,     2,     2,     3,     3,     1,    -2,     0,     0,     0,    -3,     1,     2,     2,     2,     3,     2,    -2,     0,     1,     0,     0,    -1,    -3,     0,     2,     3,     2,     0,    -1,     2,     1,     1,     3,    -2,    -1,     0,     0,    -4,     0,     1,     1,     3,     2,     3,     4,     2,     1,    -1,     0,    -3,    -1,    -1,     0,     3,     2,     2,     0,    -2,    -2,     0,     2,    -2,     1,     0,    -1,    -5,     0,     1,     2,     2,     2,     2,     4,     0,     1,     0,     0,    -2,    -1,     1,     3,     3,     2,     2,     1,    -1,    -2,    -2,    -2,     0,     1,    -1,    -1,     0,     1,     2,     0,     1,     2,     3,     4,     0,     0,     0,     2,     0,     0,     1,     2,     3,     2,     1,     1,     0,     0,    -2,    -2,    -3,     0,    -1,    -2,     0,     1,     4,     1,     1,     2,     2,     2,    -2,     0,     1,     0,     1,    -2,     0,     0,     0,     3,     5,     2,     0,    -1,    -3,    -2,    -4,     0,     0,    -2,     1,     2,     4,     3,     3,     3,     3,    -1,    -1,    -2,     0,     2,    -2,     0,    -1,     0,     0,     2,     1,     2,     0,    -1,    -3,    -4,    -5,     0,     0,    -3,     0,     1,     4,     3,     2,     3,     3,     0,    -3,    -4,     1,     1,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     1,     1,    -2,    -5,    -3,     1,    -1,     2,     0,     1,     2,     2,     4,     3,     0,    -1,    -1,    -2,     1,     0,     1,    -1,     0,    -1,     0,     0,     0,     0,     2,     1,    -2,    -6,    -2,     1,     0,     1,     1,     1,     1,     2,     3,     3,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,     0,     2,     2,    -1,     1,     1,     2,    -2,    -1,    -4,     0,     0,     0,     0,     0,     1,     2,     2,     3,     3,     2,     0,     1,     1,     1,     0,    -1,     0,     0,     1,     2,     2,     0,     1,     1,    -3,     0,    -2,    -1,     0,     0,    -3,     0,     1,     1,     2,     1,     3,     2,     1,     3,     1,     0,     0,     0,    -1,    -1,    -1,     0,     1,    -2,    -1,    -1,    -3,     0,     2,     0,     0,     0,     1,     0,    -2,     0,     1,     2,     2,     1,     0,     1,     1,     1,     1,    -1,    -4,    -3,    -1,    -1,    -1,    -3,    -2,    -2,    -1,     1,     2,     0,    -1,     0,    -1,     0,    -2,    -1,     2,     1,     1,     2,     2,     1,     1,    -1,     1,     0,    -2,    -2,    -1,    -2,    -2,    -2,    -1,    -1,     1,    -4,    -1,     0,     0,     0,     0,     2,    -4,    -3,     0,     1,    -1,    -2,     2,     1,     1,     1,     0,     1,     1,     3,     2,     0,     1,     1,     3,     1,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -4,    -4,    -1,     0,    -1,    -1,     2,    -1,     1,     2,     1,     1,     0,    -1,    -1,    -2,    -2,     1,    -2,     0,     0,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,     0),
		    76 => (    0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     1,     1,     2,     1,     1,     1,     1,     1,    -1,    -1,    -1,     0,     0,     0,     3,     1,     1,     1,     0,     0,     0,     0,     0,     0,     1,     1,     3,     1,     0,     2,     3,     0,    -1,     0,     0,     1,    -1,    -1,    -1,     1,     0,     1,     1,     4,     5,     4,     4,     2,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -4,    -4,    -4,    -2,    -2,    -3,     1,     4,     4,     3,     1,     4,     4,     0,    -3,     0,     1,     0,    -1,     0,     1,     1,    -1,    -2,    -2,     0,    -1,    -2,    -3,    -4,    -5,    -4,    -2,    -2,    -2,     0,     0,     3,     0,     3,     1,    -1,     2,     2,    -1,     0,    -1,    -2,     1,     1,    -1,    -1,    -1,     0,    -2,    -3,    -3,    -3,    -2,    -1,    -2,    -1,     0,     0,    -1,     1,     2,     3,     4,     3,     4,     2,    -1,     0,     0,     0,     1,     1,    -1,    -1,    -2,     0,    -2,    -2,    -1,    -2,    -4,    -4,    -3,    -1,    -1,     1,     0,    -1,     1,     3,     4,     2,     2,     4,     0,     0,     0,     0,     2,     1,    -2,     0,     0,     1,    -3,    -3,    -3,    -5,    -3,    -5,    -2,     0,     1,    -1,    -1,     0,    -2,    -1,     1,     2,     1,     4,     0,     0,     0,    -1,     2,     0,    -3,    -1,    -1,     0,    -4,    -4,    -5,    -4,    -4,    -3,     1,     0,     1,     0,     0,    -1,    -1,    -1,    -3,    -2,     3,    -2,     0,    -1,     0,    -2,     3,     0,    -3,     0,     1,    -1,    -3,    -4,    -4,    -4,    -2,     1,     1,     1,     0,     1,    -1,    -1,    -1,    -2,    -3,    -2,    -2,    -1,     0,    -1,     0,    -1,     2,    -1,    -2,    -1,    -1,    -3,    -7,    -5,    -4,    -1,     0,     1,    -1,    -2,    -3,    -4,    -1,    -1,    -2,    -3,    -2,    -2,    -1,    -2,     0,     0,     1,    -2,     1,     0,    -3,    -3,    -3,    -6,    -4,    -4,    -2,     0,     1,     0,    -2,    -5,    -6,    -4,    -4,    -2,    -2,    -2,    -3,     0,    -1,    -1,    -1,     0,    -1,    -2,     1,    -1,    -2,    -3,    -4,    -4,    -4,     0,    -1,     1,     0,    -1,    -2,    -3,    -6,    -4,    -3,    -2,    -1,    -1,     0,    -1,    -2,    -1,     1,     0,     0,    -1,    -1,    -1,    -2,    -2,     0,    -1,    -1,    -1,     1,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -4,    -2,     0,     0,     0,    -2,    -1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     2,    -2,     1,    -1,     1,     0,     0,    -2,     1,     0,    -1,     0,     0,    -3,    -5,    -4,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,     1,     1,    -1,     1,    -1,     1,     2,     0,    -1,    -1,     0,     1,     0,    -2,    -3,    -3,    -4,    -2,    -1,    -1,    -1,    -2,     0,     0,    -1,    -1,     0,    -2,    -1,     0,     1,     0,     0,     0,     1,     1,     0,     1,    -1,    -2,     1,     0,    -2,    -4,    -2,    -1,    -2,     0,    -1,    -1,     0,     0,    -1,    -3,    -1,    -3,    -2,     0,     1,     0,     3,    -1,    -1,    -3,    -2,    -1,    -2,    -3,     2,     2,     0,    -2,    -1,    -1,    -2,    -1,    -1,    -3,     0,     0,     0,     0,     2,    -1,    -2,    -1,     0,     0,     0,    -1,    -2,    -2,     0,     1,     0,     0,     3,     4,     3,     0,    -1,    -2,    -1,     0,    -3,     0,     0,     0,     0,    -1,     1,    -1,    -2,     0,    -2,     1,    -1,    -2,    -1,    -3,     0,     2,     1,     1,     3,     2,     2,     0,    -2,    -2,     0,     0,     0,    -1,     0,     0,    -1,    -2,     2,     0,     2,     1,    -1,     0,     0,    -1,    -1,     0,     3,     1,    -1,    -1,     0,     1,     0,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,    -2,    -1,     1,     0,     0,     0,     2,    -2,     1,     3,     2,     2,     1,     0,     0,    -2,    -2,    -2,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -4,    -1,     2,    -1,     0,     2,     3,     1,    -2,    -3,    -1,    -3,    -2,    -2,    -2,    -1,    -1,    -2,    -1,    -2,     0,     0,    -1,    -1,     0,    -1,    -2,    -1,    -2,     1,     1,     0,     1,     2,     2,     0,    -1,    -1,    -1,    -4,    -3,    -2,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     1,     0,     0,    -2,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,     0,     0,    -2,    -3,    -3,    -2,    -1,     0,     0,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,    -1,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -1),
		    77 => (    0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,    -2,    -3,    -2,     1,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -2,    -2,    -1,    -2,    -1,    -1,     0,    -2,    -2,    -4,    -1,    -2,    -1,    -1,    -2,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,    -2,    -1,    -1,    -4,    -3,    -3,    -4,    -6,    -7,    -5,    -4,    -7,    -5,    -6,    -5,    -3,    -3,    -1,    -5,    -3,    -2,    -1,     0,    -1,    -1,     1,    -1,    -3,     0,     3,     3,     2,     4,     4,     0,     2,     1,     1,    -1,     0,    -1,    -2,     0,    -1,    -3,    -5,    -5,    -4,    -5,    -4,    -1,     0,     0,     0,     0,    -1,    -1,     2,     2,     3,     4,     0,     1,     2,     3,     3,     4,     1,     3,     2,     2,     2,     2,     1,     2,     0,    -1,    -2,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -2,     2,    -1,     1,     0,     2,     4,     4,     1,     2,     1,     3,     0,     1,     2,     0,     0,     0,     1,    -1,    -1,    -1,    -2,     1,     0,    -1,    -1,    -3,    -2,    -2,    -3,    -3,    -3,     0,     0,    -1,     0,     1,     0,     1,    -1,     0,    -2,    -1,    -3,    -3,    -3,    -1,    -2,    -2,     0,     0,    -1,     1,     0,    -2,    -4,    -3,    -6,    -2,    -3,    -2,    -2,    -3,    -1,    -2,     0,    -3,     0,    -1,    -2,    -2,    -2,    -2,    -2,    -1,    -2,     1,     0,    -1,    -2,    -2,     0,    -2,     0,    -2,    -3,    -2,    -3,    -2,    -5,    -6,    -6,    -2,    -1,     1,    -1,    -1,     0,    -4,    -1,    -3,    -2,    -1,    -2,     1,     0,    -1,    -2,     0,    -2,    -2,    -2,    -4,    -5,    -4,    -6,    -4,    -7,    -4,    -3,    -1,     0,    -1,    -2,    -2,    -1,    -1,     2,     2,    -2,    -4,    -2,     2,     0,     0,    -1,     1,     0,    -2,    -3,    -5,    -4,    -6,    -4,    -5,    -4,    -3,    -2,    -1,     0,    -3,    -4,    -1,    -2,     0,     1,    -1,     0,     0,    -1,     2,     0,     0,     1,     0,    -1,    -2,    -1,     0,    -2,     0,    -2,    -1,    -1,     0,     0,     0,     1,    -2,     0,    -1,     2,     2,    -1,    -2,    -2,     0,    -2,    -2,    -1,     0,     0,    -1,     2,     0,     1,     2,     0,     0,     1,     1,     2,     1,     1,     1,     1,     0,     1,     4,     0,     0,     1,    -4,    -3,    -2,    -2,     1,     0,     0,    -1,     0,     2,     2,     2,     2,     2,    -1,     1,     0,    -1,     0,     0,     1,     3,     2,     0,    -1,    -2,     0,    -2,    -5,    -5,    -3,    -1,    -1,     1,     0,    -1,    -1,     0,     0,     0,    -3,     0,     0,     0,    -2,     0,     1,     0,     2,     1,     0,     0,    -1,     0,    -1,    -3,    -4,    -5,    -3,    -2,    -2,     0,     0,    -1,    -1,    -2,    -1,     2,    -2,    -1,     0,    -1,     1,     0,    -1,     1,    -1,    -2,    -2,     0,     0,     2,    -1,     1,    -1,     1,     1,     2,    -3,     0,     0,    -1,    -2,     0,    -2,    -2,    -1,     0,    -3,    -2,     2,     1,    -1,    -1,    -1,    -5,    -3,    -1,     0,    -2,    -2,    -3,    -2,    -1,     2,     3,    -3,     0,     0,     0,    -1,     1,    -2,     0,    -4,    -4,    -1,    -2,     0,    -2,    -1,    -1,    -3,    -7,    -3,     0,    -1,    -5,    -7,    -3,    -4,    -2,     2,    -2,    -1,     0,     1,     1,     0,    -2,    -1,    -1,    -3,    -2,    -1,     0,     1,    -2,    -2,    -1,    -3,    -4,    -2,    -5,    -5,    -2,    -3,    -3,    -2,    -4,    -4,    -1,    -1,     0,     0,     0,     0,    -1,     1,     0,     0,    -1,     0,     0,     0,     2,     1,    -1,    -1,    -2,    -1,    -3,    -2,    -4,    -3,    -1,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,     2,     0,    -1,     1,     1,     0,     0,     0,     0,     1,    -3,     0,     1,     0,    -1,    -4,    -5,    -3,    -1,     0,    -3,    -1,    -1,     0,     0,     0,    -1,    -4,     0,    -3,     0,     0,     0,    -2,    -1,    -1,     0,     2,    -1,    -1,    -3,    -4,    -2,    -2,    -4,    -2,    -2,     0,     0,     0,    -2,     0,     0,     0,    -1,    -3,    -1,    -2,     0,     2,     1,     0,    -3,     0,     1,     2,    -1,     2,    -4,    -4,    -1,    -1,    -4,    -4,    -3,     1,    -1,    -2,    -1,     0,     0,    -1,     1,     1,     1,     1,    -3,     1,     2,    -3,     0,     1,     2,    -1,    -1,    -3,    -5,    -2,    -1,    -2,    -3,    -2,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -2,    -1,    -2,     0,     3,     3,     2,     0,     0,     2,     2,     2,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     1,     0,    -1,     0,     1,     1,     1,     0,     0,     0,     1,     1,     0,     0,     0,     1,     1,     0,     0,     0),
		    78 => (   -1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     1,     0,     1,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,    -1,    -2,    -4,    -3,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -2,    -1,    -3,     2,     1,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -2,     0,    -1,    -1,    -1,     0,     1,     0,    -1,    -2,     0,     0,     0,     0,     0,    -2,    -3,     0,     0,    -1,    -3,    -3,    -4,    -1,    -1,     0,    -3,    -1,     2,     2,    -1,    -1,    -1,    -2,    -2,     0,    -1,     1,    -1,     1,    -1,     0,     0,    -2,    -2,     1,     1,    -2,    -3,    -3,    -2,    -2,    -1,    -1,     0,     0,     0,     1,     1,     0,     0,    -1,    -1,     0,    -1,    -1,    -2,     0,     1,    -2,    -3,    -1,    -2,     0,     1,     0,     0,    -2,    -2,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -3,    -1,     0,    -2,    -1,     1,     0,     0,     1,     1,     0,     0,    -2,     0,     2,     1,     0,     2,    -2,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -1,     0,    -1,    -1,     1,     0,     0,     0,     1,     0,    -1,    -1,     0,     2,     1,    -2,     1,    -1,    -2,    -1,    -1,     0,     0,     1,     0,     0,     0,    -1,    -2,     0,    -1,    -3,     1,    -1,     1,     0,     0,    -2,    -1,    -1,     0,     2,     1,    -2,     1,     0,    -1,     0,     0,    -1,    -2,     0,    -1,    -3,     0,    -1,    -2,     1,    -1,    -3,    -3,     0,     0,    -2,     0,     0,    -1,    -2,    -3,     1,    -2,     1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -1,     2,    -2,     0,     0,    -1,     0,    -1,    -3,    -2,     1,    -1,    -2,    -1,    -1,    -2,    -3,    -1,     1,     0,     0,     1,     1,    -1,    -3,    -2,     1,     0,     0,     3,    -3,     0,     0,    -2,    -1,    -2,    -1,    -2,     0,     0,    -2,    -2,    -1,    -1,    -3,    -3,     2,     1,     1,     1,     1,     0,     0,     1,    -2,    -1,    -1,    -1,    -4,     0,     0,    -2,    -1,    -2,    -2,    -2,     0,    -1,     0,    -3,    -2,    -3,    -4,    -2,     0,    -1,     0,     2,     1,     0,     1,    -1,    -1,    -2,    -2,    -2,     0,     0,     0,     0,    -1,     0,    -1,    -3,    -1,    -1,     0,     0,    -1,     0,    -4,    -1,    -2,    -3,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,    -1,    -6,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -2,    -1,     0,     0,    -2,     0,    -3,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -1,     0,    -5,    -2,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -2,    -1,    -1,    -2,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -3,    -2,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -3,    -3,    -2,    -3,     0,     2,     1,    -1,    -2,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -2,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -2,    -2,    -1,    -2,     0,     1,     1,     0,     1,    -2,     0,    -1,    -1,    -2,     0,    -1,     0,     0,     0,    -1,     0,     0,    -2,    -2,     0,    -1,    -1,    -2,    -3,     0,    -1,    -1,     1,     1,     0,     2,     2,    -1,     0,    -1,    -2,    -1,    -1,     0,     0,     0,    -3,    -2,     0,     0,    -1,     0,     0,    -2,    -1,    -1,    -1,     1,     0,    -1,     0,    -1,    -2,     0,    -1,     1,     0,    -1,    -3,    -2,    -2,    -1,     0,    -1,    -2,     1,    -2,    -1,    -1,     0,    -1,    -2,    -2,    -3,     0,     2,     0,    -2,     0,    -1,    -2,    -3,     0,     2,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -3,     0,    -1,    -1,     0,    -1,     0,    -2,    -1,    -1,    -1,     1,     1,     1,     0,    -1,    -2,    -2,     2,     1,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,    -2,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -1,    -2,     0,     1,     1,     3,     1,     0,     0,     3,     0,    -1,    -3,    -1,    -1,    -1,    -1,    -1,     0,    -3,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -1,    -2,    -1,    -1,    -1,     0,     0,     1,     1,     1,    -3,    -3,    -3,    -2,    -1,     0,    -1,    -2,    -1,    -1,     0,     0,     1,    -2,    -1,     0,     0,    -1,    -2,    -2,    -2,    -2,    -4,    -1,     1,     0,     2,    -3,    -4,    -3,    -2,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     1,    -1,     0,    -1,    -1,    -1,     0,    -2,    -2,    -3,    -2,    -3,    -5,    -2,    -1,     0,     0,    -1,    -3,    -2,    -2,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,    -2,    -2,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0),
		    79 => (    0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -1,    -2,    -2,    -2,    -2,     0,     1,     2,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -1,    -2,    -2,     2,     1,     2,     0,    -2,    -2,    -3,    -4,    -4,    -4,    -2,    -2,     0,     0,    -2,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -4,    -5,    -3,     3,     0,     0,    -1,     1,     4,    -1,    -1,    -1,     2,    -2,    -2,    -1,    -2,    -2,    -2,     0,     0,    -2,    -1,     0,    -1,    -3,     0,    -4,    -2,    -2,    -1,    -2,     1,     1,     2,     1,     1,     1,    -1,    -3,    -4,    -1,    -2,    -1,    -1,    -1,    -1,    -1,     1,     0,    -1,     0,     0,    -4,    -4,    -8,     3,    -5,     1,     3,     2,     1,     1,    -1,    -1,    -4,    -7,    -3,    -2,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -3,    -1,    -1,    -1,    -2,    -5,    -6,     3,    -1,     2,     3,     3,    -2,    -4,    -1,    -3,    -1,    -2,     1,    -1,    -2,    -1,    -2,    -2,    -2,    -4,     0,     0,    -2,    -1,    -1,    -3,    -3,    -7,    -1,     3,     0,     2,     0,    -4,    -3,    -3,     0,    -1,     1,    -3,     1,     0,    -2,     1,    -2,    -1,    -3,    -2,    -1,     0,    -1,     0,     0,    -2,    -1,    -3,     2,     3,     2,    -1,     1,    -2,     1,     5,     3,     0,     2,     3,     2,    -2,    -5,    -2,    -3,    -1,    -2,     0,    -2,    -1,    -1,     0,     0,    -1,    -2,    -1,     0,     2,     1,     0,     0,     3,     3,     4,     2,     3,     4,     1,     0,    -2,    -2,    -3,    -3,    -1,    -2,     0,    -2,     1,     0,    -1,     0,    -1,    -2,    -3,    -2,    -1,    -1,    -1,     1,     0,     2,     0,     0,     1,     1,     0,     1,    -1,    -2,     0,    -5,    -4,    -2,    -2,    -1,     0,    -1,    -1,    -3,    -2,    -2,    -3,    -1,    -1,     1,    -3,    -1,     0,     2,     0,     3,     2,     0,    -5,    -2,    -2,    -3,    -1,    -2,    -2,    -2,    -2,     0,     0,    -1,    -2,    -2,    -1,    -1,    -3,    -1,    -4,    -1,    -3,    -2,     0,     2,    -2,    -1,     1,     1,    -2,    -3,    -2,    -1,     2,    -1,     0,    -2,    -1,    -1,     0,     0,    -1,    -2,     0,    -1,    -1,    -6,    -5,     0,     1,     2,     2,    -1,     0,    -2,     1,     1,    -4,    -3,    -4,     1,     2,    -1,     1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,    -1,    -3,    -7,    -6,    -4,     0,    -1,    -4,    -3,    -2,     0,    -2,    -2,    -6,    -4,    -1,     1,     0,     1,    -2,     0,    -1,     0,     0,    -2,     0,     0,     1,     1,    -2,    -2,    -5,    -6,    -9,    -5,    -3,    -1,    -2,    -1,    -2,    -2,    -5,    -3,    -1,    -2,    -2,     1,    -1,    -1,    -1,     2,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -4,    -8,    -3,    -2,    -1,    -3,    -1,    -1,    -3,    -4,    -6,    -3,    -3,    -4,    -2,     0,    -1,    -1,     1,    -1,     0,     0,    -1,    -3,    -4,     2,    -2,    -3,    -4,    -5,    -2,    -1,    -1,    -2,    -2,    -3,    -1,     0,    -5,     1,     0,    -1,    -1,    -1,    -1,     1,     0,    -1,    -1,    -1,    -1,     1,    -3,     1,     1,    -1,     0,    -2,    -1,    -1,    -2,    -3,    -2,    -2,     0,    -1,    -4,     0,     1,     0,     2,     1,     0,     0,     0,     0,    -2,    -1,     1,     2,    -4,     0,     2,     4,     1,     0,    -1,    -1,    -3,    -3,    -3,    -1,     0,     0,    -1,    -2,     0,     2,     2,     2,    -2,     0,     0,    -1,    -4,    -2,     0,    -1,    -4,    -3,     2,     3,     0,     2,     0,     0,    -1,    -2,     0,    -1,     1,     0,     0,    -2,    -1,     1,     3,    -3,    -1,    -1,     0,     1,     0,    -2,     0,    -2,    -2,    -3,     0,     2,     2,     3,     1,     1,     2,     1,     0,    -1,     1,     0,     1,    -3,     1,     1,     2,    -1,     0,     0,     0,     0,     0,    -3,     0,     0,    -1,     0,     1,     0,     1,     0,    -2,    -2,     0,    -1,     1,     0,    -3,    -3,     2,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     1,    -1,     0,     0,     2,     3,     0,     1,    -2,    -2,    -2,    -2,    -1,     0,     1,     2,    -3,    -4,     2,     0,     2,     2,     0,     0,     0,     0,     0,     1,     0,     1,     1,     0,    -1,     0,    -5,     0,     3,     1,     0,     0,     4,    -1,    -4,    -3,    -2,    -2,     0,     0,    -1,     1,     1,     0,    -1,     0,     0,     1,     1,    -1,    -1,    -1,     0,     1,    -1,    -1,    -1,     2,     0,    -1,     0,     2,     3,    -2,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0),
		    80 => (    0,     1,    -1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,    -1,    -1,     1,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     1,     1,     0,     1,     0,     0,    -1,     0,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     4,     3,     0,     0,     1,    -1,    -1,     0,    -3,    -2,    -4,    -4,    -4,    -2,    -3,    -2,    -3,    -2,    -2,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     1,     5,     3,     1,    -1,    -1,    -2,    -2,    -2,    -1,    -1,     2,     0,    -1,     0,    -1,    -1,     0,     1,    -4,    -3,    -3,     0,    -1,    -2,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -1,    -1,    -2,    -3,    -1,    -1,     1,    -2,     0,     2,     1,     2,     1,     4,    -1,     0,    -2,    -3,     0,     0,     0,    -1,     1,     0,     0,     1,    -4,    -4,    -4,    -4,    -6,    -3,     0,    -1,    -1,    -1,     1,     1,     1,     3,     2,     5,    -1,     0,    -2,    -2,    -1,    -1,     0,    -1,    -1,     1,     3,     0,     0,    -3,    -6,    -5,    -5,    -1,     2,     0,     1,    -3,    -1,     0,     0,    -1,     3,     2,    -2,    -4,    -5,    -3,     0,     0,     0,     0,    -1,     2,     3,     1,    -1,    -2,    -1,    -2,     1,     0,     0,    -2,     0,    -1,    -1,     0,     2,     1,    -2,     2,     1,    -1,    -1,    -4,     1,     1,    -1,     1,    -1,     0,     2,     2,    -2,    -2,    -3,    -4,    -4,    -1,    -1,     2,    -2,     1,    -1,     1,     1,     1,     2,     2,     1,    -3,    -3,    -4,    -1,     0,     0,     2,     0,    -2,     2,    -1,    -2,    -1,    -5,    -2,    -3,    -1,    -1,     2,     1,    -2,     0,     1,     0,     1,    -1,     1,     3,     2,     1,    -3,     0,     0,     0,     1,     0,    -2,    -1,    -4,    -2,    -2,     1,    -2,    -1,     2,     0,     0,     1,     0,    -2,    -4,    -1,     3,     2,     3,     2,     2,     1,    -5,    -1,     0,     2,    -1,    -1,    -3,    -3,    -2,     2,     1,    -1,    -1,     0,     0,    -2,    -1,    -2,    -5,    -6,    -5,     0,     1,     1,     0,     0,    -1,     0,    -3,     0,     1,     2,    -1,    -1,    -1,    -2,    -2,     0,     0,    -1,     2,     2,     2,     2,     1,    -1,    -8,    -8,    -2,     1,    -2,    -1,     1,     4,     0,    -1,    -2,     0,     1,     1,     1,    -2,    -2,    -1,     0,     1,     1,     1,     0,     2,     1,     1,     0,    -2,   -10,    -4,     2,     0,    -2,    -3,     0,     8,     2,     2,    -2,    -1,     0,     0,     0,    -5,    -1,    -1,     1,     3,     0,     1,    -2,     0,    -1,    -1,    -8,    -7,    -7,    -3,    -2,    -1,    -1,     1,     1,     3,     1,    -1,    -4,     0,     0,     0,    -1,    -6,     1,    -2,     0,     3,     1,     1,    -3,    -1,     2,     0,    -6,    -4,    -1,     0,    -2,    -1,    -4,     1,     1,     2,     4,    -2,    -4,    -1,     1,     0,     0,    -4,     1,     0,     0,     3,     2,    -2,    -2,     0,    -2,    -4,    -2,     0,     0,    -1,     1,    -2,    -1,    -2,    -1,     0,     2,    -3,    -2,     0,     0,    -1,    -2,    -2,     1,     2,     1,     3,    -1,     1,     0,    -2,    -5,    -4,    -2,    -1,    -2,     0,     0,     1,     1,    -3,    -2,     1,     2,    -4,    -2,     0,    -1,     0,    -1,     0,     1,     0,     1,     2,     3,     2,    -3,    -5,    -4,    -2,     0,     0,    -1,     0,     1,    -2,     0,    -1,     1,     1,     0,    -2,    -1,    -1,     1,     1,    -3,    -1,     4,     0,     0,     2,     1,     2,    -3,    -5,    -2,    -3,     0,     1,    -2,     1,    -2,    -1,    -3,    -1,     1,     0,     1,    -2,     0,     0,     0,     1,    -5,     1,     3,     1,     2,     0,     1,     1,    -1,     1,    -1,    -1,    -1,    -3,    -1,    -1,    -1,    -3,    -4,    -1,     0,     0,     0,    -2,     1,     1,     0,     1,    -5,     1,     1,     1,     2,     3,     1,     1,     0,     0,    -2,    -1,     0,     1,     0,     0,    -2,    -3,    -4,    -5,    -3,    -1,     2,    -1,     1,     1,     0,     0,    -5,     0,     0,     2,     3,     1,     1,     1,     1,    -1,    -2,     0,     2,     0,    -4,    -3,    -2,    -2,    -5,    -3,    -1,     0,     2,     0,     0,     1,     0,     0,    -1,    -4,    -4,     1,     0,     0,     1,     2,     2,     2,     0,     1,     1,    -3,    -4,    -3,    -4,    -3,    -5,    -2,     1,     0,    -3,     0,     0,     0,     0,     0,    -1,    -1,     4,     5,     0,    -1,     0,     2,     4,     3,     4,    -4,    -3,    -4,    -7,    -6,    -3,    -4,    -2,     0,    -1,     0,     2,     0,     0,    -1,     0,    -1,     0,     0,    -2,    -5,    -4,    -4,    -4,    -2,    -3,    -4,    -5,    -4,    -2,    -4,    -4,    -4,    -5,    -4,     0,    -1,    -1,    -1,     0,     0,    -1,     0,     1,     0,     0,    -1,    -1,    -3,    -5,    -1,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -3,    -3,    -4,    -5,    -1,    -3,    -1,    -1,    -1,     0,     0,    -1,     0,    -1,    -1,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0),
		    81 => (   -1,     0,     1,     1,     0,     0,     0,    -1,    -1,     0,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,    -1,     1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     3,     4,     8,     6,     3,    -2,     0,    -3,    -2,    -2,     0,     0,     0,     0,     0,     0,     1,     1,    -1,    -2,    -4,    -1,     3,     1,    -2,    -3,    -3,    -1,     1,     5,     5,     1,     0,    -2,     0,     3,    -1,     0,    -2,     0,     0,     0,     0,     1,     2,     1,     3,     1,    -1,    -1,     4,     3,     2,     0,     0,    -2,     0,     1,     1,     1,    -1,    -1,     2,     3,     1,     2,     0,    -2,    -1,    -2,     0,    -1,     0,     0,     3,     7,     3,     2,     2,     1,     0,    -3,    -3,     1,     2,     1,    -1,     1,     0,     1,     2,     2,     2,     1,     0,    -1,    -2,    -2,     0,     0,    -4,     0,     1,     1,     3,     1,    -2,    -2,     1,    -1,     0,    -1,     0,    -1,    -2,     2,     1,     3,     2,    -1,     1,     0,     0,     0,    -1,     0,    -1,     0,    -5,    -4,    -4,     0,     2,     2,    -3,     1,     2,    -2,     0,    -3,    -1,     2,    -1,     1,     2,     3,     1,     0,     1,    -1,    -1,     0,    -2,    -1,     0,     0,    -5,    -3,    -4,    -1,     1,     0,    -1,     1,     1,     1,     1,    -3,    -3,     1,     2,     0,     2,    -3,    -2,    -1,     1,    -2,     0,     0,    -2,     0,     0,     0,    -5,    -2,    -3,    -3,     0,     1,     2,     0,     0,     4,     3,    -2,    -3,    -1,    -2,    -2,    -2,    -1,    -1,    -1,    -2,     0,    -1,     0,     0,    -1,     0,     0,    -4,    -1,    -5,    -2,    -4,     0,     2,     3,     1,     4,     1,    -1,    -2,    -1,    -3,    -2,    -1,    -4,    -2,    -3,     0,     0,    -1,    -1,     1,     0,     0,     1,    -1,     0,    -4,    -2,    -4,     0,    -2,     1,     0,     2,     1,    -1,     0,    -3,     0,    -3,    -3,    -3,    -2,    -2,     0,     0,    -1,     0,     0,     1,     0,     0,    -1,    -1,    -3,    -3,     1,     2,     1,     0,    -1,     0,     0,    -2,    -3,    -1,    -1,    -3,    -1,    -3,    -5,    -2,    -1,    -1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -3,     1,     2,     2,     3,    -1,    -2,     0,    -1,    -3,    -1,     2,    -1,    -2,    -2,    -7,    -3,    -3,    -2,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -3,     3,     2,    -1,    -1,    -4,    -5,    -3,    -2,    -2,     1,     1,     0,    -2,    -3,    -5,    -4,    -5,    -3,    -2,    -1,    -2,     0,     0,    -1,     0,     0,     1,    -1,    -2,    -1,    -1,    -3,    -4,    -5,    -5,    -5,     0,     2,     0,    -1,    -2,    -3,    -6,    -4,    -4,    -3,    -3,    -7,    -1,     0,    -1,     0,     0,     1,    -2,    -1,    -1,    -2,    -2,    -5,    -3,    -3,    -5,    -4,     0,     3,     2,    -1,    -3,    -2,    -5,    -4,    -5,    -2,    -4,    -2,    -1,    -1,    -1,     0,     0,     0,    -3,    -1,    -1,    -2,    -4,    -4,    -4,    -4,    -9,    -5,    -4,     1,    -1,    -1,    -2,     0,    -2,    -3,    -2,     0,    -2,    -4,    -4,     0,    -1,    -1,     0,     0,    -1,    -1,    -3,    -6,    -4,    -6,    -4,    -4,   -11,   -10,    -5,     0,    -2,    -1,     1,    -1,    -1,     2,     1,     3,    -1,    -7,    -2,    -2,    -1,     0,     0,    -1,    -1,    -2,    -6,    -3,    -1,     0,    -2,    -3,    -5,    -3,    -3,    -2,     1,     3,     0,    -2,     0,     1,     0,     0,     1,     0,     0,    -2,    -1,     0,    -1,    -2,     2,     0,    -4,    -2,     1,     1,     2,     4,     0,    -1,     0,     1,     1,     3,     2,     5,     4,     3,     0,     1,     1,     1,     0,    -2,     0,     1,     1,    -2,     2,     3,     1,     3,     3,     3,     3,     2,     2,     0,     1,     1,     3,     1,     3,     5,     1,     2,     0,    -2,    -1,     1,     2,    -2,     0,     1,     0,    -6,    -4,     2,     4,     1,     0,     1,     1,     1,     1,     1,     1,     0,     1,    -1,     1,     1,     3,     3,     1,    -5,    -3,     1,     0,     0,     0,     1,     0,    -1,    -2,     1,    -1,     1,    -1,     0,    -1,    -2,     0,     0,     2,    -2,    -3,    -5,    -4,    -1,     1,     2,     3,    -1,    -3,    -3,    -3,     2,     0,     0,     0,     0,     0,    -1,    -2,    -2,     0,     1,     1,    -1,     0,    -4,    -3,    -6,    -5,    -4,    -3,    -2,    -1,     1,     1,    -1,    -2,    -3,     0,     0,     1,     0,     0,     1,    -1,     0,     0,    -1,     0,     0,    -3,    -1,    -2,    -2,    -3,    -2,    -4,    -3,    -3,    -4,    -3,    -4,    -3,    -3,    -1,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -3,     0,     0,    -1,    -2,    -1,    -3,    -1,    -3,    -2,    -2,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1),
		    82 => (    0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,    -1,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     1,     0,    -1,    -2,    -1,    -2,    -2,    -2,    -4,    -2,     0,     2,     0,    -2,    -5,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     0,     1,     0,    -3,    -3,     1,     0,    -1,     0,     4,     3,     2,     1,     1,     0,     2,     0,     0,    -2,    -3,    -2,    -1,    -1,     0,     1,     1,     0,     0,     0,     0,     0,    -4,    -5,    -1,     0,     1,    -1,     2,     1,     1,    -1,     1,     3,     1,     1,     0,    -2,    -2,    -1,     1,    -2,    -6,     1,     1,     0,     0,     0,     0,    -1,     1,     1,    -2,     0,    -1,    -3,     1,     3,     0,     0,     2,     2,     1,     1,     1,     3,     0,     0,    -1,    -3,    -1,    -2,    -1,    -1,     0,     0,    -1,     1,     0,     0,     1,     1,    -3,     0,     1,    -2,    -1,     1,     0,     0,    -1,     2,    -1,     1,    -1,    -1,    -1,    -2,    -1,    -4,     0,    -2,    -1,     0,     0,     0,    -1,    -2,     0,     0,     2,    -2,    -2,     1,    -1,    -3,     2,     0,     1,     3,     0,     1,    -2,    -1,     0,    -1,    -2,    -5,     2,    -1,    -1,     0,     0,     0,    -1,    -2,    -1,     1,     0,    -2,    -2,     2,     0,     0,    -2,     0,     1,     0,     0,    -3,    -1,     1,     2,     0,    -5,    -2,     1,    -2,    -1,    -1,     1,    -1,    -2,    -1,    -3,    -2,     0,     1,     1,     2,     1,    -3,    -2,    -3,     0,     0,     1,     1,     2,     0,     0,     0,    -2,    -4,    -5,    -2,    -1,     0,    -1,    -1,    -2,    -1,    -4,    -4,    -4,    -5,    -1,     0,    -3,    -4,     0,    -1,    -3,    -1,     1,     2,    -2,    -1,     3,     0,    -2,    -2,    -3,    -2,    -1,    -1,     0,    -1,    -3,    -3,    -4,    -4,    -9,   -12,   -11,    -9,    -7,    -2,    -3,    -1,    -3,     0,    -1,     1,     0,     0,    -1,     0,    -1,    -4,    -3,    -1,    -1,     0,    -2,    -2,    -3,    -3,    -4,    -6,    -7,   -10,    -8,    -7,    -4,    -3,    -4,    -1,    -3,    -2,    -4,    -4,     0,     0,     0,     1,    -1,    -4,     0,    -1,    -1,     1,    -2,    -4,    -3,    -5,    -4,    -4,    -5,    -1,    -1,    -1,     1,    -1,    -1,     1,    -2,    -3,    -4,    -3,    -1,    -1,     1,     3,    -3,    -3,     4,     0,    -1,    -1,    -2,     0,    -1,    -3,    -2,     1,     5,     2,    -1,    -1,     1,     4,     3,     1,     1,     0,     0,    -2,    -2,     0,     2,     4,     0,    -1,     2,     0,     0,     0,    -2,    -3,     3,     2,     0,     3,     5,     4,     3,     4,     3,     3,     4,     4,     0,     2,    -3,    -2,    -1,     1,     0,     1,     1,    -1,     2,     2,     2,     0,    -1,     1,     7,     3,     4,     2,     2,     2,     2,     3,     1,     2,     1,    -2,     1,    -1,     1,    -1,     0,    -2,    -1,    -1,     2,     0,     3,     6,     3,     0,     0,     1,     3,    -1,     4,     6,     3,     1,     2,     2,     0,    -2,     1,     1,     1,     1,     1,     0,     0,    -2,    -2,    -1,    -1,    -2,     4,     6,     2,     0,    -1,     0,    -2,     2,     1,     4,    -1,     2,    -1,    -2,     1,     0,    -1,     3,     2,     2,     0,     0,    -2,     0,    -4,    -3,    -4,    -5,     1,     1,     4,     0,     0,    -2,     1,     0,     3,     3,     0,     0,    -1,    -2,    -1,     0,     1,    -1,     0,     2,     1,     2,     3,     1,    -1,    -2,    -2,     1,     3,     2,     3,     0,    -2,    -2,    -1,     2,     2,     2,     2,     1,     1,    -2,     0,     0,    -1,    -2,     0,     1,     0,     2,     3,     0,     2,     2,     1,     3,     3,     3,     2,     0,    -2,     0,     0,     1,     4,     1,     0,    -1,    -2,    -1,    -3,    -3,    -3,    -3,    -1,     0,    -2,    -2,     0,    -1,     0,    -1,     1,     4,    -1,     1,     0,    -1,     2,     0,     1,     2,     1,     1,     1,     2,    -2,    -2,    -1,    -1,    -3,    -2,    -2,    -2,    -1,    -2,     0,     1,     2,     1,     2,     1,    -2,    -1,     0,    -1,     0,     0,     1,     2,    -2,    -2,    -1,    -1,    -2,    -1,     0,    -1,    -3,    -4,    -1,    -2,    -3,    -3,    -1,     0,     1,    -1,    -1,    -1,    -4,    -4,     0,     0,    -1,     1,     3,     3,     0,    -3,    -1,    -2,    -4,    -1,    -2,     0,    -5,    -3,    -4,    -2,    -2,    -3,    -5,    -2,     0,     2,    -3,    -3,    -2,    -3,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -2,    -3,    -5,    -6,    -4,    -3,    -6,    -4,    -4,    -4,    -2,    -2,    -5,    -6,    -3,    -5,    -3,     1,     2,     2,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -4,    -2,    -1,    -1,    -4,    -3,    -2,    -3,    -4,    -2,    -5,    -4,    -2,    -3,    -1,    -1,     1,     2,     0,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -1,     0,     0,     0,     0,    -2,    -1,    -4,    -3,    -2,    -2,    -1,    -1,    -1,    -1,     1,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     0),
		    83 => (    1,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     1,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -3,    -2,    -2,    -1,    -3,    -1,    -2,    -1,    -1,    -1,     0,     1,     0,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -3,    -4,     2,     0,    -1,    -2,    -3,    -3,    -2,     0,     0,    -3,    -4,    -5,    -4,    -4,    -1,     1,     0,     0,     0,     0,    -1,    -1,    -1,     1,     3,     7,     7,     3,     3,     3,     2,     1,    -1,     3,     4,     3,     3,     6,    10,     1,    -6,    -7,    -3,    -2,     0,     0,     1,     0,    -4,     0,     1,     2,     1,     4,     5,     0,     3,     1,     2,    -1,     1,     0,     2,     3,     2,     3,     1,    -3,    -4,   -13,   -10,    -4,    -3,     0,     0,     1,    -1,     0,     0,     2,     5,     6,     1,     1,     2,    -1,    -2,     0,    -1,     0,     3,    -2,    -1,     2,     0,    -1,    -1,     1,     1,    -5,    -2,     0,     0,     1,     1,     0,    -1,     4,     7,     5,     3,     3,     1,     0,    -2,     1,     0,     2,     2,     1,     1,     0,     0,    -1,     0,     1,     2,    -6,    -3,    -1,     0,     0,     0,     1,    -1,     1,     6,     8,     4,     0,     1,     4,     1,    -2,     1,     0,     2,    -1,    -2,     1,    -1,    -1,    -2,    -1,     2,    -5,    -3,    -1,    -2,    -1,    -2,     0,     1,     4,     1,     2,     1,    -1,    -1,    -3,    -3,    -2,    -1,     3,     2,     2,    -3,     2,     0,    -2,     2,     0,    -2,    -3,    -3,     0,     0,    -1,    -6,    -1,     6,     6,     3,     3,     3,    -1,     1,    -2,    -2,    -1,    -2,    -1,     0,     3,     2,    -1,     1,    -1,     4,     3,    -7,    -3,    -2,     0,    -1,     0,    -7,     0,     1,     3,     4,     5,     0,    -1,    -3,    -4,    -2,    -3,    -1,    -2,     0,     2,     3,     1,    -3,    -2,     1,     5,    -3,    -3,    -3,     0,    -1,    -2,    -3,     3,     5,     5,     3,     1,     2,    -1,    -1,    -3,    -3,    -1,     0,    -3,     0,     1,     1,    -2,    -3,    -2,     0,    -1,    -8,    -6,    -3,    -1,    -1,    -1,    -3,     1,     4,     5,     4,     2,     1,    -2,     1,    -1,    -2,    -2,    -2,     0,     1,     0,     1,     1,    -2,    -4,    -2,     0,    -5,    -4,    -1,     0,     1,    -1,    -3,     0,     5,     4,     2,     2,     4,     0,     2,    -1,    -2,    -1,    -1,     2,    -6,    -2,     3,     2,    -2,    -2,    -3,     2,    -1,    -6,    -1,    -1,     0,     1,    -1,     1,     2,     4,     4,     0,     2,     0,    -1,    -1,     0,    -2,     1,    -3,    -3,    -1,     2,     2,     1,     1,    -1,     2,    -1,    -8,    -4,     0,    -1,     2,    -1,     1,     2,     5,     3,    -3,    -2,    -3,     0,    -2,    -1,    -2,    -2,    -1,    -3,    -3,    -1,     3,     0,     1,     2,     4,     4,    -8,     1,    -2,     0,     0,     1,     5,     5,     4,     1,     2,    -4,     0,     0,    -3,    -5,    -1,     0,    -1,    -3,    -2,     3,     4,     1,    -2,     2,     0,     3,    -9,    -4,    -2,     0,     1,    -1,     3,     3,     1,    -1,     1,    -1,    -1,    -2,    -2,     0,     0,    -3,    -2,     1,     1,     2,     4,    -1,     0,    -2,    -1,    -2,    -8,    -2,    -1,    -1,     1,     0,     2,     4,     3,     0,     0,    -1,    -3,     0,    -1,    -2,     2,     0,     2,     0,     2,     4,    -2,     1,    -2,    -1,    -5,    -1,    -7,     0,    -2,     0,    -1,     1,     1,     2,     3,    -1,    -2,    -3,    -5,    -2,    -3,    -1,     1,     3,     2,     0,     2,     2,    -1,     1,    -1,    -1,    -2,     1,    -4,    -3,    -2,     0,     1,    -3,     1,     2,     2,     0,    -1,    -3,     0,    -2,    -2,    -1,     0,     2,     2,     5,     3,    -1,    -1,     2,     2,     2,     2,     0,    -5,    -2,     0,    -1,    -1,     1,     0,     1,    -3,     2,     3,     0,    -1,    -2,     0,     1,     2,     4,     4,     3,     1,     2,     3,     0,     2,     3,    -1,    -4,    -5,    -3,     0,    -1,     0,     3,     2,    -3,     2,     3,     4,    -1,     1,     2,     1,    -1,     1,     2,     1,    -2,     1,    -1,     3,     0,     2,     5,     1,    -3,    -4,    -2,    -1,     0,     0,     1,     0,    -2,    -1,     2,     4,     1,     1,     1,     2,     0,    -1,    -1,     2,     1,     0,    -1,    -2,     0,     5,     5,     2,     5,     2,    -3,     1,     0,     0,     3,     5,     4,     0,     3,     3,     2,     4,     1,    -1,    -1,     0,     1,    -1,     0,     0,    -2,     1,     7,     4,     2,     3,    -5,    -3,    -1,     0,     1,     0,     1,    -1,     0,     4,     3,    -1,     1,     2,    -2,    -1,     1,     4,     0,    -1,    -1,     1,     2,     2,    -2,    -5,    -6,    -6,    -5,    -1,    -1,    -1,     0,     0,     0,    -1,    -6,     3,     1,     0,     2,    -1,    -1,    -3,    -3,    -2,    -2,     0,     5,     6,     5,     1,    -1,    -2,    -7,    -3,     0,     0,     0,     1,     0,     0,     0,     0,    -1,    -2,    -2,    -1,    -1,    -4,    -3,    -3,    -2,    -4,    -3,    -2,     0,    -1,     0,    -3,    -4,    -1,    -1,    -1,     1,     0,     0,     0),
		    84 => (    0,     0,     1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -2,    -3,    -2,    -2,    -3,    -3,    -1,    -3,    -3,     0,    -2,    -1,    -3,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -4,    -3,    -4,    -6,    -5,    -7,    -7,     1,     2,     0,    -4,    -3,    -4,    -6,    -4,    -7,    -3,    -3,    -2,    -1,    -2,     1,     0,     0,     0,     0,    -7,    -4,    -5,    -3,    -4,    -3,    -6,    -5,    -6,    -3,    -7,    -1,    -1,    -4,    -2,    -2,     0,     3,     0,    -3,    -4,    -2,    -1,    -1,     0,     0,     1,    -3,    -6,    -1,     0,     1,     0,    -3,     0,    -1,    -4,     0,    -1,    -2,    -3,    -1,     0,    -1,     0,     0,    -2,     1,     1,     2,    -1,    -4,    -1,    -1,    -1,    -3,     0,     0,    -1,     0,    -1,     2,    -1,     2,     0,     3,    -2,    -1,    -3,    -2,     2,    -1,     0,    -3,    -1,     0,     0,    -2,     2,    -2,     0,     0,     0,    -2,    -3,     1,     3,     2,    -3,    -1,    -3,     0,     1,     0,    -2,    -5,    -5,    -4,    -3,    -4,    -2,    -5,     0,     0,     0,    -1,    -1,     0,    -2,     1,    -6,    -2,     0,     1,     2,    -3,    -3,    -5,    -2,    -1,     0,    -3,    -3,    -4,    -5,    -4,    -1,    -2,    -3,    -3,    -2,    -2,    -2,     1,     3,     3,    -4,    -2,    -5,     3,     1,     3,     1,    -4,    -5,    -5,    -2,    -4,    -3,    -2,    -1,    -6,    -4,    -3,    -1,    -1,    -1,    -2,    -3,    -2,    -1,     2,     3,     0,    -1,     0,    -4,     3,     1,    -2,     0,    -3,    -2,    -3,    -3,    -4,    -1,     0,    -2,    -4,    -1,    -2,    -1,     0,     2,     1,     3,     2,     2,     3,    -2,    -4,    -1,     1,    -3,     2,     1,    -2,     2,    -1,    -3,    -1,     0,     0,     0,     2,    -1,    -2,     2,     2,     4,    -1,     0,     2,     1,     1,     0,     0,     1,    -2,    -1,     0,    -3,     0,     0,     0,     4,     0,     0,     1,     4,     3,     2,     4,    -1,     0,     3,     4,     1,    -2,    -1,     0,     1,     2,     2,    -1,    -1,    -4,    -4,     0,     0,     2,     2,    -1,     3,     2,     2,     2,     3,     3,     3,     3,     1,    -1,     0,     0,    -1,    -2,     0,    -1,     2,     3,     2,     4,     2,     2,    -4,     0,    -1,     0,     4,     2,     3,     1,     2,     0,     2,     2,     5,     4,     2,     0,    -1,     2,     1,    -2,     0,     1,     3,     2,     3,     2,     6,     5,    -3,     0,     1,    -6,     2,     5,     4,     2,     2,     3,     2,     2,     1,     3,     0,    -1,    -2,     2,     4,    -2,     3,    -1,     4,     2,    -2,     0,     3,     3,    -1,     0,     1,     6,     3,     0,     3,     1,    -1,     1,     1,     2,     1,     1,     1,    -1,     2,     3,     1,     0,     3,     0,     0,     3,     2,    -1,     2,     6,    -1,     0,     0,    -1,     4,     1,     3,     3,     3,     2,     1,     0,    -1,     1,     0,    -1,     4,     1,     2,     4,     5,     1,     1,     0,     0,     0,     2,     4,    -1,     0,    -1,     2,    -1,     4,     3,     1,     2,     0,     1,     0,     0,     0,     1,     1,     1,     2,     1,     0,     2,    -2,     0,     1,     1,     1,     1,     3,     0,    -3,     0,     3,     1,     3,     0,    -1,    -1,     1,     2,     0,     2,     1,     3,     3,     0,     0,     1,     1,    -1,    -1,     0,    -1,    -2,    -1,    -4,    -1,    -1,     0,    -2,    -2,     5,     0,     4,     1,    -3,     1,     0,    -2,     0,     0,    -1,     2,     0,    -1,    -2,    -2,    -4,    -3,    -2,    -4,    -4,    -1,    -3,    -1,    -1,     0,    -1,    -3,     3,     2,     0,     0,     0,     1,    -3,    -6,    -3,    -4,    -2,    -1,    -3,    -1,    -3,    -4,    -3,    -6,    -4,    -3,    -4,    -1,    -6,    -1,     0,     0,    -1,    -5,     1,     2,     1,    -3,    -5,    -1,    -3,    -4,    -2,    -3,    -3,    -4,    -2,     0,    -2,    -3,    -4,    -1,    -3,    -2,    -3,     1,    -4,    -4,     0,    -1,     0,     0,    -4,    -6,    -1,     0,    -5,    -5,    -4,    -1,    -1,    -3,    -3,    -2,    -1,    -2,    -3,    -2,    -1,    -3,     1,     0,     2,    -2,    -1,    -1,    -1,     0,     0,     0,    -5,    -2,    -6,     0,     2,     0,    -3,     2,    -2,    -1,    -1,    -2,    -1,    -2,     0,    -2,    -1,    -2,     1,    -1,    -3,    -4,     0,     0,     1,     0,     0,     0,    -1,    -5,     0,     1,     2,     2,     1,    -2,    -1,    -4,     1,     2,    -2,     0,    -2,    -5,    -3,    -1,     1,    -1,    -2,    -7,    -1,    -2,     0,     0,     0,    -1,    -1,     1,    -3,     1,     0,    -1,    -3,    -1,    -1,    -4,    -4,    -2,    -5,    -1,    -2,    -2,    -4,    -1,     0,     2,    -1,    -4,    -2,    -1,     0,     0,     0,     0,    -4,    -2,    -1,    -4,    -4,    -2,    -2,    -6,    -4,    -3,    -7,    -6,    -4,    -6,    -2,    -1,    -6,    -8,    -8,    -7,    -2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -5,    -5,    -3,    -4,    -5,    -2,    -3,    -6,    -3,    -4,    -5,    -4,    -3,    -1,     0,     0,     0,    -1),
		    85 => (    0,     0,     1,    -1,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,    -1,     0,    -1,     1,     0,     0,    -1,    -2,    -2,    -3,    -2,    -2,    -3,    -2,    -3,    -4,    -2,    -2,    -1,     0,    -1,     0,     0,     0,     0,     1,    -1,    -1,    -1,    -1,    -2,    -1,    -6,    -5,    -7,    -6,    -5,    -5,    -5,    -1,    -1,     1,     1,    -1,     1,     1,    -1,     1,    -2,    -1,     0,     0,     0,     0,    -2,     2,     3,    -2,    -7,    -5,    -1,     1,     2,    -3,    -4,    -1,    -2,     4,     3,     1,     5,     4,     4,     8,     6,     5,    -2,     2,     1,     0,     0,     0,    -2,     2,    -7,    -6,    -3,    -2,    -7,    -2,     2,    -2,    -2,    -3,     1,     3,     3,     5,     9,     4,     5,     6,    10,     4,    -3,     1,    -2,    -2,     0,     0,    -3,     3,    -7,    -2,    -2,    -2,     0,     2,     3,     0,    -2,    -3,     1,     1,     3,     4,     5,     6,     7,     1,     4,     1,    -2,    -2,    -3,    -4,     0,     0,    -1,    -7,    -1,     4,     4,     2,     3,     1,     1,     0,     0,    -3,     0,     0,     1,     0,     4,     6,     4,     0,     3,     3,     5,     5,     1,     1,     0,    -1,    -1,    -8,    -4,    -2,     2,     1,     0,     0,     0,     3,    -2,    -1,    -1,    -5,    -1,    -2,     3,     5,     2,     2,     7,     6,     6,     1,     3,     4,    -2,    -2,    -3,    -8,    -3,    -3,     1,     2,    -1,     0,    -3,     1,     2,     0,    -2,    -4,    -5,    -1,    -2,     5,     3,     3,     6,     5,     4,     1,     2,     3,     0,     0,    -3,    -4,    -2,    -2,    -1,     1,     1,    -2,     1,     0,     0,     0,    -3,    -5,    -5,    -4,    -1,     4,     0,     1,     3,     4,     4,     2,     0,     0,     0,    -1,    -2,    -7,     1,     0,    -3,    -3,     0,     2,    -3,     2,     2,    -2,    -3,    -2,    -6,    -4,     1,     1,     1,     3,     3,     5,     6,     1,    -2,    -2,     0,    -1,     0,    -5,     1,    -2,     0,    -2,     1,    -1,    -1,     0,     1,    -2,    -4,    -2,     2,     1,     0,     1,    -3,    -1,     2,     4,     5,     4,    -2,    -1,     0,     0,    -1,    -4,     4,    -1,    -1,     2,     2,     2,     5,     0,     4,    -1,    -1,    -3,    -1,    -1,    -1,    -3,    -3,    -2,     0,     1,     1,     4,     6,    -2,     1,     0,     0,    -4,     0,     1,    -1,     3,     0,     0,     2,     2,     3,    -1,    -2,    -1,    -1,    -2,    -4,     1,    -1,     2,    -3,    -4,    -4,    -3,     4,    -2,     0,     0,    -1,    -5,     3,     1,     4,    -1,     0,     2,     2,     2,    -1,     0,     1,     0,     0,    -2,     1,     0,     2,    -1,     2,     0,    -1,    -5,    -5,    -2,     1,     0,    -3,    -1,     3,     5,     0,     2,    -1,     1,     2,    -1,    -1,     0,    -1,    -5,    -2,     1,    -1,    -1,    -1,    -1,     0,     1,     1,    -2,    -4,    -1,     0,    -1,    -3,    -1,     1,     4,     5,     2,     1,     1,    -1,    -2,    -2,     0,    -1,    -3,    -4,     0,     2,     1,    -2,     2,     3,     0,    -3,    -6,    -6,    -2,     0,    -1,    -4,    -1,     3,     5,     2,     7,     4,     0,     0,    -1,    -5,    -1,     1,    -2,    -1,    -2,     1,     1,     2,     0,     2,     0,    -2,    -6,    -9,    -6,    -1,    -1,    -4,     0,     1,     2,     6,     5,     4,     2,    -3,    -1,    -4,    -5,     2,     1,    -1,    -3,    -1,    -1,     3,    -1,     0,     0,    -3,    -6,    -5,    -5,     0,    -2,     2,     3,     0,     3,     5,     2,     0,     1,     1,     1,    -2,    -3,     1,     2,     1,     1,    -1,     0,    -2,     1,     0,     2,     2,    -1,    -6,    -4,     0,    -1,     4,     3,     4,     7,     3,     0,     1,     3,     1,     1,    -1,     1,     0,     3,     1,     1,     1,     1,    -1,     0,     0,     2,    -3,     1,    -8,     0,     0,    -1,    -3,     0,     2,     4,     7,     1,    -1,     0,    -1,    -2,     1,     0,    -1,    -2,     0,     0,     1,     0,     1,     1,     1,     0,    -2,     1,     1,     0,     0,     0,    -6,    -3,    -1,     1,    -1,     3,     0,     1,    -1,     2,    -1,    -1,     2,     1,     1,     3,    -1,     3,     1,    -1,    -2,     1,     1,     2,     5,     0,     0,     0,     2,    -1,     1,     0,     2,     1,    -1,    -1,     3,     2,     2,     3,     2,     2,     1,     1,    -5,    -2,     1,    -1,    -3,    -1,     3,     3,     6,    -1,     0,    -1,    -3,    -2,    -4,     0,     0,     0,     2,     3,     1,     1,     2,     3,     3,     2,     3,     1,     1,     0,    -1,    -1,    -1,    -3,     1,    -6,    -3,     0,     0,    -1,    -1,     3,    -6,    -6,     0,    -1,     0,    -1,     0,     0,     0,     1,    -2,     3,     3,     3,     1,     3,     3,     3,     6,     5,     4,    -1,     0,    -1,     0,     1,     0,    -2,    -4,    -4,    -6,    -8,    -4,    -2,    -1,     2,     3,     8,     4,     6,     2,     0,    -2,     1,     0,     0,     0,    -4,    -2,     0,     0,     0,     0,     0,    -1,     0,     1,     1,    -1,    -1,    -1,    -1,     0,     0,     1,    -1,    -6,    -3,    -1,    -1,    -2,    -2,    -4,    -5,    -4,    -3,    -1,     0,     0,     1),
		    86 => (    0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     2,     2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,     2,     2,     2,     2,     3,     1,     3,     2,    -3,     0,     0,     2,     2,     2,     3,     1,     1,     0,    -1,     0,     0,     0,     0,    -1,     1,     0,     1,     0,     2,     2,     3,     3,     2,     1,     3,     2,     1,     0,     2,     2,     3,     3,     5,     5,     3,     1,     1,     2,    -1,    -1,    -1,     0,    -2,     0,     0,     2,     4,     5,     4,     4,     5,     4,     2,     4,     3,    -1,     0,     3,     3,     0,     1,     4,     5,     4,     3,    -1,     0,     0,     0,     0,    -4,    -2,     2,     4,     5,     4,     1,     3,     5,     3,     4,     0,     1,    -2,     2,     3,     1,     2,     4,    -2,     0,     2,     2,     2,    -1,     1,     0,     0,    -3,    -3,     2,     3,     2,     3,     3,     4,     4,     1,     2,     0,     1,     0,     2,     1,    -2,    -2,     0,    -1,     2,     2,     2,     4,     1,     1,     0,     0,     0,    -1,     2,     1,     3,     1,     1,     4,     5,     1,    -1,    -1,    -1,    -1,     0,    -1,     1,     1,     1,     3,     1,     2,     2,     2,     0,    -1,     0,     0,     0,    -2,     1,     1,     0,     3,     2,     4,     2,     0,     0,    -2,     0,    -2,     0,     1,     4,     1,     3,     1,    -1,    -2,     1,     0,    -2,    -3,     0,     0,    -2,    -3,     3,     1,    -1,     1,     2,     2,     2,     0,     1,    -2,     1,    -1,    -2,     4,    -2,     1,     2,     4,    -3,    -4,    -4,    -6,    -4,    -5,     0,    -1,    -3,    -3,     1,    -1,    -1,     0,     2,     0,     0,     1,     1,    -1,     0,    -2,    -3,    -4,    -3,     2,     2,    -1,    -4,    -3,    -1,    -5,    -2,    -4,     0,     0,    -2,    -4,     1,    -2,    -2,    -2,    -1,     0,     1,    -2,     1,     0,     0,    -3,    -4,    -4,    -2,     1,     0,    -2,    -4,    -4,    -4,    -1,    -2,    -6,     0,     0,    -2,    -5,     0,     0,     0,    -2,    -4,    -2,    -1,     1,     2,    -1,    -2,    -2,    -1,    -1,     1,     1,     0,    -2,    -3,    -2,    -2,    -1,    -5,    -2,     0,     0,     0,    -3,    -1,     0,    -1,    -3,    -6,     0,     0,     1,     0,    -1,    -1,     0,     2,     5,     4,     1,    -1,     1,    -2,     4,     1,    -2,    -5,    -2,     0,     0,    -1,    -3,    -1,    -2,    -2,    -6,    -7,    -3,    -1,    -1,    -1,     1,    -1,     1,     2,    -1,    -1,     1,    -1,     1,     0,     5,    -2,    -3,    -4,     0,    -1,     0,    -1,    -3,    -3,    -1,    -4,    -4,    -5,    -2,     0,     0,     0,    -1,     0,     1,     0,    -2,    -3,    -2,    -2,     0,     2,     3,     0,    -1,    -1,     0,     0,    -1,    -1,    -3,    -4,    -3,    -3,    -1,    -7,    -6,    -2,     0,    -1,    -1,    -2,     1,     1,    -3,    -2,     1,    -1,     0,     0,     0,     0,     1,    -3,    -5,     0,    -1,    -2,    -6,    -1,     1,    -2,    -1,    -5,    -2,    -1,     0,    -2,    -3,    -1,     0,     1,     0,     1,     0,    -1,     1,     0,     0,     1,     1,    -3,    -4,     0,     0,    -1,    -5,     1,    -2,     0,     1,     0,     1,     1,     2,    -2,    -4,    -2,    -1,     1,     0,     1,     0,     0,    -1,     0,     3,     3,     2,    -2,    -6,     0,     0,    -1,    -6,    -1,    -2,    -1,     0,     1,     3,     4,     3,     2,    -1,    -1,     1,     1,     3,     3,     1,     2,     2,    -1,     2,     2,     3,    -2,    -3,     0,    -2,    -5,    -5,     0,    -1,     2,     2,     3,     1,     6,     5,     4,     1,     2,     0,     0,    -1,     0,     1,     1,     0,     0,    -1,     0,     0,    -2,    -1,     0,    -1,    -1,    -4,    -1,    -2,    -2,     5,     4,     4,     6,     5,     5,     3,     4,     4,     0,    -2,    -1,    -3,     1,     0,    -1,    -1,    -4,    -1,    -4,     0,     1,     0,    -3,    -2,    -2,    -3,    -2,     3,     9,     5,     4,     2,     3,     3,     4,     1,    -1,    -1,    -1,     2,     1,    -1,    -1,    -1,    -6,    -5,    -3,    -1,     0,     0,    -1,    -2,    -4,    -6,    -4,     0,     2,     4,     3,     3,     2,     0,     0,    -1,    -2,    -1,    -1,     0,     2,     1,    -1,    -2,    -8,    -4,    -3,     0,     1,     0,     0,    -3,    -2,    -3,    -3,    -3,    -3,     0,     0,    -1,     0,    -1,    -1,     1,     1,    -3,    -1,     3,     2,    -1,    -3,    -5,    -6,    -2,    -2,    -1,     0,     0,     0,     0,    -2,    -1,    -1,    -3,    -6,    -6,    -6,    -8,    -4,    -5,    -4,     0,     3,     4,     3,    -2,    -1,    -5,    -3,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,    -1,    -2,    -3,    -4,    -3,    -2,    -3,     0,     2,     1,    -2,    -2,    -3,    -2,    -2,    -1,    -5,    -2,    -3,    -4,    -1,     0,     1,     0,    -1,     0,     0,     0,    -1,    -2,     0,     0,     0,     0,    -1,    -1,     0,     1,    -1,    -1,     0,     1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0),
		    87 => (    0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -2,    -2,     0,    -3,    -5,    -4,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -3,    -5,    -1,    -1,     0,    -4,    -1,    -2,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -1,    -1,    -3,    -5,    -3,    -3,    -2,    -2,    -3,    -3,    -2,    -3,    -3,    -2,    -2,    -3,    -1,    -1,    -2,     0,     0,    -1,     0,     0,     0,     0,     0,     0,    -3,    -2,    -2,    -6,    -6,    -5,   -11,    -4,    -2,     0,    -1,    -2,    -5,    -4,    -4,    -4,    -4,     3,     0,    -3,    -4,    -2,    -1,     0,     1,    -1,     0,    -5,    -2,     5,     1,     3,     2,     2,    -2,    -6,    -6,     0,    -2,    -4,    -2,    -4,    -5,    -3,    -2,    -1,    -2,    -6,    -2,    -4,     0,     0,     0,     0,     3,     3,     3,     5,     3,     3,     2,     2,     5,     0,     0,    -3,    -3,    -3,    -2,    -1,    -3,     0,     0,     0,     2,    -5,    -1,    -3,    -2,    -1,     0,     1,     3,     0,     5,     5,     6,     7,     1,     6,     6,     3,     2,     2,     1,    -1,    -2,     0,     1,     0,     1,     0,     5,     1,    -1,    -3,    -1,    -2,    -2,    -1,     0,     1,     1,     2,     1,     5,     1,     3,     3,     3,     4,     1,     2,     2,     0,    -1,    -1,     0,     0,     0,     4,     0,    -3,    -5,    -3,    -2,    -1,     0,     4,     2,     2,     0,     0,     2,     2,     0,     0,     1,     5,     3,     4,     2,     1,     0,    -1,     0,     1,     0,     3,     1,    -5,     1,     4,     8,     0,    -2,     2,    -1,    -2,    -1,    -1,    -2,     1,     0,    -1,    -2,    -3,     0,    -1,     0,     0,     2,     2,    -1,     1,    -2,    -2,    -2,    -2,     3,     4,     7,     0,    -1,     1,    -2,    -2,    -4,    -2,    -1,    -2,    -1,    -4,    -1,    -4,    -5,    -2,     0,    -1,    -1,    -2,    -1,     0,    -3,     0,     1,    -4,    -5,    -4,     1,     0,     1,    -2,    -3,    -2,    -4,    -4,    -4,    -5,    -6,    -8,    -3,    -4,    -3,    -2,     1,     1,     0,     1,     1,     1,    -1,    -2,    -2,    -9,    -1,    -4,     1,     0,     0,     1,    -3,    -6,    -2,    -2,    -3,    -4,    -3,    -3,    -3,    -1,    -3,    -1,     3,    -1,     1,     1,     0,    -4,     2,    -2,     0,    -4,    -3,    -4,    -2,    -1,     1,    -1,    -1,    -2,    -1,     0,     0,    -2,    -2,     1,     0,     1,     1,     2,     1,    -2,     3,     2,     3,     0,     2,     0,     1,     0,    -3,    -3,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,    -3,    -1,    -2,    -1,     0,     1,     0,     1,    -2,     2,     2,     0,    -3,     4,     0,     2,    -1,    -3,    -1,    -2,     1,    -1,     0,    -2,    -1,    -1,    -1,    -1,    -1,     0,     2,    -1,     1,     2,     0,     0,     0,     0,     1,     0,     1,     0,    -1,    -2,     1,    -6,    -4,    -1,     0,     1,    -4,    -3,    -4,    -2,     2,     2,     0,     2,     3,     1,     2,     0,     0,    -1,     1,    -1,    -3,    -1,     1,     0,     0,    -1,     0,    -2,     1,    -3,     1,     0,    -1,    -2,    -3,     0,    -2,     3,     0,     0,     1,     0,     0,     0,    -2,    -2,    -2,    -1,    -3,    -1,    -1,    -3,    -1,    -1,    -2,    -3,     2,    -3,     0,     1,    -1,     0,    -2,    -4,    -1,     0,     0,    -1,    -2,     1,     0,     1,     0,    -1,    -3,    -2,    -5,    -3,    -4,    -5,    -2,    -1,     3,    -1,    -3,    -1,    -1,     2,    -1,    -2,    -6,    -5,    -3,     0,     1,    -1,    -2,     1,    -1,     0,    -1,    -2,    -1,    -6,    -6,    -4,    -4,    -4,    -5,     0,     1,    -4,    -4,    -1,     0,    -1,    -1,    -4,    -2,    -3,    -3,    -6,    -4,    -3,    -1,    -2,     0,     0,    -2,    -2,    -2,    -4,    -5,    -4,    -4,    -3,    -4,     0,    -1,    -2,    -1,     0,    -1,     0,    -1,    -6,     0,    -1,    -2,    -1,    -5,    -4,    -1,    -1,    -1,    -1,    -3,     0,    -1,     0,    -2,    -2,    -3,    -9,    -7,    -5,    -3,    -1,    -4,    -1,     0,     0,    -2,    -7,    -1,     0,     1,     1,    -5,    -2,     0,     0,     0,     0,     0,     0,    -1,     0,    -4,    -1,    -3,    -4,    -7,    -3,    -3,    -1,    -4,     0,     0,     0,     1,    -1,     2,     2,    -1,    -1,    -1,    -2,    -3,     0,    -1,     0,     0,    -1,    -2,     3,    -3,    -1,     1,     1,    -4,    -3,    -2,    -1,    -1,     0,     0,     0,    -2,     2,    -2,    -2,    -2,     4,     2,    -1,    -3,    -2,    -1,    -1,     0,    -3,     0,     0,    -1,     0,    -2,    -1,    -1,    -1,    -4,    -1,    -1,     1,     0,     0,    -1,    -2,    -8,    -6,    -7,    -2,     0,    -2,    -2,    -4,    -3,    -1,     0,     3,     0,    -2,     0,    -3,     0,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     1,     3,     4,     3,    -1,    -2,    -2,     3,     3,     4,     4,    -1,     0,     0,    -2,     0,     0,     0,     0,     0),
		    88 => (    0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -2,    -3,    -6,    -7,    -6,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,     0,    -2,    -2,    -3,    -4,    -3,    -1,     0,    -3,    -4,     1,     2,     0,    -3,    -4,    -4,     0,    -1,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -5,    -4,    -5,    -3,    -2,     1,     2,     2,     0,    -1,    -3,    -4,    -6,    -3,    -1,     1,     2,     0,     1,     2,    -2,    -1,     0,    -1,     0,     1,     0,    -3,    -6,    -4,    -4,     2,     1,     4,     4,     1,    -4,     0,    -2,    -2,     1,     0,    -3,    -2,     1,    -3,     1,     2,     2,     1,    -1,     0,     0,    -2,    -2,    -5,    -4,    -5,     0,    -2,     1,     3,     3,     1,     2,     0,     2,     3,     3,     1,     0,     0,    -1,    -4,    -3,     2,     1,    -2,    -2,     0,     1,    -4,    -4,     1,    -3,    -5,    -3,     0,    -1,     1,     1,    -1,     0,     2,     3,     2,     1,     1,    -2,    -1,     0,     1,     1,     0,     2,     0,    -1,     0,    -4,    -2,     1,     2,    -2,    -3,     0,     1,     1,     0,     0,    -1,    -1,     0,     4,     4,     1,     0,    -2,     1,     1,     3,     4,     1,     1,     0,    -3,    -2,    -3,    -2,     5,     3,     0,     1,     1,    -3,     1,     1,     0,    -1,     1,     1,     2,     2,     1,     1,    -1,    -1,    -2,     0,     2,    -1,     1,     2,     0,     0,    -2,    -3,     3,     6,     0,     0,    -2,    -1,     1,     0,    -2,    -1,    -1,     0,     2,    -1,    -2,    -1,     1,     0,     0,    -2,     0,    -1,     4,     5,    -4,    -1,    -2,    -4,    -2,     3,     0,    -1,     0,    -2,    -3,    -3,    -3,    -2,     2,     2,    -1,    -5,    -3,    -3,    -2,     0,    -2,     1,     1,     2,     1,     4,    -3,     1,    -1,    -3,    -1,     2,     0,     2,    -1,    -2,    -1,    -4,    -2,     0,     2,     0,    -5,    -5,    -3,    -2,    -1,    -1,    -1,    -1,     3,     1,    -3,     2,    -3,     0,     0,    -1,     1,    -3,     0,    -4,    -4,    -3,    -3,    -1,     2,     2,     1,     2,     0,    -2,    -3,    -1,    -2,     1,     0,     1,     0,    -2,    -7,    -7,    -4,     0,     0,     0,    -1,    -3,    -2,    -3,    -3,    -2,     4,     4,     3,     4,     2,     0,     1,     0,    -1,     1,    -1,     1,     3,     2,     0,    -4,    -6,    -5,     0,    -1,     0,    -1,    -2,    -3,     0,     1,    -1,     2,     4,     4,     5,     4,     3,     0,     1,     0,    -1,     0,     2,     3,     3,    -1,    -3,    -2,     0,    -3,    -1,    -1,     0,    -1,    -1,    -4,    -1,     3,     3,     3,     5,     6,     3,     3,     4,     1,     1,     1,     0,     2,     2,     2,     1,     1,    -3,    -3,     4,    -5,    -2,    -1,     0,    -2,    -2,    -3,    -2,    -1,     3,     1,     4,     5,     4,     2,     0,     0,     0,     2,     5,     4,     1,     3,     2,     0,     0,     0,     2,    -6,    -2,     0,    -1,    -3,    -2,     1,    -3,    -3,     0,     0,     0,     2,     1,    -1,    -2,    -1,     3,     0,     1,     2,     1,     1,    -1,    -1,     1,     1,    -2,    -1,    -3,    -1,    -1,    -3,    -5,    -2,    -3,    -1,    -2,    -2,     0,    -1,    -2,    -2,    -1,     2,    -1,     0,    -2,     0,    -1,    -4,    -3,    -1,     2,    -1,    -4,     0,    -1,     0,     0,    -2,    -6,    -3,    -5,    -4,    -4,    -4,    -3,    -2,    -2,     0,     2,     3,     1,     2,    -1,    -1,    -3,    -2,     0,     1,     1,    -2,    -5,    -3,    -2,    -1,     0,    -3,    -5,    -3,    -3,    -3,    -1,     0,    -3,    -2,    -2,     2,     3,     4,     3,     1,     1,    -2,     0,     1,     1,     0,     0,    -4,    -4,    -3,     0,    -1,    -1,    -3,    -1,    -2,     0,     0,     0,     0,     0,    -2,     3,     7,     3,     2,     4,     2,     2,     0,     0,     1,    -2,    -1,     0,    -2,    -2,    -4,    -1,    -1,    -1,    -2,     0,     3,     1,     0,    -2,    -2,     0,     1,     3,     2,     1,     5,     4,     1,    -1,    -1,    -2,     1,    -2,     1,     2,    -2,    -3,    -3,    -1,     0,     0,    -1,     0,     1,     1,    -1,    -3,    -2,     3,     3,     0,     2,     5,     4,     3,     1,    -2,    -1,     0,     2,     0,     2,     2,    -5,    -4,    -2,     0,     0,     0,    -2,    -1,    -1,    -2,    -2,    -3,    -2,     0,    -1,     1,     4,     6,     4,     0,    -1,    -2,     1,     5,     4,     1,    -3,    -2,    -6,    -3,    -1,     0,     0,     0,    -2,     0,    -6,    -4,     0,    -2,    -4,    -4,    -1,     3,     3,     3,     1,     1,    -4,    -1,     0,     1,    -2,    -6,    -5,    -3,    -3,    -1,    -2,     0,     0,     0,     0,    -3,    -2,    -2,    -4,    -3,     3,     2,    -2,    -1,    -1,     1,     0,    -5,    -2,    -2,    -3,    -4,    -7,    -5,    -3,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,    -3,    -5,    -2,    -1,    -1,    -3,    -5,    -4,    -4,    -3,    -2,    -1,     0,     0,    -1,     0,     1,     0,     0,     0),
		    89 => (    0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -3,    -2,     0,     0,    -1,     0,    -2,    -2,     0,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,    -3,    -1,     0,     0,    -1,    -1,     0,    -1,    -2,     0,    -1,    -3,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,    -1,     0,     0,    -1,     0,     1,     1,    -1,    -2,    -3,    -2,    -3,    -1,    -1,     0,    -2,    -2,    -3,    -3,    -3,    -2,    -3,    -4,    -3,    -2,    -2,    -1,     0,     0,    -1,     0,     1,     0,     1,     0,    -1,    -2,    -1,    -3,     1,    -2,    -1,    -1,    -3,    -5,    -4,    -2,    -2,    -1,    -1,    -2,    -4,    -5,    -2,    -1,    -1,     0,    -3,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -4,    -2,    -2,    -2,     0,    -1,     0,    -2,    -1,    -2,     0,    -1,    -3,    -2,     0,    -1,    -1,     0,     0,     0,    -1,    -2,     0,    -1,    -3,    -2,    -6,    -3,    -2,    -2,    -1,     1,     4,     2,     1,     2,     0,     0,     1,     0,    -2,    -2,    -1,    -2,    -1,    -1,     0,     0,    -1,     0,    -2,    -3,    -4,    -4,    -6,     0,    -1,     2,     2,     0,    -1,     2,     0,     0,    -1,     0,     0,    -1,    -2,    -2,    -3,    -1,     0,    -1,    -2,    -2,    -1,    -2,    -1,    -4,    -3,    -6,    -2,    -3,     1,     0,    -2,     0,     0,    -5,    -2,     0,    -1,    -1,     0,    -2,    -2,    -3,    -5,    -1,    -1,     0,     0,     0,    -1,    -2,    -4,    -5,    -3,    -4,     0,     1,     0,     2,    -1,    -1,     1,    -3,    -3,    -1,     3,     1,     1,    -2,    -2,    -1,    -2,    -5,     0,    -2,     0,    -1,    -2,     0,    -1,    -1,    -2,     1,     1,     0,    -3,    -2,    -4,    -3,    -2,    -2,    -4,    -3,     3,     0,    -1,    -3,    -1,     0,    -2,     0,    -1,    -2,     0,    -4,     0,     2,     0,    -2,    -2,     0,     1,    -1,    -2,    -5,    -3,    -1,    -1,    -2,    -2,     0,    -2,     0,     0,    -1,    -1,     2,    -3,    -1,    -1,    -2,    -1,    -1,     1,     1,     1,     1,     1,     0,     2,    -1,    -2,    -5,    -1,    -3,    -5,    -3,    -2,    -1,    -3,    -1,     0,     2,     0,     1,    -5,    -2,    -1,    -1,    -1,    -3,    -2,     3,     2,     1,     1,     0,    -1,    -4,    -2,    -2,    -4,    -3,    -1,    -1,     1,    -3,    -3,    -1,     0,     2,     0,    -2,    -4,    -2,    -1,     0,    -1,    -2,    -3,     0,     2,     1,     1,     1,     3,    -3,    -2,    -5,    -4,    -3,    -2,     1,     0,    -2,     2,     2,     0,     0,     1,    -4,    -3,    -2,     1,     0,     0,     0,    -3,    -1,     0,     0,     2,     1,     1,    -3,    -1,    -5,    -4,    -4,    -2,    -2,    -2,    -3,     1,     1,     3,     1,     1,    -6,    -5,    -1,     1,     0,     1,     0,    -3,    -2,     1,    -2,     3,     0,     0,    -1,     2,    -1,     0,    -1,    -2,    -3,    -4,    -2,     3,     1,     2,    -1,    -1,    -5,    -2,    -2,     0,     0,     0,     0,    -2,    -2,     2,    -2,     0,     2,    -2,     0,    -1,    -1,    -1,    -3,    -1,     0,     0,     0,     1,     1,     1,    -1,    -1,    -3,    -1,    -1,    -2,    -1,     0,     0,    -2,    -1,     2,     2,     2,     0,    -2,     0,     3,     1,     2,     0,     1,    -1,    -2,     1,     2,     1,    -1,     1,     1,    -2,    -5,     0,    -2,    -2,     0,     0,    -1,    -1,     1,     4,     3,     5,    -1,     0,     3,     6,     1,    -1,    -2,     0,     0,     0,     3,    -2,    -1,    -1,    -1,    -2,    -2,     1,    -3,     0,     0,    -1,    -1,    -1,     0,     2,     1,    -1,     1,     1,     0,     0,     0,    -2,    -4,    -2,    -1,     1,     3,    -1,    -1,     0,    -1,    -1,     3,     1,    -2,     0,     0,     0,    -2,    -2,    -3,    -1,     1,     2,     1,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     0,     1,     0,     1,    -2,     0,     0,     4,    -1,    -5,     1,     0,     0,    -1,    -1,    -2,    -2,    -3,    -3,     0,     0,    -2,    -3,    -1,    -3,     2,     1,    -1,    -1,     0,     0,     1,     0,     1,    -1,     3,     1,    -4,     0,     0,     0,    -1,     1,    -2,    -2,    -2,    -3,    -3,    -5,    -6,    -5,    -4,    -1,     1,     3,    -2,    -1,    -2,     2,     1,     1,     4,     0,     4,     1,    -2,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -2,    -3,    -5,    -4,    -1,     3,    -1,     0,     0,    -1,     1,     1,     2,     3,     4,     3,     3,     1,     0,     0,     0,     0,     2,    -1,    -1,     1,    -1,    -2,    -2,    -2,     0,     1,     2,     3,     0,    -2,    -3,    -3,    -1,     4,     5,     3,     5,     2,     2,    -1,    -1,     0,     0,     0,     0,     1,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -2,    -1,    -4,    -5,    -3,    -1,     0,     4,     2,     2,     2,     0,     0,     1,     1,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -2,    -1,    -2,    -4,    -2,    -2,    -1,    -2,     0,    -1,     0,     0,     0,     0),
		    90 => (   -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -1,    -1,     1,     1,     1,     0,     0,     0,    -1,    -1,     1,     0,     0,     0,     0,     0,     1,    -1,    -1,    -2,    -2,     1,     0,     0,     0,    -2,    -1,    -1,    -1,    -1,     2,     2,     1,     2,     2,     0,     0,    -1,     0,    -1,    -1,     0,     1,     0,    -1,     0,     0,    -1,     1,    -2,    -1,    -1,    -1,    -1,     0,     0,    -1,    -1,     0,    -1,     0,     2,     2,     0,    -1,    -1,    -1,    -1,     0,    -2,     1,     0,    -1,    -1,    -1,    -2,     1,     1,     0,    -1,    -1,     0,    -1,    -1,    -1,    -1,     1,     1,     0,     1,     2,     1,    -1,    -1,    -1,    -3,    -1,     0,     0,    -1,    -1,    -1,     0,     1,     2,     0,    -1,     1,     1,     0,     1,     1,     0,     2,     1,     1,     3,     1,     0,     1,     2,     0,     0,     0,    -2,     0,     0,    -1,     1,    -1,     1,     1,     1,     2,     1,    -2,    -1,     0,     1,    -1,     0,    -1,     0,     1,     0,     1,     2,     2,     1,     1,    -1,    -1,    -1,    -1,    -1,     0,     1,     0,     3,     0,    -1,     0,     1,     1,    -1,    -3,    -3,    -3,    -2,    -3,    -1,    -1,     0,     0,     0,     3,     2,    -1,     1,    -1,     0,     0,     0,     0,     0,     0,     0,     2,     2,     2,     2,     0,    -3,    -2,    -3,    -2,    -1,     0,    -3,    -2,    -2,    -1,    -1,    -1,     2,     0,    -1,    -1,    -1,     0,     0,     2,     0,    -1,     2,     2,     1,    -1,     0,    -3,    -3,    -4,    -3,     0,     1,     1,    -2,    -2,    -3,    -4,    -3,    -2,     0,     0,     2,     0,     0,     0,     0,     0,     0,    -1,     2,     1,     1,    -1,     0,    -2,    -3,    -4,    -3,     0,    -1,    -1,    -4,    -4,    -3,    -3,    -3,    -1,     0,    -1,     1,     1,     0,     1,     1,     0,     0,     0,     3,     0,     3,    -1,    -2,    -3,    -5,    -5,    -2,    -1,    -1,    -2,    -4,    -3,    -3,    -3,    -3,    -2,     0,     1,     1,     0,     0,    -1,     0,     0,     0,    -2,     3,     2,    -1,    -2,    -3,    -4,    -3,    -3,    -3,    -2,    -1,    -3,    -3,    -3,    -3,    -3,    -3,    -1,    -2,    -1,    -2,     1,    -1,     0,     0,     0,     0,     0,     3,     1,    -1,    -2,    -2,    -3,    -3,    -3,    -2,    -2,    -2,    -1,    -1,    -2,    -2,    -3,    -3,    -1,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,     0,     2,     2,     2,     0,    -1,    -2,    -2,    -2,    -2,    -2,     1,    -1,    -1,    -4,    -4,    -4,    -1,    -3,    -1,     2,     0,     1,    -1,     1,     0,     0,    -1,     1,     3,     2,     2,     2,    -1,    -2,     0,     0,    -1,    -2,    -1,    -2,    -4,    -4,    -4,    -3,    -2,     0,     1,     0,    -1,     1,    -3,     1,     0,     0,    -1,     0,     4,     1,     1,     2,     0,    -1,     0,    -1,    -1,    -1,    -3,    -1,    -3,    -3,    -4,    -3,    -1,     1,     0,     1,     0,    -1,    -1,     0,     1,     0,     1,     0,     2,     0,     1,     1,    -1,     0,     1,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,     0,     1,     0,     0,    -1,     0,    -2,    -1,     0,    -1,     0,     1,     0,     2,    -1,     2,     1,     0,    -2,    -1,     1,    -1,     0,     1,     0,     1,     2,    -2,     0,     0,     0,     1,    -1,     0,    -2,     0,     0,     0,     0,    -1,     0,     0,    -2,     0,     2,     0,     0,    -1,     1,    -1,     0,     0,     0,    -1,     0,     0,     1,     1,     0,    -1,     0,    -1,     0,     1,     1,     1,     0,     0,    -1,    -1,    -1,    -2,     2,     1,    -1,     0,     1,    -1,     0,    -1,    -1,     1,     1,     0,     1,     1,    -1,    -1,    -1,    -2,     0,     1,     1,     1,     0,     0,    -1,    -1,    -1,     1,     2,    -1,    -1,     0,     0,     1,    -1,    -1,     0,    -1,     0,    -1,     1,     0,     0,     0,    -1,    -2,    -2,    -1,     0,     0,     0,    -1,    -1,    -1,     0,     2,     2,     1,    -1,     0,     0,    -1,     1,     1,     1,     0,     1,     1,    -1,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     1,     3,     3,     1,     0,     0,    -1,    -1,    -2,     0,     0,    -1,    -3,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,    -2,     0,    -1,     0,    -1,     0,     0,    -1,    -1,    -1,    -2,    -5,    -3,    -3,    -3,    -2,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,     0,     0,     0,    -1),
		    91 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     1,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     3,     2,     2,    -2,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,    -1,     0,     1,    -2,    -2,    -2,    -2,    -1,     1,     1,     2,     5,     3,     3,     1,     2,    -3,    -3,    -3,     0,     0,    -1,     0,     0,     0,     4,     2,     0,    -2,    -4,     2,     1,     1,    -3,    -4,    -2,     0,     0,     0,     1,     0,     0,    -3,    -1,    -2,    -2,    -2,    -2,     0,     0,     0,     0,     0,     4,     4,     3,     0,    -1,     1,     3,     2,     1,     0,    -3,     1,    -1,     1,    -1,     0,     0,    -3,    -3,    -1,     3,     2,     2,    -1,    -1,    -2,     0,    -1,     1,     1,     4,     4,     1,     1,     2,     0,    -1,     0,    -1,    -1,    -3,    -1,    -1,    -1,    -1,    -1,    -3,     1,     3,     4,     3,    -3,    -1,    -2,    -1,     0,    -2,     0,     4,     2,     1,     0,    -3,    -2,    -1,    -1,     1,    -1,    -1,    -2,    -3,    -2,    -1,    -5,    -1,     2,     3,     3,     1,     0,    -1,    -1,     0,     0,    -2,    -2,    -2,    -2,    -3,     2,    -5,    -1,     4,     3,     3,    -1,     1,    -2,    -4,    -2,    -1,    -3,    -1,     2,     3,     4,     1,    -2,    -2,    -1,    -1,     0,    -3,    -2,    -2,    -2,    -2,     3,    -4,    -1,     4,     0,     3,     0,    -1,    -1,    -2,    -3,    -3,    -3,     2,     2,     2,     1,     1,    -1,    -3,    -1,     0,     0,    -3,     0,    -2,    -2,    -2,     4,    -1,     1,     2,     0,    -2,    -3,    -2,    -2,    -3,    -5,    -3,    -4,     0,     0,     2,     1,     0,    -1,    -2,    -1,     0,     0,    -2,     0,    -2,    -1,    -2,     1,     1,    -2,     3,     0,     0,     0,    -1,    -2,    -4,    -4,    -1,    -1,     0,     0,     2,     2,    -1,     0,     1,     1,    -1,     0,     0,     0,     0,    -2,    -3,     2,    -2,    -1,     0,    -2,    -1,    -2,     2,     0,    -3,    -1,    -1,    -1,    -1,    -2,     2,     1,    -1,     0,     0,     3,    -1,     0,    -2,     0,     1,    -1,    -1,    -2,    -3,    -3,     0,     0,    -1,    -2,     1,    -1,    -1,    -1,    -1,    -1,    -1,    -2,     0,     1,    -2,     1,     2,     3,     0,     0,    -1,     0,    -1,    -1,     0,    -1,     0,    -1,    -1,    -1,     1,    -1,     0,     0,    -2,    -1,    -3,    -1,    -2,    -2,    -2,    -5,    -2,     2,     1,     1,     0,     1,     1,     1,    -1,    -2,     1,    -1,    -1,    -2,    -4,    -6,    -2,     2,     1,     1,     0,    -1,    -1,    -4,    -3,    -3,    -4,    -2,    -1,    -3,     0,     0,     0,     0,     0,     0,    -1,    -4,    -2,    -2,    -3,    -4,    -7,    -6,    -2,     1,     2,    -2,    -3,     1,     0,    -3,    -4,    -2,    -4,    -2,    -5,    -4,    -3,    -1,     0,    -1,     0,     0,    -1,    -1,    -2,    -2,    -3,    -1,    -3,    -2,    -3,    -1,     3,     1,    -1,     1,     1,    -1,    -1,     0,     0,    -2,     3,    -4,    -3,    -1,     1,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     2,     1,    -2,    -1,     2,     0,     1,    -1,     1,     0,     2,     2,     2,    -1,     0,    -3,    -2,    -2,     0,    -1,     0,    -2,    -1,     0,    -3,     0,     2,     3,     2,    -3,    -3,    -2,     1,     0,     1,     2,     0,     1,    -2,    -1,     1,     0,     1,     0,    -2,     0,    -1,     0,     1,    -2,    -1,     0,     4,     4,     5,     5,     4,     1,    -4,     0,    -1,     2,     3,     0,     1,    -2,     0,     0,     2,     5,     2,     2,    -2,    -1,     1,     0,     0,    -1,     1,     3,     4,     4,     3,     3,     2,     0,    -1,     0,     1,     0,     2,     0,     0,     1,     3,     3,     4,     2,     1,     0,    -1,     0,     1,     1,    -1,     0,    -1,    -3,    -1,     0,     0,    -1,    -1,    -3,    -1,     1,    -2,     0,    -3,    -2,     0,     1,     1,     0,     2,     1,     0,     2,    -1,     0,     2,     1,    -2,    -1,    -1,     2,     0,    -1,    -3,    -3,    -3,    -3,     1,     0,     0,     1,    -3,    -1,     0,     0,     0,     0,    -3,    -2,    -1,     0,     1,     0,    -1,     0,    -1,    -1,     1,     3,     3,     1,     0,     0,     1,     0,     3,     1,    -2,    -2,    -2,     1,    -1,    -1,     2,     0,    -1,    -2,    -2,    -2,     3,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,     1,     1,    -1,     0,    -2,    -4,    -2,    -2,    -1,    -4,     0,    -3,    -1,    -1,    -3,     2,     3,     0,    -1,     0,     0,    -1,    -1,    -1,     0,    -1,    -2,    -1,    -2,    -1,     0,     2,     2,    -2,    -3,    -2,    -2,    -2,    -4,    -3,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -3,    -3,    -2,    -1,    -1,    -1,     0,    -1,    -2,    -3,    -2,    -2,    -2,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,     0,    -1,    -2,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0),
		    92 => (    0,     1,     1,     0,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,    -1,     1,     1,     1,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,    -1,     1,    -1,    -2,    -3,    -4,    -1,    -1,     0,     2,     2,     0,    -2,    -5,    -3,    -3,    -2,     0,     1,     0,     0,     0,     0,     0,     0,    -1,    -2,     0,     1,     0,     0,     4,     4,     5,     0,     1,     3,     6,     5,     2,    -2,    -4,    -2,    -1,    -2,    -1,     0,     0,     1,     1,     0,     0,     0,    -3,    -4,     2,     2,     3,     0,    -3,    -4,    -6,    -7,     0,    -1,     0,     0,    -2,    -5,    -4,    -3,    -1,     0,    -3,    -4,     0,    -1,     0,     0,     0,    -1,    -3,     0,     1,     6,     5,     3,     6,     2,    -1,    -2,    -2,    -1,     1,    -2,    -1,     1,    -1,    -1,    -3,     0,    -3,    -5,     0,    -3,    -1,     0,     0,    -2,    -1,     0,    -2,    -2,     0,     4,     1,     3,     0,     1,     1,     1,     1,     0,     1,     2,     2,     1,     3,    -1,    -2,    -4,     1,    -5,    -1,     0,     0,     0,     0,     1,    -1,    -1,    -1,     2,     0,     1,    -3,     1,    -2,     0,     0,     2,     1,     2,     1,     0,     1,    -1,    -2,    -7,    -1,    -5,    -1,    -1,     0,     2,     0,     2,     5,     2,     1,     2,    -1,    -4,    -2,     0,     1,    -1,     1,     2,    -2,     1,    -1,     1,     3,     3,    -5,     1,     3,    -3,    -2,    -3,     3,     2,     1,     0,     4,     2,    -1,     1,     1,    -1,     1,     1,     0,     0,    -3,    -2,    -1,    -2,     1,     0,    -2,     0,     3,    -1,    -2,    -5,    -2,     0,    -2,     1,     2,    -3,     0,     0,    -2,     0,    -1,     0,     2,     2,     2,    -1,     0,    -1,     0,     0,    -1,     0,    -1,     3,     0,    -2,    -7,    -1,    -1,     1,     0,    -1,     1,    -1,     3,     5,     1,     1,    -2,     3,    -1,     0,     0,    -1,     0,    -1,     3,    -2,    -2,     0,     1,    -1,    -4,    -3,    -2,    -2,    -2,     0,    -3,     0,     0,    -1,     1,     2,     2,     1,     2,     2,    -1,    -2,    -3,    -1,    -3,    -1,    -2,     0,     1,     1,     0,    -3,    -3,     1,     1,    -2,    -3,     0,    -1,    -5,     0,    -2,     0,     4,     2,     0,     3,    -1,    -3,    -2,    -1,    -3,    -3,    -3,    -2,     2,     4,    -1,     3,     3,    -3,     3,     1,     0,    -1,     0,    -3,    -2,    -1,    -1,     2,     7,     2,    -1,     0,    -1,     0,    -1,     1,    -3,    -2,    -3,    -1,     1,     2,    -1,     1,     3,     6,     4,     5,     5,    -1,     0,     0,    -1,     1,     2,     3,     5,     5,    -3,     2,     0,    -4,    -2,    -3,    -2,    -1,    -1,     0,     0,     2,    -4,     2,     5,     8,     7,     3,     3,     1,     0,    -2,     4,     4,     0,     1,     2,     2,     3,     1,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -2,    -1,    -2,     1,     3,     3,     2,    -1,     3,     6,     4,     0,     0,     5,     4,    -3,    -2,     0,     4,     2,     4,     2,     0,     2,     0,    -1,    -1,    -1,    -2,    -1,     1,    -1,     9,     7,     4,     1,     5,     6,     3,     0,    -1,     4,     3,    -1,    -2,     1,    -1,    -1,    -1,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,     3,     9,     5,     2,     1,     2,     2,     2,     0,     0,     1,     2,    -1,    -1,     0,    -2,     1,    -1,    -2,     0,     1,     0,    -3,    -2,    -2,    -3,     0,     2,     8,     7,     5,     4,     3,     3,    -1,     1,     0,    -2,     1,    -1,     0,     0,    -1,     0,     1,     1,     2,     2,    -1,    -2,     1,     2,    -1,    -3,     1,     4,     5,     7,     5,     2,     0,    -2,     1,     3,    -1,    -1,     4,    -2,    -1,     0,     0,     0,     0,     2,     3,     3,     0,     0,    -2,     0,    -3,    -1,     2,     5,     7,     8,     3,     3,     1,     1,     1,    -1,     0,     0,     4,    -2,     3,    -1,     1,     0,     3,     5,     3,     0,     1,     1,    -3,     0,    -1,    -3,     6,     9,     7,     6,     8,     1,    -1,     1,    -1,     0,     0,     0,    -1,    -3,    -1,     1,    -2,     0,     3,     2,     1,     1,    -2,     0,    -2,    -1,     0,     2,     8,     8,     7,     5,     5,     2,    -3,     1,     0,     0,    -1,     0,     0,    -4,     0,     1,     2,     1,     1,     4,     2,     1,     1,     1,    -2,    -1,     5,     9,     7,     5,     7,     7,     5,     3,    -3,     0,     0,    -1,     0,     0,    -3,    -1,    -2,    -4,     2,    -2,     0,     2,     2,     1,    -4,    -6,    -1,     1,     6,     8,    11,     7,     4,     6,     4,    -1,     1,     0,     1,     0,     1,     0,    -1,    -1,    -4,    -7,     2,    -2,    -2,    -3,    -4,    -4,    -5,    -5,     1,     1,     1,     4,     7,     2,     0,     1,    -3,    -2,    -1,     0,     1,     0,     1,     1,     0,    -1,    -1,    -2,    -4,    -6,    -3,    -7,    -8,    -6,    -6,    -8,    -8,    -7,    -7,    -6,    -5,    -8,    -2,    -1,    -3,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -1,    -3,    -4,    -3,    -3,    -4,    -2,    -2,    -2,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     1),
		    93 => (    0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,    -3,    -3,     4,     1,    -1,    -2,    -4,    -2,    -2,    -2,    -2,    -1,    -4,    -3,    -4,    -2,     0,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,     1,     2,    -2,    -4,    -5,    -4,    -5,    -6,    -7,    -4,    -3,    -4,    -5,    -3,    -3,    -2,    -1,    -3,    -1,    -1,     0,     0,    -1,     0,     0,     0,     1,     4,     4,    -2,    -1,    -5,    -1,    -1,    -1,    -4,    -6,    -6,    -5,    -5,    -5,    -5,    -4,    -1,    -2,    -2,    -1,    -2,     0,     1,     1,     0,     0,     1,     2,     3,     0,    -1,     0,     2,     3,     2,     2,    -1,    -2,    -1,    -2,    -2,    -4,    -5,    -3,    -3,    -3,    -1,    -1,    -3,    -1,     1,     0,     0,     0,     2,     1,    -2,     1,     3,     0,     2,    -1,     2,     1,    -2,    -2,    -3,    -4,    -3,    -2,    -5,    -4,    -3,    -3,    -3,    -2,     0,    -2,     0,     0,     1,     0,     2,     0,    -1,     3,     1,     2,     0,    -1,    -3,     0,     0,    -1,     2,    -3,    -4,    -5,    -6,    -4,    -3,    -3,    -3,    -2,     0,    -1,    -1,     0,     0,    -2,     1,     0,     0,    -1,    -3,    -1,    -1,    -3,     0,     3,     4,     4,     3,    -1,    -5,    -6,    -6,    -5,    -2,    -3,    -3,    -2,    -1,    -1,     0,     0,    -2,    -2,     0,    -1,     1,    -2,    -1,    -3,    -1,    -1,     2,     3,     4,     4,     0,    -3,    -7,    -7,    -7,    -4,    -2,    -2,    -1,    -2,    -2,    -2,     0,     0,    -3,    -1,     3,     0,     2,     0,    -1,    -2,     0,     0,     2,     3,     2,     1,    -2,    -3,    -7,    -8,    -6,    -5,    -5,    -2,     0,    -1,    -1,    -1,     0,     0,    -4,     0,     4,     3,     1,    -1,     0,    -1,     1,     2,     1,     2,     0,    -2,    -2,    -3,    -3,    -3,    -4,    -3,    -4,    -3,    -1,     0,    -3,    -2,     0,     0,    -3,    -4,     3,    -1,     0,    -3,    -2,     2,     1,     3,     3,     2,     0,     0,     0,    -3,    -3,     1,     0,     0,     2,     3,     2,    -2,    -2,    -1,     0,     0,    -1,    -3,     3,     2,     1,     0,    -1,     1,     2,     2,     2,     2,     2,     1,    -1,     0,     0,     1,     0,    -1,     1,     2,     3,     3,    -3,    -2,     0,    -1,     1,     0,     2,    -3,    -2,    -2,    -1,     1,     2,     1,     0,    -1,     0,    -2,    -1,     1,    -2,     0,     3,     0,     0,     0,     5,     2,    -3,    -1,    -1,     0,     2,     0,     1,    -3,    -3,    -2,     0,     1,     0,    -1,    -2,    -2,    -2,     0,    -2,     0,     0,     0,     2,     3,     2,     2,     2,     0,    -3,     0,     0,     0,     1,     0,     0,    -3,    -5,    -2,    -3,     1,     3,    -2,    -3,    -2,    -4,    -5,    -2,    -2,    -2,     0,     1,     3,     3,     3,     0,     0,    -2,    -2,    -1,     1,     0,    -1,     2,    -1,    -2,    -2,    -4,    -2,    -2,    -5,    -3,    -3,    -3,    -5,    -5,    -3,    -3,    -4,     2,     1,     4,     2,     2,     0,    -2,    -1,     0,     0,     0,     1,     0,     0,    -1,    -3,    -2,     0,    -1,    -5,    -2,    -1,    -2,    -2,    -4,    -2,     0,    -1,     0,     1,     2,     2,     0,     1,    -2,    -1,    -2,     1,     0,    -1,    -1,    -2,    -1,    -1,     1,     0,    -1,    -2,    -1,     1,     1,     1,    -1,     1,     2,    -1,     0,     0,     1,     1,    -1,     1,     0,    -3,    -1,     1,     0,    -1,    -3,    -2,    -2,    -3,     0,     1,     1,    -1,     1,     1,     2,     2,     2,     3,     0,    -1,    -1,     2,     2,     1,     0,     1,    -1,    -1,     0,    -1,     0,     0,     0,     2,    -1,    -4,    -3,    -2,    -1,    -2,    -2,    -2,    -1,     1,     0,     0,    -1,    -2,     0,     0,    -3,    -1,     1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,    -3,    -3,    -3,    -3,    -2,    -3,     0,     0,    -2,    -1,    -3,    -3,    -1,    -1,    -1,    -1,    -1,     1,    -2,    -1,     0,     0,     0,     0,     1,    -2,     0,    -1,    -1,     0,    -1,    -1,    -2,     0,     1,    -1,    -2,    -1,    -2,    -1,    -3,    -1,    -2,    -2,    -1,    -3,    -1,    -1,     0,     0,     0,     0,     1,    -1,    -2,    -1,     1,     2,     1,     0,     0,     4,     1,    -2,     0,    -1,    -2,    -3,    -2,    -1,    -2,     0,    -1,    -3,    -2,    -1,     0,     0,     1,     0,     0,    -2,     0,    -1,     0,     1,     1,     0,    -1,    -1,    -1,     2,     1,    -1,    -2,    -2,     0,    -1,    -4,    -3,    -3,    -4,     0,     0,     0,     1,     0,     1,     0,    -1,    -1,    -2,    -1,    -2,    -3,    -3,    -1,    -3,    -2,     0,    -3,    -1,     0,     0,    -2,    -2,    -2,    -1,    -3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -1,    -2,    -2,    -3,     0,     0,     0,    -2,    -1,    -1,    -1,     0,     0,     0,     1,     0),
		    94 => (    0,    -1,     0,     0,     0,     1,     0,     0,     0,     0,     1,     0,    -1,     0,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     1,     0,     0,     0,     0,    -1,    -2,    -1,    -2,    -2,    -2,    -3,    -2,    -1,    -3,    -3,    -2,     0,     0,    -3,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,    -3,    -5,    -1,    -2,    -3,    -2,    -3,    -4,    -7,    -5,    -3,    -4,    -2,    -1,    -2,    -3,    -3,    -3,    -1,    -2,    -2,    -3,    -2,    -1,     0,     0,     0,     0,    -4,    -6,    -1,    -4,    -4,    -2,    -3,    -4,    -2,    -2,    -5,    -3,    -2,     2,    -2,    -4,     0,    -1,     0,     1,     1,    -3,    -2,     0,     1,     1,     0,    -2,    -3,     0,    -2,    -4,     0,     0,    -1,    -4,     0,     2,    -2,    -2,    -5,    -2,    -3,    -3,     3,     2,     2,     0,    -2,    -3,     1,    -1,     0,     0,     0,    -2,    -3,    -3,    -2,    -3,     0,     1,     1,     4,    -1,    -1,    -2,    -4,    -5,    -2,     1,     6,     1,     0,     1,    -2,    -2,    -3,     1,    -2,     0,     0,     0,    -1,    -1,    -2,    -2,    -1,     0,    -1,    -1,    -4,    -2,    -2,    -1,    -6,    -9,    -2,     0,     3,     3,     5,     5,    -2,    -1,    -3,    -2,    -1,    -2,     1,    -1,    -2,     0,    -2,     0,    -1,     3,    -1,    -2,    -3,     1,     2,    -2,    -7,    -6,    -1,     1,     2,     2,     2,     1,    -2,    -2,    -4,    -3,    -1,    -2,    -2,    -3,     2,     0,    -1,     0,     1,     2,    -2,    -3,    -3,     1,     0,    -3,    -4,    -3,    -3,     5,     1,     2,     0,    -3,    -3,    -4,    -3,    -1,    -3,    -1,     0,    -3,     2,    -1,    -2,    -2,     0,    -1,    -1,    -1,    -4,     0,    -1,    -1,    -3,    -4,     0,     3,     1,    -1,     0,     2,     1,    -3,    -3,    -1,    -1,    -1,     0,    -2,     2,     3,     0,    -2,    -3,     0,     1,    -2,     1,     0,    -1,    -1,    -3,    -6,    -2,     2,     1,    -1,    -2,     2,    -2,    -5,    -5,    -1,     0,    -1,     0,    -4,    -1,     2,    -3,     0,    -1,    -1,     2,     0,     1,     2,     1,    -2,    -6,    -5,     0,     2,     0,     0,    -2,    -4,    -4,    -4,    -7,    -3,    -1,    -3,     0,    -2,     1,     0,    -2,     0,     3,     1,     0,    -1,     3,     1,     2,    -4,    -5,    -4,     0,     0,     1,    -1,    -3,    -4,    -4,     0,     1,     1,    -2,    -3,     0,    -2,    -1,    -1,    -1,     0,     3,     1,     0,     1,     2,     2,    -1,    -4,    -5,    -4,    -1,     1,     2,    -2,    -3,     1,     2,     2,    -2,    -1,    -3,     1,     0,     0,    -4,    -1,     4,     2,     0,     1,    -1,     3,     4,     3,     0,    -1,    -1,    -3,     0,     0,     1,     1,     1,     2,     0,     0,    -1,    -3,    -2,     0,     0,     0,     5,     0,     3,     1,    -1,    -1,     0,     1,     3,     2,     2,     0,    -2,    -3,    -1,     0,    -1,     2,     0,     2,     5,    -1,    -4,    -5,    -2,     0,     0,    -1,     0,    -3,    -2,    -3,     1,     0,    -1,     0,    -1,    -4,    -2,    -2,    -3,    -1,    -1,     0,     1,    -1,     2,     1,     0,    -5,    -1,    -2,    -3,    -1,     0,     1,     1,    -4,     0,    -1,     0,     2,     2,    -1,     0,    -1,    -5,    -1,     0,     2,    -1,     1,     1,    -1,     1,     2,    -2,    -2,    -3,     2,    -1,    -2,    -1,     0,     1,    -3,     1,     2,     1,     2,     0,    -1,    -1,    -2,    -5,    -1,     1,     3,     0,     1,     1,     1,     3,     0,    -4,    -1,    -3,    -2,    -1,     0,     0,     0,    -3,     0,    -1,     1,     3,     0,     0,     1,     0,    -5,    -5,    -1,    -1,     3,     0,    -2,     2,     1,     2,     2,    -2,    -2,    -3,    -4,     0,    -1,     0,     0,    -1,    -1,     1,    -2,     0,     1,     0,    -2,    -4,    -1,     0,     0,     0,     1,     0,     1,     2,     2,     2,     3,    -3,    -1,     0,    -1,     0,     0,     0,     0,    -3,    -1,     0,    -1,     1,     1,     1,    -3,    -3,    -3,    -1,     0,     0,     1,    -1,     2,     1,     1,     2,     2,     2,    -2,     2,    -1,    -2,     0,     1,     1,     0,    -3,    -5,     2,     1,    -1,    -3,    -5,    -7,    -3,    -2,     0,    -1,    -1,    -1,    -2,     1,     2,     2,     3,     1,    -1,     0,     4,     1,     0,     0,     0,     0,    -2,    -3,    -3,    -1,    -1,    -1,    -5,    -6,    -3,    -3,    -2,     0,     0,     2,    -3,     0,     2,     3,     5,    -3,    -2,     0,     1,     1,     0,     1,     0,     0,    -1,    -2,     0,     0,    -1,    -2,    -3,    -4,    -3,    -2,    -1,    -3,    -2,     0,    -1,     0,    -1,     1,    -1,    -3,     0,    -3,    -2,    -1,     0,     0,     1,    -2,    -1,    -2,     0,    -1,     0,    -1,    -3,    -4,    -2,     0,    -2,    -5,     0,     1,    -1,    -3,    -6,    -3,    -4,    -5,    -2,    -3,    -2,    -2,     0,     0,     0,     0,    -1,    -2,     0,     0,    -1,    -1,    -3,    -5,    -1,    -2,    -4,    -5,    -3,    -6,    -4,    -4,    -4,    -6,    -4,    -5,    -1,    -1,     0,     0,     0,     1,    -1,     1,     0,    -1,     0,    -1,    -1,    -1,    -2,    -3,    -3,    -2,    -1,    -2,     0,    -3,    -4,    -3,    -2,    -3,    -2,    -3,    -1,     0,     0,     0,     0),
		    95 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,     0,     0,    -1,     1,     0,     0,     0,     0,     1,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,    -2,    -2,    -2,    -2,    -3,    -2,    -1,     1,     0,     0,     0,     1,     2,     1,     1,     2,    -1,     0,     0,     0,     0,     0,    -1,     1,     0,    -1,    -3,    -4,    -1,     0,     2,     1,     2,     4,     5,     2,    -1,    -3,     4,    -1,    -1,     1,    -1,    -2,    -2,     1,     1,     0,     0,     0,    -1,     0,    -2,    -2,     2,     0,    -3,     3,     0,     2,     2,    -2,    -3,    -1,     1,    -1,     1,     3,    -2,     1,     2,     3,     5,     5,     2,    -1,     0,     0,    -1,     0,     0,     1,    -1,    -3,     0,     4,     4,     0,    -3,    -3,    -2,    -1,     2,     0,     1,     0,     1,     2,     3,     2,     4,     3,     3,    -1,     0,    -1,    -1,    -1,     1,     1,    -2,    -1,     3,     1,     1,    -3,    -3,    -1,     1,     4,     1,     3,     2,    -1,     1,     2,     3,    -1,     2,     2,     3,     0,     0,     0,     0,    -2,     0,     0,    -2,     2,     2,     3,     2,     0,    -3,    -1,     3,     3,     5,     4,     1,     1,     1,     1,    -1,    -2,    -2,     2,     2,     1,     0,     0,    -3,    -3,    -3,    -2,     0,     1,     4,     3,     3,    -2,    -1,    -3,    -1,     1,    -1,     1,     1,    -2,    -1,    -3,    -2,    -2,    -2,    -2,     4,     1,     0,    -1,    -3,    -3,    -2,    -1,     0,     1,     2,     2,     1,     2,    -4,    -6,    -6,    -8,    -9,   -11,    -6,    -8,    -8,    -7,    -5,    -4,    -4,    -2,     4,     2,     0,     0,    -1,    -3,    -1,     0,    -1,     0,     2,     2,     1,    -1,    -4,    -5,    -6,    -5,    -5,    -9,   -10,    -9,   -11,   -10,    -9,    -4,    -2,    -1,     1,     2,     0,     0,     0,    -1,     0,    -1,     0,    -1,     1,     1,    -2,    -1,    -1,    -2,     0,     1,     2,     0,    -3,    -3,    -5,    -6,    -7,    -6,    -4,    -1,     0,     1,     0,     0,     0,     2,     0,     2,     2,     1,     3,     0,     2,     0,    -1,    -2,    -2,     1,     1,     1,     1,    -1,     0,     1,    -3,    -2,    -3,    -2,     0,     0,     0,     0,     0,     1,     2,     1,    -2,    -1,    -1,     1,     0,     1,    -1,    -2,    -2,    -3,     0,     0,     1,     0,     0,     0,     1,     2,    -1,    -1,    -2,    -3,     0,    -1,    -1,     0,     3,     1,     3,     0,    -1,     2,     0,    -1,    -1,    -3,    -2,     0,    -1,    -2,    -1,    -2,     0,    -1,     2,     1,     5,    -2,    -3,    -2,     0,     1,    -1,    -4,    -3,    -4,     1,    -3,     0,    -1,     2,     2,    -1,    -1,    -2,    -2,    -1,    -4,    -2,     0,     1,    -1,     0,     0,     4,     0,    -3,    -3,    -1,    -1,     0,    -2,    -4,    -3,    -2,    -1,    -2,     1,     1,     0,    -1,    -2,     0,    -1,    -1,    -2,    -4,    -2,    -1,     1,     1,     1,     0,    -2,    -5,    -4,     0,    -1,    -2,     2,     0,    -2,     1,     0,    -2,    -1,     0,     0,     0,    -2,    -3,    -4,    -2,    -2,    -1,     2,     1,     1,     1,     0,     0,     0,    -5,    -4,     0,     0,     2,     3,    -1,     1,    -1,     0,     0,    -3,     0,    -1,    -2,    -3,    -6,    -3,    -3,    -3,    -1,     0,     0,     2,    -2,    -2,     0,     0,    -5,    -4,     0,     0,     4,     3,     1,     0,    -2,    -3,    -5,    -3,    -2,    -4,    -2,    -7,    -3,    -4,    -4,     1,     1,     2,     3,     1,     0,    -2,     3,     0,    -1,    -3,     0,     0,     2,     2,     2,    -1,    -2,    -2,    -2,     0,    -1,    -1,    -1,     1,    -1,     2,     1,     2,     2,     1,     0,     1,     0,    -1,    -1,    -1,    -3,     0,    -1,     0,    -1,     1,     2,     0,     1,     0,    -2,    -4,     0,    -1,    -1,     0,    -2,     3,     1,     3,     1,    -1,     0,     2,     2,     3,     1,     3,    -1,     0,     0,     0,    -2,     1,    -1,     1,     0,    -1,    -1,    -2,    -3,    -1,    -1,    -1,    -2,     2,     2,     1,     1,     0,     0,     0,     1,     5,     1,     5,     5,     0,     0,    -1,     2,     2,     0,     0,    -1,    -1,     2,     0,    -1,     0,    -1,     0,     1,    -1,    -1,    -1,    -1,    -2,     3,     1,     3,     2,     1,     4,     6,    -1,     0,     0,     0,     2,     3,     2,     3,    -1,    -1,     2,    -1,    -2,     0,     2,     1,     3,    -3,     0,     0,     1,     1,     1,    -1,    -4,    -1,    -1,    -1,     0,    -1,     0,     1,     3,    -3,    -2,     4,     2,     3,     4,     3,    -1,     4,     3,     3,     2,    -2,     0,     2,     3,     3,     2,     5,     3,     2,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,     0,     0,     1,     0,     3,     2,     1,    -5,    -2,    -1,     1,    -3,    -2,     1,    -1,    -1,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,    -1,    -2,    -3,    -3,     0,     0,     0,     0,     0),
		    96 => (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     3,     3,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     1,     1,     2,     4,     2,     2,     1,     4,     5,    -2,     1,     2,     3,     3,     1,     3,     1,     1,     1,     0,     0,     0,     0,     0,     0,     0,     0,     4,     4,     3,     3,     1,     2,     3,     4,     6,     4,     2,     2,     3,     3,     1,     0,     1,    -1,    -1,    -1,     1,     1,     0,     0,     0,     0,     0,     5,     0,     1,     4,     5,     3,     2,     3,     1,     1,     5,     3,     2,    -1,    -3,    -2,     0,     1,    -2,    -1,    -1,     0,    -1,     0,     0,     0,     0,    -1,     6,     0,     4,     3,     0,     0,     1,     1,     1,     2,     0,     0,    -2,    -2,    -1,    -1,    -2,    -5,    -3,    -4,    -4,    -4,    -3,     0,     1,     0,     0,    -1,    -1,     2,     1,     0,    -2,    -2,     1,     1,     0,     3,     0,    -4,     0,    -4,    -1,    -2,    -3,    -5,    -6,    -7,    -5,    -3,    -2,     1,     1,     0,    -1,    -1,    -3,     1,    -1,    -2,    -4,    -3,     3,     1,     2,     2,     0,    -1,    -4,    -3,    -4,    -7,    -7,    -5,    -7,    -7,    -6,    -3,    -1,     0,    -2,     0,     0,     0,    -4,     2,     1,    -3,    -4,     0,     0,     2,     2,     1,     0,    -3,    -5,    -7,    -7,    -9,    -6,    -4,    -1,    -7,    -7,    -5,    -2,     1,    -3,     0,     0,     0,    -3,     2,     0,    -1,    -1,     2,     1,     0,     0,    -1,     0,    -6,   -10,    -7,    -4,    -4,     0,     0,     1,    -2,    -4,    -5,    -4,     0,    -3,     0,    -1,     0,    -1,     3,    -1,    -2,    -1,     2,    -1,    -1,     1,     0,    -7,    -4,    -3,    -1,     0,     0,     3,     4,     3,     2,     1,     0,    -4,    -3,    -1,     0,    -1,     0,    -1,     1,     1,    -2,     0,     2,    -2,     1,    -1,    -1,    -7,    -5,     0,     1,     3,     3,     1,     2,     1,    -1,     0,     1,    -1,    -4,    -5,     0,     1,    -1,    -2,     2,     2,    -3,     1,     0,    -1,    -1,    -2,    -3,    -6,    -3,     0,     2,     2,     2,     2,     2,     0,     0,    -1,     1,     0,    -2,    -2,     0,     0,    -1,    -3,     1,     0,    -1,     0,     1,    -1,    -1,    -1,    -3,    -2,     2,    -2,     2,    -1,     2,     2,     2,     1,     3,     2,     3,     1,    -3,    -3,     0,     0,    -1,    -3,    -1,     2,     1,    -2,     0,    -1,     1,    -3,    -5,    -1,     0,     0,     2,     0,    -3,     2,     0,     2,     2,     4,     3,     1,    -2,     1,     0,     0,    -1,    -3,    -2,     1,     3,    -1,     2,    -1,     1,     0,    -2,     0,     0,     2,     1,     0,     3,    -2,     1,     1,     3,     3,     1,     6,    -1,     0,     0,     0,    -1,    -2,    -3,    -1,     3,     0,     0,     0,     0,     0,    -1,     2,     2,     1,    -1,    -1,     1,    -2,     1,     2,    -1,     0,     1,     4,     0,    -4,     0,     0,    -1,    -3,    -1,     0,     2,     0,    -1,     0,     2,     3,    -2,     0,     2,     0,     1,     0,    -3,     1,    -1,     0,    -2,     1,     3,     4,     0,    -2,     0,     0,     0,    -3,    -2,    -1,     0,    -1,     2,    -2,     0,    -2,    -1,     1,     2,     2,    -1,    -2,    -2,     0,    -3,    -1,    -1,     0,     4,     4,     0,    -2,     1,     0,     0,    -3,     2,    -1,    -3,     1,     0,    -2,    -5,    -3,    -2,     0,     1,    -1,    -1,     0,    -1,    -1,    -1,    -1,     1,     2,     2,     1,    -1,    -1,     0,    -1,     0,    -1,     3,    -2,    -2,     1,     1,     0,     0,    -3,    -3,    -2,     3,     2,     2,    -1,    -3,    -1,     0,    -1,    -1,     0,     0,     2,    -2,     0,     0,    -1,     0,    -2,     2,     0,    -3,    -1,    -3,    -1,     1,    -2,    -3,    -1,     1,     5,     3,     1,     3,    -2,     2,    -1,    -2,    -3,    -1,     2,     0,     0,     0,     0,     0,    -1,     1,     0,     0,     1,    -2,    -1,    -1,    -2,    -3,     1,     2,     2,     1,     1,    -2,    -3,     1,    -2,    -1,    -3,    -3,     0,     1,     0,     1,     0,    -1,    -1,    -1,     0,     1,    -3,    -6,    -4,    -3,    -5,    -2,     0,     0,    -2,    -3,    -1,    -2,    -3,    -2,    -5,    -5,    -5,    -6,    -1,     1,     0,     0,     0,     0,    -1,    -1,     0,    -1,    -2,    -2,    -5,    -6,    -5,    -4,    -1,    -1,    -4,    -8,    -8,    -7,    -4,    -1,    -4,    -4,    -3,    -5,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,     0,     0,     1,     0,    -2,    -4,    -4,    -5,    -2,    -4,    -5,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -4,    -2,    -2,    -2,    -1,     1,     0,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -1,     0,    -1,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,    -1),
		    97 => (    0,     0,     1,    -1,     1,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     0,    -1,     0,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -3,    -4,     0,    -1,     0,     0,     0,     0,    -1,     0,     0,     0,     1,     0,    -1,    -1,    -1,     0,     0,    -1,    -1,    -2,    -2,    -5,    -1,     0,    -1,    -2,    -1,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -3,    -3,    -6,    -6,    -5,    -6,    -7,    -6,    -7,    -4,    -2,    -1,    -1,     0,    -2,    -3,    -3,    -5,    -1,    -1,    -1,     0,     0,     0,     0,    -1,    -1,    -3,    -5,    -5,    -5,    -8,    -9,    -8,    -4,    -4,    -4,    -4,    -3,    -6,    -4,    -3,    -3,    -3,    -2,    -4,    -7,    -7,    -4,    -1,     1,     0,     0,     0,    -4,    -7,     1,    -3,    -1,     1,     1,    -2,    -2,     0,     2,     3,     0,     3,     1,     0,    -3,    -6,    -4,    -2,    -8,    -5,    -7,    -3,     0,     0,     0,     2,     2,     2,    -2,    -2,    -1,    -2,     0,    -1,     0,     1,     0,     1,     2,    -1,    -1,    -1,     1,     3,     2,     2,    -3,    -5,    -4,    -4,    -2,    -1,     3,     3,     1,     2,    -3,    -1,     1,    -1,     0,    -1,     1,     1,     1,     1,    -1,    -1,     5,     0,    -1,     0,     0,    -1,    -1,     0,    -4,    -5,    -3,    -3,     6,     1,     0,     1,     0,    -2,     1,     1,     3,     2,     1,     0,    -1,    -2,     0,    -1,     2,     3,     1,     2,     0,    -2,    -2,    -2,    -6,    -7,    -2,     1,     3,    -1,     1,     2,     1,     2,     1,     2,     4,     4,     1,    -3,    -1,     1,     1,     0,     2,     2,     0,     2,     0,     1,    -2,    -3,    -1,     0,     6,     0,     3,     2,     0,     2,     2,     0,     2,     3,     2,     2,    -2,    -4,    -1,     2,     4,     2,     0,     2,     1,     3,     0,    -1,    -2,    -2,     2,     0,     5,     0,     0,     4,     1,    -1,     0,     0,     1,     2,     1,    -2,    -2,     2,     3,     6,     4,     3,     0,     2,    -1,     1,    -2,     0,     1,     1,    -5,    -3,     3,     0,     2,     4,     1,    -2,    -2,     0,     0,     2,     0,     1,     3,     3,     3,     6,     5,     3,     2,     0,    -3,    -1,     0,     4,     0,     1,     3,     2,     3,     0,     1,     4,     0,    -3,    -2,     1,     0,     0,     1,     0,     2,     3,     2,     6,     4,     3,     1,    -3,    -2,    -4,    -1,     1,    -1,     0,     3,    -1,    -2,    -1,     1,     2,    -3,    -4,     0,    -1,    -2,     0,     1,    -1,     1,     0,     1,     4,     1,     1,     2,    -1,    -1,    -2,    -4,    -1,     1,     2,    -3,    -3,     0,     0,     0,     1,    -2,    -3,    -1,     0,    -1,    -4,    -4,    -2,    -1,    -2,     0,    -1,    -2,     0,     1,     4,    -1,     1,     0,     3,     2,     2,     1,    -1,    -2,     0,    -1,     0,    -2,    -1,     0,     0,    -1,     0,     2,     2,    -2,    -4,    -2,    -2,    -1,    -1,     4,     7,     5,     1,     4,     3,     4,     3,    -3,    -3,    -2,     0,    -1,    -1,    -1,     0,     1,     0,    -2,     0,     0,     0,    -3,    -5,    -2,     0,     0,     3,     5,     6,     1,     3,     2,     4,     3,     0,     2,    -1,    -3,     1,     0,     1,    -1,     0,     2,     2,    -1,    -2,    -3,    -1,    -2,    -3,    -2,    -1,     0,     1,     6,     4,     2,     1,     1,     2,     1,     0,     1,     0,    -2,    -1,     1,     0,     0,     1,     1,     1,     1,     1,    -3,    -1,    -1,    -2,    -3,    -2,    -2,     4,     7,     2,     2,     0,     1,     0,     0,     2,    -1,    -3,    -1,     0,     2,    -1,    -2,    -4,     1,     0,     2,     1,     0,    -1,    -1,    -2,     0,     0,     1,     0,     1,     0,     0,     0,     0,    -2,    -1,     2,    -2,    -3,     0,     0,     0,     0,    -1,    -3,     2,     2,     2,     1,     3,     2,     0,     1,     1,    -1,     1,     0,    -2,    -3,    -2,    -1,     1,    -1,    -1,    -3,    -2,    -1,     0,     0,     0,    -2,    -3,    -3,     1,     4,     2,     0,     0,     1,    -1,     1,     1,    -1,    -3,     0,    -3,    -3,    -3,    -3,    -2,    -5,    -4,    -3,     0,    -3,     0,     0,     1,    -1,    -5,    -3,     2,     4,     2,     1,     0,     3,     0,    -1,     0,    -5,    -4,    -2,    -4,    -5,    -4,    -3,    -3,    -5,    -5,    -2,     0,    -2,     0,     0,     0,     0,    -1,     0,     3,     1,     2,     0,     0,     0,     1,     0,     0,    -3,    -3,    -2,    -2,    -5,    -5,    -4,    -1,    -4,    -5,    -3,    -2,     0,     1,     0,    -1,    -2,     3,     0,     0,     0,     1,    -2,     1,     1,    -1,    -1,     1,    -4,    -4,     0,    -3,    -4,    -5,    -3,    -1,     0,    -3,    -1,    -1,     0,     0,    -1,     0,     0,    -3,    -2,    -3,    -2,    -2,     0,     4,    -1,    -1,     0,     0,     0,     1,    -1,    -3,    -1,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,     0,     1,    -1,     0,     1,     2,     0,    -2,    -1,     0,     0,    -3,    -1,    -1,    -3,     1,     0,     4,     1,    -1,     0,     2,     0,     2,     0,     0,     0,     0),
		    98 => (    0,     0,     0,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,     1,     0,     0,     1,     0,     0,     0,     0,     0,    -1,    -1,    -1,    -2,    -2,    -2,    -1,     1,    -1,    -1,     0,    -1,     0,     0,     0,     0,     0,     1,    -1,     0,     0,     0,     0,     0,    -1,    -4,    -5,    -5,    -2,     0,    -1,    -3,    -3,    -1,     0,     0,    -1,    -1,    -2,    -1,     0,     0,     0,     0,     1,     1,    -1,     0,    -1,    -2,    -1,    -6,     2,     3,     4,     2,     4,     4,     3,     1,     0,     1,    -1,    -3,    -2,    -4,    -2,     0,    -1,    -1,    -1,     0,     0,    -1,     1,    -1,    -4,    -4,    -1,     1,     1,     2,    -1,    -3,     0,    -1,    -1,    -1,     0,     0,     0,     1,     0,     1,    -4,    -2,    -1,     0,     0,    -1,     0,     0,     0,    -3,    -4,    -7,    -2,     1,     2,    -2,     0,     1,    -3,    -2,     2,     0,     1,     2,     1,     0,     2,     0,    -2,    -2,    -2,    -1,     1,    -1,     0,     0,    -4,    -2,    -2,    -2,     0,     5,     3,     2,     2,     1,     0,     1,     1,     2,     2,     0,    -2,     2,    -1,     0,    -2,    -1,    -2,    -2,     0,     0,    -1,    -2,    -1,    -3,    -1,     0,     3,     4,    -3,    -1,     1,    -2,    -1,    -2,    -2,    -1,    -2,     0,     0,     1,    -1,    -3,    -2,    -2,    -1,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -4,    -4,     1,     5,    -2,    -1,     2,     1,    -1,    -3,    -3,    -1,    -5,     1,     0,     1,    -1,    -1,    -1,    -3,     0,     1,     2,     0,     0,     0,    -1,    -1,    -5,    -4,    -1,    -1,    -2,     0,     3,     3,     1,    -2,    -2,    -1,    -1,     2,    -3,    -1,     0,     1,    -1,    -1,    -1,     1,    -4,    -4,     0,    -1,    -2,    -2,    -2,    -5,     1,    -2,    -6,    -1,     2,     6,     6,     4,     1,     0,     0,     1,     1,    -3,     3,     2,     0,    -2,    -4,    -5,    -4,    -4,     0,    -1,    -1,    -3,    -2,    -2,     0,     0,    -2,     0,    -5,     0,     3,     5,     3,     0,    -1,    -3,    -1,    -1,    -1,    -1,    -2,    -2,    -5,    -3,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -3,    -5,    -5,    -6,    -6,     0,     0,     1,     4,     1,     0,     1,     1,     0,     1,     1,     0,    -1,    -3,    -2,    -1,     0,     0,    -1,     0,    -2,    -1,    -1,    -3,    -5,    -7,    -5,    -4,    -3,     0,     0,     2,     1,    -1,     0,    -2,    -3,     0,     1,    -4,    -3,    -2,    -2,    -1,     0,     0,     0,    -3,    -2,     1,     0,    -2,    -2,    -4,    -1,     2,     1,     1,    -1,    -2,     0,     0,     0,    -3,    -1,     2,    -1,    -3,    -3,    -2,    -4,    -2,    -1,     0,    -2,    -2,    -3,    -1,    -2,     0,    -1,     1,     0,     1,    -1,    -2,    -2,    -1,     2,    -1,    -3,     0,     0,     1,    -3,    -2,    -2,    -2,    -4,    -2,     0,    -1,    -1,    -1,    -2,     0,     2,     2,     1,     3,     1,     0,    -2,    -1,    -4,     0,    -4,     3,    -2,     2,     2,     1,    -1,    -1,    -1,    -1,    -5,    -2,     0,     0,    -2,    -4,     1,     1,    -1,     2,     2,     0,    -1,     0,    -1,    -5,    -4,    -1,    -3,    -1,     1,     3,     1,     3,     3,     0,    -2,    -2,    -1,    -3,    -1,     0,    -1,    -1,     4,     0,     1,     3,    -1,    -2,    -2,     1,    -2,    -4,    -2,    -1,    -5,    -2,     1,     2,     2,     2,     1,     1,    -4,    -2,     0,    -2,     0,    -1,    -2,     3,     3,     4,     3,     1,    -3,    -2,     0,     1,    -4,    -3,    -3,    -1,    -2,     0,    -2,     0,     1,     2,     0,    -2,    -3,    -1,    -5,    -2,    -1,     0,    -2,     0,     3,     1,     2,     1,    -1,    -4,    -1,     1,    -3,    -1,    -1,     1,     2,    -2,    -2,    -1,     2,     2,     1,    -2,    -2,     0,    -4,    -1,    -2,    -1,    -2,    -2,     1,     0,     0,     0,    -2,     0,    -1,     0,     1,    -2,     2,    -1,    -1,    -2,    -4,     1,     2,     2,    -1,    -2,    -2,    -1,    -3,    -1,    -2,    -1,    -2,    -3,    -2,     0,     4,     3,    -2,    -1,     1,     1,     2,    -2,    -1,    -3,    -2,    -1,    -2,    -1,     0,    -1,    -4,    -1,     0,     0,    -2,     0,    -1,     1,    -1,    -1,    -3,     2,     1,     3,     1,    -2,    -1,    -2,     0,     0,     0,    -1,    -1,    -3,    -1,     0,    -2,    -5,    -2,    -1,     0,     2,    -3,     0,    -1,     0,    -1,    -1,    -3,    -3,     1,     1,     1,     0,    -2,    -2,     0,     0,     1,     2,     3,    -2,     0,     0,     0,    -2,    -2,     0,    -3,     0,    -1,     0,     0,     0,     0,     0,    -1,    -2,     0,    -1,    -3,    -2,    -3,    -3,    -3,    -3,    -3,    -4,    -3,    -2,    -1,     0,     0,    -1,    -1,    -1,    -1,     0,    -1,     0,     0,    -1,     0,    -1,    -1,    -1,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -3,    -4,    -2,    -2,    -1,    -1,    -2,    -4,    -4,    -2,     0,     0,     0,     1,     0,     0,     0,     1,     0,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     0,    -2,    -1,    -1,    -1,    -1,    -1,    -1,     0,     0,     1,     0,     0,     0,    -1,     0),
		    99 => (    0,     0,     0,     0,    -1,     0,     0,    -1,    -1,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     1,     0,    -1,     0,     0,     0,     0,     0,     0,    -1,     0,     0,     1,     0,     0,     0,     0,    -1,    -1,    -2,    -2,     0,     0,     0,     0,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    -1,     0,    -1,     0,     0,    -1,     0,     0,     0,     0,     0,    -1,    -1,    -1,     0,     0,     0,    -1,     0,     0,     0,     0,    -1,    -1,    -1,    -1,    -1,    -2,    -2,    -1,     0,     0,    -1,    -1,     0,     0,    -1,    -1,    -1,    -2,    -1,    -2,    -1,    -2,    -1,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -3,     0,     0,     0,     0,    -1,    -3,    -2,    -1,    -3,    -2,    -3,    -1,    -3,    -5,    -1,     0,     0,     0,    -3,    -1,     0,     1,     0,     0,    -1,     0,     0,     0,    -1,    -1,    -1,    -1,    -2,    -3,    -3,    -4,    -5,    -3,    -1,     0,     1,    -2,    -2,    -2,    -1,     0,    -1,    -1,     0,     0,     0,     0,    -1,     0,    -1,    -2,    -2,    -3,    -1,    -2,     0,     0,     0,     0,     0,    -2,    -3,    -1,    -2,    -3,    -2,    -2,    -1,    -1,     0,    -1,    -2,     0,     0,    -1,    -1,    -1,    -2,    -4,    -5,    -5,    -2,    -2,     1,     0,     1,     0,     1,     2,    -2,    -1,    -2,    -2,    -4,    -2,     1,    -1,     0,    -1,    -1,    -2,    -2,    -1,    -1,    -3,    -3,    -4,    -5,    -3,    -3,     0,     1,     1,    -1,     0,     0,     2,    -2,    -1,     1,     0,     0,    -2,     0,     0,    -3,    -1,     0,     0,    -2,    -2,    -2,    -3,    -2,    -3,    -1,     1,    -1,     0,     1,     1,     1,     1,     4,     1,    -1,     0,     2,     1,     0,     0,     0,    -1,    -2,    -1,    -1,    -1,    -3,    -2,     0,    -1,    -2,    -3,    -1,     1,    -2,    -3,     1,     1,     1,     3,     0,     2,    -1,     2,     2,    -1,     0,    -1,    -2,    -2,    -2,    -1,    -2,     0,    -5,     3,     0,    -1,    -1,    -2,     0,     0,    -1,    -4,     0,     1,     2,     1,     0,    -2,    -3,     0,     0,     0,    -1,     0,    -1,    -3,    -3,    -1,    -1,     0,    -2,     1,     3,     2,     0,     1,     0,    -2,    -5,    -3,    -1,    -1,    -2,     0,     0,    -1,     0,    -1,     1,     0,     2,     0,    -1,    -3,    -2,    -2,     0,     0,    -2,    -1,     2,     1,     1,     2,     0,    -2,    -6,    -2,    -1,    -4,    -4,    -2,     0,     0,    -2,     0,     0,    -1,     2,     1,    -1,    -4,    -2,    -1,     0,     0,    -2,    -2,     2,     2,     2,     0,     0,    -4,    -4,    -1,    -1,    -3,    -3,    -3,    -1,    -1,    -2,     0,     1,     1,     2,    -1,    -3,    -3,    -2,     0,     0,     0,     0,    -3,     2,     3,     1,     1,     0,    -2,    -4,    -1,    -2,    -3,     0,     0,     0,     0,    -3,     0,     0,    -1,     1,     1,    -3,    -4,    -2,     0,    -1,     0,    -1,    -2,     2,     4,     2,     4,     1,     1,     1,     1,    -3,     0,     0,     0,     0,    -4,    -2,    -2,    -3,     0,    -1,     2,     2,    -3,     0,    -2,    -1,     0,    -1,    -5,     0,     0,     0,     1,     2,     4,     3,     2,     3,     2,     0,    -1,    -2,    -3,    -3,     0,    -2,    -1,    -1,     2,    -1,    -3,    -1,    -2,    -2,     0,     0,    -5,     1,    -1,    -2,     0,     1,     0,     0,     3,     1,     0,    -4,    -1,     0,    -1,    -1,     0,    -3,    -1,    -1,     2,     2,    -1,     0,    -3,    -1,    -1,    -1,    -3,     2,     0,    -3,    -2,    -2,    -3,    -3,    -1,    -1,     0,    -4,     1,     0,    -2,    -2,    -1,    -4,     0,    -2,    -1,     2,     3,     2,    -2,     0,    -1,     0,    -1,     2,     2,    -1,    -2,    -2,    -4,    -2,    -3,    -2,    -4,    -3,     1,     1,    -2,    -3,    -1,    -2,     1,     0,    -1,     2,     3,     5,    -3,     0,     0,     0,    -2,     1,     1,     0,    -2,    -2,    -2,    -3,    -2,    -1,    -1,    -2,     2,    -1,    -6,    -2,    -1,    -1,    -1,     2,    -2,     0,     1,     3,    -3,     0,     0,     0,    -2,    -1,    -3,    -1,    -1,    -2,    -1,    -2,    -1,    -2,     0,     0,     3,    -4,    -4,    -1,     0,    -1,     0,     0,     0,     0,    -1,    -3,    -1,     0,     0,     0,    -2,    -1,    -1,     0,    -1,    -1,    -1,     0,    -1,     0,     0,     0,     1,    -2,     0,     1,     0,    -1,     2,     0,     3,     1,     0,    -1,    -1,     0,     0,     0,    -1,     0,    -2,    -1,     0,     1,    -2,    -3,    -1,    -1,     0,    -1,     1,     1,     2,    -1,     0,     0,     2,     1,     2,     1,     0,    -1,    -1,     0,     0,    -1,     3,    -2,     0,     2,     1,     0,    -3,    -1,    -1,     0,    -1,    -2,     2,     2,     1,    -1,    -1,     1,     3,     2,     2,     0,    -1,    -1,     0,    -1,     0,     0,     1,     4,     2,     2,     2,     0,     0,     2,    -2,    -1,    -1,    -3,     0,     1,     0,     0,     0,     2,     3,     4,     2,     0,     1,     0,     1,     0,     0,     0,    -1,     0,    -1,    -1,     1,     3,     2,     2,     0,     1,    -1,    -2,     0,    -1,    -1,     0,    -2,    -1,    -1,     0,     1,    -1,     1,     0,     0,     0)
        );

 ---------------------------------INFO-
 -- COEF =5.3922606

 -- MIN =-15.999999
 -- MAX =10.598255

 -- SUMMIN =-1136.8025
 -- SUMMAX =826.5192
 ---------------------------------INFO-

-- Fonction d'accès à un élément de la matrice
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer;

end WeightMatrix01;


package body WeightMatrix01 is
  function get_ML01(
    framebuffer : framebuffer_ML01;
        y           : integer;
        x           : integer
    ) return integer is
    begin
        return framebuffer(y , x);
    end function;

end package body WeightMatrix01;
